module circuit ( clk, rst, input_s1, input_s2, output_s1, output_s2, Key, 
        enc_dec, done );
  input [63:0] input_s1;
  input [63:0] input_s2;
  output [63:0] output_s1;
  output [63:0] output_s2;
  input [127:0] Key;
  input clk, rst, enc_dec;
  output done;
  wire   k_0_p_0_, roundHalf_Select_Signal, roundEnd_Select_Signal,
         controller_n2, controller_n1, controller_MoreControl,
         controller_roundCounter_n6, controller_roundCounter_n5,
         controller_roundCounter_n4, controller_roundCounter_n3,
         controller_roundCounter_n2, controller_roundCounter_n1,
         controller_roundCounter_CO,
         controller_roundCounter_mux_eachroundcounter_out_1_,
         controller_roundCounter_N1,
         controller_roundCounter_counterMUX_MUXInst_0_n2,
         controller_roundCounter_counterMUX_MUXInst_2_n6,
         controller_roundCounter_counterMUX_MUXInst_3_n6,
         controller_roundCounter_Adder_inst_c3,
         controller_roundCounter_Adder_inst_c2,
         controller_roundCounter_Adder_inst_c1,
         controller_roundCounter_Adder_inst_Cout,
         controller_roundCounter_EachRoundMUX_MUXInst_0_n6,
         controller_roundCounter_EachRoundMUX_MUXInst_1_n6,
         controller_roundCounter_FA2_Cout,
         controller_roundCounter_EachRoundMUX2_MUXInst_0_n7,
         controller_roundCounter_EachRoundMUX2_MUXInst_1_n7, prince_n267,
         prince_n266, prince_n265, prince_n264, prince_n263, prince_n262,
         prince_n261, prince_n260, prince_n259, prince_n258, prince_n257,
         prince_n256, prince_n255, prince_n254, prince_n253, prince_n252,
         prince_n251, prince_n250, prince_n249, prince_n248, prince_n247,
         prince_n246, prince_n245, prince_n244, prince_n243, prince_n242,
         prince_n241, prince_n240, prince_n239, prince_n238, prince_n237,
         prince_n236, prince_n235, prince_n234, prince_n233, prince_n232,
         prince_n231, prince_n230, prince_n229, prince_n228, prince_n227,
         prince_n226, prince_n225, prince_n224, prince_n223, prince_n222,
         prince_n221, prince_n220, prince_n219, prince_n218, prince_n217,
         prince_n216, prince_n215, prince_n214, prince_n213, prince_n212,
         prince_n211, prince_n210, prince_n209, prince_n208, prince_n207,
         prince_n206, prince_n205, prince_n204, prince_n203, prince_n202,
         prince_n201, prince_n200, prince_rounds_n402, prince_rounds_n401,
         prince_rounds_n400, prince_rounds_n399, prince_rounds_n398,
         prince_rounds_n397, prince_rounds_n396, prince_rounds_n395,
         prince_rounds_n394, prince_rounds_n393, prince_rounds_n392,
         prince_rounds_n391, prince_rounds_n390, prince_rounds_n389,
         prince_rounds_n388, prince_rounds_n387, prince_rounds_n386,
         prince_rounds_n385, prince_rounds_n384, prince_rounds_n383,
         prince_rounds_n382, prince_rounds_n381, prince_rounds_n380,
         prince_rounds_n379, prince_rounds_n378, prince_rounds_n377,
         prince_rounds_n376, prince_rounds_n375, prince_rounds_n374,
         prince_rounds_n373, prince_rounds_n372, prince_rounds_n371,
         prince_rounds_n370, prince_rounds_n369, prince_rounds_n368,
         prince_rounds_n367, prince_rounds_n366, prince_rounds_n365,
         prince_rounds_n364, prince_rounds_n363, prince_rounds_n362,
         prince_rounds_n361, prince_rounds_n360, prince_rounds_n359,
         prince_rounds_n358, prince_rounds_n357, prince_rounds_n356,
         prince_rounds_n355, prince_rounds_n354, prince_rounds_n353,
         prince_rounds_n352, prince_rounds_n351, prince_rounds_n350,
         prince_rounds_n349, prince_rounds_n348, prince_rounds_n347,
         prince_rounds_n346, prince_rounds_n345, prince_rounds_n344,
         prince_rounds_n343, prince_rounds_n342, prince_rounds_n341,
         prince_rounds_n340, prince_rounds_n339, prince_rounds_n338,
         prince_rounds_n337, prince_rounds_n336, prince_rounds_n335,
         prince_rounds_n334, prince_rounds_n333,
         prince_rounds_constant_MUX_n56, prince_rounds_constant_MUX_n55,
         prince_rounds_constant_MUX_n54, prince_rounds_constant_MUX_n53,
         prince_rounds_constant_MUX_n52, prince_rounds_constant_MUX_n51,
         prince_rounds_constant_MUX_n50, prince_rounds_constant_MUX_n49,
         prince_rounds_constant_MUX_n48, prince_rounds_constant_MUX_n47,
         prince_rounds_constant_MUX_n46, prince_rounds_constant_MUX_n45,
         prince_rounds_constant_MUX_n44, prince_rounds_constant_MUX_n43,
         prince_rounds_constant_MUX_n42, prince_rounds_constant_MUX_n41,
         prince_rounds_constant_MUX_n40, prince_rounds_constant_MUX_n39,
         prince_rounds_constant_MUX_n38, prince_rounds_constant_MUX_n37,
         prince_rounds_constant_MUX_n36, prince_rounds_constant_MUX_n35,
         prince_rounds_constant_MUX_n34, prince_rounds_constant_MUX_n33,
         prince_rounds_constant_MUX_n32, prince_rounds_constant_MUX_n31,
         prince_rounds_constant_MUX_n30, prince_rounds_constant_MUX_n29,
         prince_rounds_constant_MUX_n28, prince_rounds_constant_MUX_n27,
         prince_rounds_constant_MUX_n26, prince_rounds_constant_MUX_n25,
         prince_rounds_constant_MUX_n24, prince_rounds_constant_MUX_n23,
         prince_rounds_constant_MUX_n22, prince_rounds_constant_MUX_n21,
         prince_rounds_constant_MUX_n20, prince_rounds_constant_MUX_n19,
         prince_rounds_constant_MUX_n18, prince_rounds_constant_MUX_n17,
         prince_rounds_constant_MUX_n16, prince_rounds_constant_MUX_n15,
         prince_rounds_constant_MUX_n14, prince_rounds_constant_MUX_n13,
         prince_rounds_constant_MUX_n12, prince_rounds_constant_MUX_n11,
         prince_rounds_constant_MUX_n10, prince_rounds_constant_MUX_n9,
         prince_rounds_constant_MUX_n8,
         prince_rounds_roundResult_Reg_s1_SFF_0_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_1_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_2_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_3_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_4_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_5_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_6_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_7_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_8_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_9_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_10_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_11_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_12_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_13_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_14_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_15_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_16_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_17_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_18_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_19_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_20_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_21_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_22_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_23_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_24_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_25_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_26_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_27_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_28_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_29_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_30_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_31_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_32_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_33_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_34_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_35_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_36_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_37_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_38_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_39_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_40_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_41_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_42_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_43_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_44_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_45_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_46_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_47_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_48_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_49_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_50_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_51_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_52_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_53_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_54_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_55_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_56_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_57_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_58_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_59_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_60_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_61_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_62_SFFInst_N3,
         prince_rounds_roundResult_Reg_s1_SFF_63_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_0_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_1_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_2_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_3_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_4_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_5_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_6_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_7_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_8_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_9_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_10_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_11_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_12_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_13_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_14_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_15_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_16_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_17_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_18_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_19_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_20_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_21_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_22_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_23_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_24_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_25_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_26_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_27_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_28_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_29_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_30_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_31_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_32_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_33_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_34_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_35_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_36_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_37_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_38_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_39_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_40_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_41_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_42_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_43_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_44_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_45_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_46_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_47_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_48_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_49_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_50_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_51_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_52_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_53_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_54_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_55_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_56_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_57_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_58_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_59_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_60_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_61_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_62_SFFInst_N3,
         prince_rounds_roundResult_Reg_s2_SFF_63_SFFInst_N3,
         prince_rounds_MUX_inst0_n11, prince_rounds_MUX_inst0_n10,
         prince_rounds_MUX_inst0_n9, prince_rounds_MUX_inst0_n8,
         prince_rounds_MUX_inst1_n12, prince_rounds_MUX_inst1_n11,
         prince_rounds_MUX_inst1_n10, prince_rounds_MUX_inst1_n9,
         prince_rounds_MUX_inst1_n8,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n53,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n52,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n51,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n49,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n48,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n47,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n46,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n45,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n44,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n43,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n42,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n41,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n40,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n39,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n38,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n37,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n36,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n35,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n34,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n33,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n32,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n31,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n30,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n28,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n27,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n26,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n25,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n24,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n23,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n22,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n14,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n13,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n12,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n11,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n10,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n9,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n8,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n7,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n29,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n28,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n27,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n26,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n25,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n24,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n23,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n22,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n14,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n13,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n12,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n11,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n10,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n9,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n8,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n7,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n32,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n31,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n30,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n29,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n28,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n27,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n26,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n25,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n24,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n23,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n22,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n14,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n13,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n12,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n11,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n10,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n9,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n8,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n7,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n32,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n31,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n30,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n29,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n28,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n27,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n26,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n25,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n24,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n23,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n22,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n14,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n13,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n12,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n11,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n10,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n9,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n8,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n7,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n31,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n30,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n29,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n28,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n27,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n26,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n25,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n24,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n23,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n22,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n14,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n13,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n12,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n11,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n10,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n9,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n8,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n7,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n2,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n1,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n55,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n54,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n53,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n52,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n50,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n49,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n48,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n47,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n46,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n45,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n44,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n43,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n42,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n41,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n40,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n39,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n38,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n37,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n36,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n35,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n30,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n29,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n28,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n27,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n26,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n25,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n24,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n23,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n22,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n14,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n13,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n12,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n11,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n10,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n9,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n8,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n7,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n2,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n1,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_n2,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_n1,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n66,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n65,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n64,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n63,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n62,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n61,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n60,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n59,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n58,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n57,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n56,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n107,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n106,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n105,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n104,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n103,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n102,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n101,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n100,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n99,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n98,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n97,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n96,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n95,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n94,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n93,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n92,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n91,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n90,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n89,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n87,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n86,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n85,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n84,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n83,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n82,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n81,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n80,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n79,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n78,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n77,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n76,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n75,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n74,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n73,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n72,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n71,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n70,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n69,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n68,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n67,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_0_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_1_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_2_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_3_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_4_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_5_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_6_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_7_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_8_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_9_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_10_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_11_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_12_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_13_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_14_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_15_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_16_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_17_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_18_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_19_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_20_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_21_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_22_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_23_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_24_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_25_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_26_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_27_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_28_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_29_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_30_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_31_SFFInst_N3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_n5,
         prince_rounds_mul_s1_n32, prince_rounds_mul_s1_n31,
         prince_rounds_mul_s1_n30, prince_rounds_mul_s1_n29,
         prince_rounds_mul_s1_n28, prince_rounds_mul_s1_n27,
         prince_rounds_mul_s1_n26, prince_rounds_mul_s1_n25,
         prince_rounds_mul_s1_n24, prince_rounds_mul_s1_n23,
         prince_rounds_mul_s1_n22, prince_rounds_mul_s1_n21,
         prince_rounds_mul_s1_n20, prince_rounds_mul_s1_n19,
         prince_rounds_mul_s1_n18, prince_rounds_mul_s1_n17,
         prince_rounds_mul_s1_n16, prince_rounds_mul_s1_n15,
         prince_rounds_mul_s1_n14, prince_rounds_mul_s1_n13,
         prince_rounds_mul_s1_n12, prince_rounds_mul_s1_n11,
         prince_rounds_mul_s1_n10, prince_rounds_mul_s1_n9,
         prince_rounds_mul_s1_n8, prince_rounds_mul_s1_n7,
         prince_rounds_mul_s1_n6, prince_rounds_mul_s1_n5,
         prince_rounds_mul_s1_n4, prince_rounds_mul_s1_n3,
         prince_rounds_mul_s1_n2, prince_rounds_mul_s1_n1,
         prince_rounds_mul_s2_n96, prince_rounds_mul_s2_n95,
         prince_rounds_mul_s2_n94, prince_rounds_mul_s2_n93,
         prince_rounds_mul_s2_n92, prince_rounds_mul_s2_n91,
         prince_rounds_mul_s2_n90, prince_rounds_mul_s2_n89,
         prince_rounds_mul_s2_n88, prince_rounds_mul_s2_n87,
         prince_rounds_mul_s2_n86, prince_rounds_mul_s2_n85,
         prince_rounds_mul_s2_n84, prince_rounds_mul_s2_n83,
         prince_rounds_mul_s2_n82, prince_rounds_mul_s2_n81,
         prince_rounds_mul_s2_n80, prince_rounds_mul_s2_n79,
         prince_rounds_mul_s2_n78, prince_rounds_mul_s2_n77,
         prince_rounds_mul_s2_n76, prince_rounds_mul_s2_n75,
         prince_rounds_mul_s2_n74, prince_rounds_mul_s2_n73,
         prince_rounds_mul_s2_n72, prince_rounds_mul_s2_n71,
         prince_rounds_mul_s2_n70, prince_rounds_mul_s2_n69,
         prince_rounds_mul_s2_n68, prince_rounds_mul_s2_n67,
         prince_rounds_mul_s2_n66, prince_rounds_mul_s2_n65;
  wire   [2:0] round_Signal;
  wire   [1:0] controller_roundCounter_zero_or_PlusOne;
  wire   [1:0] controller_roundCounter_feedback1;
  wire   [3:0] controller_roundCounter_zero_or_PlusOne_count;
  wire   [3:0] controller_roundCounter_CountPlusOne;
  wire   [3:1] controller_roundCounter_mux_count_out;
  wire   [1:0] controller_roundCounter_eachroundcounter;
  wire   [63:0] prince_SR_Inv_Result_s1;
  wire   [63:0] prince_rounds_mul_input_s2;
  wire   [63:0] prince_rounds_mul_input_s1;
  wire   [63:0] prince_rounds_SR_Inv_Result_s1;
  wire   [63:0] prince_rounds_sub_Inv_Result_s1;
  wire   [63:0] prince_rounds_Sbox_Input_s2;
  wire   [63:0] prince_rounds_Sbox_Input_s1;
  wire   [63:0] prince_rounds_round_inputXORkeyRCON_s1;
  wire   [63:0] prince_rounds_SR_Result_s2;
  wire   [63:0] prince_rounds_SR_Result_s1;
  wire   [63:0] prince_rounds_mul_result_s2;
  wire   [63:0] prince_rounds_mul_result_s1;
  wire   [63:1] prince_rounds_round_Constant;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_0_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_1_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_2_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_3_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_4_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_5_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_6_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_7_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_8_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_9_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_10_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_11_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_12_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_13_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_14_e_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_h_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_g_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_f_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_e_si;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_h_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_g_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_f_s;
  wire   [8:1] prince_rounds_sub_sBoxCombined_PRINCE_15_e_s;

  XOR2_X1 keys_U1 ( .A(Key[65]), .B(Key[127]), .Z(k_0_p_0_) );
  AND2_X1 controller_U4 ( .A1(round_Signal[0]), .A2(controller_n2), .ZN(done)
         );
  NOR2_X1 controller_U3 ( .A1(round_Signal[1]), .A2(controller_n1), .ZN(
        controller_n2) );
  NAND2_X1 controller_U2 ( .A1(round_Signal[2]), .A2(roundEnd_Select_Signal), 
        .ZN(controller_n1) );
  OR2_X1 controller_U1 ( .A1(roundEnd_Select_Signal), .A2(
        controller_MoreControl), .ZN(roundHalf_Select_Signal) );
  OR2_X1 controller_roundCounter_U10 ( .A1(controller_MoreControl), .A2(
        controller_roundCounter_n6), .ZN(controller_roundCounter_N1) );
  NOR2_X1 controller_roundCounter_U9 ( .A1(
        controller_roundCounter_eachroundcounter[0]), .A2(
        controller_roundCounter_n5), .ZN(controller_roundCounter_n6) );
  NAND2_X1 controller_roundCounter_U8 ( .A1(
        controller_roundCounter_eachroundcounter[1]), .A2(
        controller_roundCounter_n4), .ZN(controller_roundCounter_n5) );
  NOR2_X1 controller_roundCounter_U7 ( .A1(controller_roundCounter_n4), .A2(
        controller_roundCounter_n3), .ZN(controller_MoreControl) );
  NAND2_X1 controller_roundCounter_U6 ( .A1(
        controller_roundCounter_eachroundcounter[1]), .A2(
        controller_roundCounter_eachroundcounter[0]), .ZN(
        controller_roundCounter_n3) );
  NAND2_X1 controller_roundCounter_U5 ( .A1(round_Signal[1]), .A2(
        controller_roundCounter_n2), .ZN(controller_roundCounter_n4) );
  NOR2_X1 controller_roundCounter_U4 ( .A1(roundEnd_Select_Signal), .A2(
        controller_roundCounter_n1), .ZN(controller_roundCounter_n2) );
  NAND2_X1 controller_roundCounter_U3 ( .A1(round_Signal[2]), .A2(
        round_Signal[0]), .ZN(controller_roundCounter_n1) );
  NOR2_X1 controller_roundCounter_counterMUX_MUXInst_0_U2 ( .A1(rst), .A2(
        controller_roundCounter_counterMUX_MUXInst_0_n2), .ZN(
        controller_roundCounter_Adder_inst_c1) );
  INV_X1 controller_roundCounter_counterMUX_MUXInst_0_U1 ( .A(round_Signal[0]), 
        .ZN(controller_roundCounter_counterMUX_MUXInst_0_n2) );
  OR2_X1 controller_roundCounter_counterMUX_MUXInst_1_U1 ( .A1(round_Signal[1]), .A2(rst), .ZN(controller_roundCounter_mux_count_out[1]) );
  NOR2_X1 controller_roundCounter_counterMUX_MUXInst_2_U2 ( .A1(rst), .A2(
        controller_roundCounter_counterMUX_MUXInst_2_n6), .ZN(
        controller_roundCounter_mux_count_out[2]) );
  INV_X1 controller_roundCounter_counterMUX_MUXInst_2_U1 ( .A(round_Signal[2]), 
        .ZN(controller_roundCounter_counterMUX_MUXInst_2_n6) );
  NOR2_X1 controller_roundCounter_counterMUX_MUXInst_3_U2 ( .A1(rst), .A2(
        controller_roundCounter_counterMUX_MUXInst_3_n6), .ZN(
        controller_roundCounter_mux_count_out[3]) );
  INV_X1 controller_roundCounter_counterMUX_MUXInst_3_U1 ( .A(
        roundEnd_Select_Signal), .ZN(
        controller_roundCounter_counterMUX_MUXInst_3_n6) );
  INV_X1 controller_roundCounter_Adder_inst_FA1_U1 ( .A(
        controller_roundCounter_Adder_inst_c1), .ZN(
        controller_roundCounter_CountPlusOne[0]) );
  XOR2_X1 controller_roundCounter_Adder_inst_FA2_U2 ( .A(
        controller_roundCounter_mux_count_out[1]), .B(
        controller_roundCounter_Adder_inst_c1), .Z(
        controller_roundCounter_CountPlusOne[1]) );
  AND2_X1 controller_roundCounter_Adder_inst_FA2_U1 ( .A1(
        controller_roundCounter_mux_count_out[1]), .A2(
        controller_roundCounter_Adder_inst_c1), .ZN(
        controller_roundCounter_Adder_inst_c2) );
  XOR2_X1 controller_roundCounter_Adder_inst_FA3_U2 ( .A(
        controller_roundCounter_mux_count_out[2]), .B(
        controller_roundCounter_Adder_inst_c2), .Z(
        controller_roundCounter_CountPlusOne[2]) );
  AND2_X1 controller_roundCounter_Adder_inst_FA3_U1 ( .A1(
        controller_roundCounter_mux_count_out[2]), .A2(
        controller_roundCounter_Adder_inst_c2), .ZN(
        controller_roundCounter_Adder_inst_c3) );
  XOR2_X1 controller_roundCounter_Adder_inst_FA4_U2 ( .A(
        controller_roundCounter_mux_count_out[3]), .B(
        controller_roundCounter_Adder_inst_c3), .Z(
        controller_roundCounter_CountPlusOne[3]) );
  AND2_X1 controller_roundCounter_Adder_inst_FA4_U1 ( .A1(
        controller_roundCounter_mux_count_out[3]), .A2(
        controller_roundCounter_Adder_inst_c3), .ZN(
        controller_roundCounter_Adder_inst_Cout) );
  MUX2_X1 controller_roundCounter_EachRoundMUX3_MUXInst_0_U1 ( .A(
        controller_roundCounter_Adder_inst_c1), .B(
        controller_roundCounter_CountPlusOne[0]), .S(
        controller_roundCounter_N1), .Z(
        controller_roundCounter_zero_or_PlusOne_count[0]) );
  MUX2_X1 controller_roundCounter_EachRoundMUX3_MUXInst_1_U1 ( .A(
        controller_roundCounter_mux_count_out[1]), .B(
        controller_roundCounter_CountPlusOne[1]), .S(
        controller_roundCounter_N1), .Z(
        controller_roundCounter_zero_or_PlusOne_count[1]) );
  MUX2_X1 controller_roundCounter_EachRoundMUX3_MUXInst_2_U1 ( .A(
        controller_roundCounter_mux_count_out[2]), .B(
        controller_roundCounter_CountPlusOne[2]), .S(
        controller_roundCounter_N1), .Z(
        controller_roundCounter_zero_or_PlusOne_count[2]) );
  MUX2_X1 controller_roundCounter_EachRoundMUX3_MUXInst_3_U1 ( .A(
        controller_roundCounter_mux_count_out[3]), .B(
        controller_roundCounter_CountPlusOne[3]), .S(
        controller_roundCounter_N1), .Z(
        controller_roundCounter_zero_or_PlusOne_count[3]) );
  DFF_X1 controller_roundCounter_Inst_Reg_s_current_state_reg_0_ ( .D(
        controller_roundCounter_zero_or_PlusOne_count[0]), .CK(clk), .Q(
        round_Signal[0]), .QN());
  DFF_X1 controller_roundCounter_Inst_Reg_s_current_state_reg_1_ ( .D(
        controller_roundCounter_zero_or_PlusOne_count[1]), .CK(clk), .Q(
        round_Signal[1]), .QN());
  DFF_X1 controller_roundCounter_Inst_Reg_s_current_state_reg_2_ ( .D(
        controller_roundCounter_zero_or_PlusOne_count[2]), .CK(clk), .Q(
        round_Signal[2]), .QN());
  DFF_X1 controller_roundCounter_Inst_Reg_s_current_state_reg_3_ ( .D(
        controller_roundCounter_zero_or_PlusOne_count[3]), .CK(clk), .Q(
        roundEnd_Select_Signal), .QN());
  INV_X1 controller_roundCounter_EachRoundMUX_MUXInst_0_U2 ( .A(
        controller_roundCounter_feedback1[0]), .ZN(
        controller_roundCounter_EachRoundMUX_MUXInst_0_n6) );
  NOR2_X1 controller_roundCounter_EachRoundMUX_MUXInst_0_U1 ( .A1(rst), .A2(
        controller_roundCounter_EachRoundMUX_MUXInst_0_n6), .ZN(
        controller_roundCounter_CO) );
  INV_X1 controller_roundCounter_EachRoundMUX_MUXInst_1_U2 ( .A(
        controller_roundCounter_feedback1[1]), .ZN(
        controller_roundCounter_EachRoundMUX_MUXInst_1_n6) );
  NOR2_X1 controller_roundCounter_EachRoundMUX_MUXInst_1_U1 ( .A1(rst), .A2(
        controller_roundCounter_EachRoundMUX_MUXInst_1_n6), .ZN(
        controller_roundCounter_mux_eachroundcounter_out_1_) );
  INV_X1 controller_roundCounter_FA1_U1 ( .A(controller_roundCounter_CO), .ZN(
        controller_roundCounter_eachroundcounter[0]) );
  AND2_X1 controller_roundCounter_FA2_U2 ( .A1(
        controller_roundCounter_mux_eachroundcounter_out_1_), .A2(
        controller_roundCounter_CO), .ZN(controller_roundCounter_FA2_Cout) );
  XOR2_X1 controller_roundCounter_FA2_U1 ( .A(
        controller_roundCounter_mux_eachroundcounter_out_1_), .B(
        controller_roundCounter_CO), .Z(
        controller_roundCounter_eachroundcounter[1]) );
  NOR2_X1 controller_roundCounter_EachRoundMUX2_MUXInst_0_U2 ( .A1(
        controller_roundCounter_N1), .A2(
        controller_roundCounter_EachRoundMUX2_MUXInst_0_n7), .ZN(
        controller_roundCounter_zero_or_PlusOne[0]) );
  INV_X1 controller_roundCounter_EachRoundMUX2_MUXInst_0_U1 ( .A(
        controller_roundCounter_eachroundcounter[0]), .ZN(
        controller_roundCounter_EachRoundMUX2_MUXInst_0_n7) );
  NOR2_X1 controller_roundCounter_EachRoundMUX2_MUXInst_1_U2 ( .A1(
        controller_roundCounter_N1), .A2(
        controller_roundCounter_EachRoundMUX2_MUXInst_1_n7), .ZN(
        controller_roundCounter_zero_or_PlusOne[1]) );
  INV_X1 controller_roundCounter_EachRoundMUX2_MUXInst_1_U1 ( .A(
        controller_roundCounter_eachroundcounter[1]), .ZN(
        controller_roundCounter_EachRoundMUX2_MUXInst_1_n7) );
  DFF_X1 controller_roundCounter_Inst_Reg1_s_current_state_reg_0_ ( .D(
        controller_roundCounter_zero_or_PlusOne[0]), .CK(clk), .Q(
        controller_roundCounter_feedback1[0]), .QN() , .QN());
  DFF_X1 controller_roundCounter_Inst_Reg1_s_current_state_reg_1_ ( .D(
        controller_roundCounter_zero_or_PlusOne[1]), .CK(clk), .Q(
        controller_roundCounter_feedback1[1]) , .QN());
  XOR2_X1 prince_U196 ( .A(input_s1[0]), .B(prince_n267), .Z(
        prince_SR_Inv_Result_s1[16]) );
  XOR2_X1 prince_U195 ( .A(input_s1[10]), .B(prince_n266), .Z(
        prince_SR_Inv_Result_s1[58]) );
  XOR2_X1 prince_U194 ( .A(input_s1[11]), .B(prince_n265), .Z(
        prince_SR_Inv_Result_s1[59]) );
  XOR2_X1 prince_U193 ( .A(input_s1[12]), .B(prince_n264), .Z(
        prince_SR_Inv_Result_s1[12]) );
  XOR2_X1 prince_U192 ( .A(input_s1[13]), .B(prince_n263), .Z(
        prince_SR_Inv_Result_s1[13]) );
  XOR2_X1 prince_U191 ( .A(input_s1[14]), .B(prince_n262), .Z(
        prince_SR_Inv_Result_s1[14]) );
  XOR2_X1 prince_U190 ( .A(input_s1[15]), .B(prince_n261), .Z(
        prince_SR_Inv_Result_s1[15]) );
  XOR2_X1 prince_U189 ( .A(input_s1[16]), .B(prince_n260), .Z(
        prince_SR_Inv_Result_s1[32]) );
  XOR2_X1 prince_U188 ( .A(input_s1[17]), .B(prince_n259), .Z(
        prince_SR_Inv_Result_s1[33]) );
  XOR2_X1 prince_U187 ( .A(input_s1[18]), .B(prince_n258), .Z(
        prince_SR_Inv_Result_s1[34]) );
  XOR2_X1 prince_U186 ( .A(input_s1[19]), .B(prince_n257), .Z(
        prince_SR_Inv_Result_s1[35]) );
  XOR2_X1 prince_U185 ( .A(input_s1[1]), .B(prince_n256), .Z(
        prince_SR_Inv_Result_s1[17]) );
  XOR2_X1 prince_U184 ( .A(input_s1[20]), .B(prince_n255), .Z(
        prince_SR_Inv_Result_s1[52]) );
  XOR2_X1 prince_U183 ( .A(input_s1[21]), .B(prince_n254), .Z(
        prince_SR_Inv_Result_s1[53]) );
  XOR2_X1 prince_U182 ( .A(input_s1[22]), .B(prince_n253), .Z(
        prince_SR_Inv_Result_s1[54]) );
  XOR2_X1 prince_U181 ( .A(input_s1[23]), .B(prince_n252), .Z(
        prince_SR_Inv_Result_s1[55]) );
  XOR2_X1 prince_U180 ( .A(input_s1[24]), .B(prince_n251), .Z(
        prince_SR_Inv_Result_s1[8]) );
  XOR2_X1 prince_U179 ( .A(input_s1[25]), .B(prince_n250), .Z(
        prince_SR_Inv_Result_s1[9]) );
  XOR2_X1 prince_U178 ( .A(input_s1[26]), .B(prince_n249), .Z(
        prince_SR_Inv_Result_s1[10]) );
  XOR2_X1 prince_U177 ( .A(input_s1[27]), .B(prince_n248), .Z(
        prince_SR_Inv_Result_s1[11]) );
  XOR2_X1 prince_U176 ( .A(input_s1[28]), .B(prince_n247), .Z(
        prince_SR_Inv_Result_s1[28]) );
  XOR2_X1 prince_U175 ( .A(input_s1[29]), .B(prince_n246), .Z(
        prince_SR_Inv_Result_s1[29]) );
  XOR2_X1 prince_U174 ( .A(input_s1[2]), .B(prince_n245), .Z(
        prince_SR_Inv_Result_s1[18]) );
  XOR2_X1 prince_U173 ( .A(input_s1[30]), .B(prince_n244), .Z(
        prince_SR_Inv_Result_s1[30]) );
  XOR2_X1 prince_U172 ( .A(input_s1[31]), .B(prince_n243), .Z(
        prince_SR_Inv_Result_s1[31]) );
  XOR2_X1 prince_U171 ( .A(input_s1[32]), .B(prince_n242), .Z(
        prince_SR_Inv_Result_s1[48]) );
  XOR2_X1 prince_U170 ( .A(input_s1[33]), .B(prince_n241), .Z(
        prince_SR_Inv_Result_s1[49]) );
  XOR2_X1 prince_U169 ( .A(input_s1[34]), .B(prince_n240), .Z(
        prince_SR_Inv_Result_s1[50]) );
  XOR2_X1 prince_U168 ( .A(input_s1[35]), .B(prince_n239), .Z(
        prince_SR_Inv_Result_s1[51]) );
  XOR2_X1 prince_U167 ( .A(input_s1[36]), .B(prince_n238), .Z(
        prince_SR_Inv_Result_s1[4]) );
  XOR2_X1 prince_U166 ( .A(input_s1[37]), .B(prince_n237), .Z(
        prince_SR_Inv_Result_s1[5]) );
  XOR2_X1 prince_U165 ( .A(input_s1[38]), .B(prince_n236), .Z(
        prince_SR_Inv_Result_s1[6]) );
  XOR2_X1 prince_U164 ( .A(input_s1[39]), .B(prince_n235), .Z(
        prince_SR_Inv_Result_s1[7]) );
  XOR2_X1 prince_U163 ( .A(input_s1[3]), .B(prince_n234), .Z(
        prince_SR_Inv_Result_s1[19]) );
  XOR2_X1 prince_U162 ( .A(input_s1[40]), .B(prince_n233), .Z(
        prince_SR_Inv_Result_s1[24]) );
  XOR2_X1 prince_U161 ( .A(input_s1[41]), .B(prince_n232), .Z(
        prince_SR_Inv_Result_s1[25]) );
  XOR2_X1 prince_U160 ( .A(input_s1[42]), .B(prince_n231), .Z(
        prince_SR_Inv_Result_s1[26]) );
  XOR2_X1 prince_U159 ( .A(input_s1[43]), .B(prince_n230), .Z(
        prince_SR_Inv_Result_s1[27]) );
  XOR2_X1 prince_U158 ( .A(input_s1[44]), .B(prince_n229), .Z(
        prince_SR_Inv_Result_s1[44]) );
  XOR2_X1 prince_U157 ( .A(input_s1[45]), .B(prince_n228), .Z(
        prince_SR_Inv_Result_s1[45]) );
  XOR2_X1 prince_U156 ( .A(input_s1[46]), .B(prince_n227), .Z(
        prince_SR_Inv_Result_s1[46]) );
  XOR2_X1 prince_U155 ( .A(input_s1[47]), .B(prince_n226), .Z(
        prince_SR_Inv_Result_s1[47]) );
  XOR2_X1 prince_U154 ( .A(input_s1[48]), .B(prince_n225), .Z(
        prince_SR_Inv_Result_s1[0]) );
  XOR2_X1 prince_U153 ( .A(input_s1[49]), .B(prince_n224), .Z(
        prince_SR_Inv_Result_s1[1]) );
  XOR2_X1 prince_U152 ( .A(input_s1[4]), .B(prince_n223), .Z(
        prince_SR_Inv_Result_s1[36]) );
  XOR2_X1 prince_U151 ( .A(input_s1[50]), .B(prince_n222), .Z(
        prince_SR_Inv_Result_s1[2]) );
  XOR2_X1 prince_U150 ( .A(input_s1[51]), .B(prince_n221), .Z(
        prince_SR_Inv_Result_s1[3]) );
  XOR2_X1 prince_U149 ( .A(input_s1[52]), .B(prince_n220), .Z(
        prince_SR_Inv_Result_s1[20]) );
  XOR2_X1 prince_U148 ( .A(input_s1[53]), .B(prince_n219), .Z(
        prince_SR_Inv_Result_s1[21]) );
  XOR2_X1 prince_U147 ( .A(input_s1[54]), .B(prince_n218), .Z(
        prince_SR_Inv_Result_s1[22]) );
  XOR2_X1 prince_U146 ( .A(input_s1[55]), .B(prince_n217), .Z(
        prince_SR_Inv_Result_s1[23]) );
  XOR2_X1 prince_U145 ( .A(input_s1[56]), .B(prince_n216), .Z(
        prince_SR_Inv_Result_s1[40]) );
  XOR2_X1 prince_U144 ( .A(input_s1[57]), .B(prince_n215), .Z(
        prince_SR_Inv_Result_s1[41]) );
  XOR2_X1 prince_U143 ( .A(input_s1[58]), .B(prince_n214), .Z(
        prince_SR_Inv_Result_s1[42]) );
  XOR2_X1 prince_U142 ( .A(input_s1[59]), .B(prince_n213), .Z(
        prince_SR_Inv_Result_s1[43]) );
  XOR2_X1 prince_U141 ( .A(input_s1[5]), .B(prince_n212), .Z(
        prince_SR_Inv_Result_s1[37]) );
  XOR2_X1 prince_U140 ( .A(input_s1[60]), .B(prince_n211), .Z(
        prince_SR_Inv_Result_s1[60]) );
  XOR2_X1 prince_U139 ( .A(input_s1[61]), .B(prince_n210), .Z(
        prince_SR_Inv_Result_s1[61]) );
  XOR2_X1 prince_U138 ( .A(input_s1[62]), .B(prince_n209), .Z(
        prince_SR_Inv_Result_s1[62]) );
  XOR2_X1 prince_U137 ( .A(input_s1[63]), .B(prince_n208), .Z(
        prince_SR_Inv_Result_s1[63]) );
  XOR2_X1 prince_U136 ( .A(input_s1[6]), .B(prince_n207), .Z(
        prince_SR_Inv_Result_s1[38]) );
  XOR2_X1 prince_U135 ( .A(input_s1[7]), .B(prince_n206), .Z(
        prince_SR_Inv_Result_s1[39]) );
  XOR2_X1 prince_U134 ( .A(input_s1[8]), .B(prince_n205), .Z(
        prince_SR_Inv_Result_s1[56]) );
  XOR2_X1 prince_U133 ( .A(input_s1[9]), .B(prince_n204), .Z(
        prince_SR_Inv_Result_s1[57]) );
  XOR2_X1 prince_U132 ( .A(prince_rounds_SR_Inv_Result_s1[16]), .B(prince_n267), .Z(output_s1[0]) );
  MUX2_X1 prince_U131 ( .A(k_0_p_0_), .B(Key[64]), .S(prince_n203), .Z(
        prince_n267) );
  XOR2_X1 prince_U130 ( .A(prince_rounds_SR_Inv_Result_s1[58]), .B(prince_n266), .Z(output_s1[10]) );
  MUX2_X1 prince_U129 ( .A(Key[75]), .B(Key[74]), .S(prince_n203), .Z(
        prince_n266) );
  XOR2_X1 prince_U128 ( .A(prince_rounds_SR_Inv_Result_s1[59]), .B(prince_n265), .Z(output_s1[11]) );
  MUX2_X1 prince_U127 ( .A(Key[76]), .B(Key[75]), .S(prince_n203), .Z(
        prince_n265) );
  XOR2_X1 prince_U126 ( .A(prince_rounds_SR_Inv_Result_s1[12]), .B(prince_n264), .Z(output_s1[12]) );
  MUX2_X1 prince_U125 ( .A(Key[77]), .B(Key[76]), .S(prince_n203), .Z(
        prince_n264) );
  XOR2_X1 prince_U124 ( .A(prince_rounds_SR_Inv_Result_s1[13]), .B(prince_n263), .Z(output_s1[13]) );
  MUX2_X1 prince_U123 ( .A(Key[78]), .B(Key[77]), .S(prince_n202), .Z(
        prince_n263) );
  XOR2_X1 prince_U122 ( .A(prince_rounds_SR_Inv_Result_s1[14]), .B(prince_n262), .Z(output_s1[14]) );
  MUX2_X1 prince_U121 ( .A(Key[79]), .B(Key[78]), .S(prince_n202), .Z(
        prince_n262) );
  XOR2_X1 prince_U120 ( .A(prince_rounds_SR_Inv_Result_s1[15]), .B(prince_n261), .Z(output_s1[15]) );
  MUX2_X1 prince_U119 ( .A(Key[80]), .B(Key[79]), .S(prince_n202), .Z(
        prince_n261) );
  XOR2_X1 prince_U118 ( .A(prince_rounds_SR_Inv_Result_s1[32]), .B(prince_n260), .Z(output_s1[16]) );
  MUX2_X1 prince_U117 ( .A(Key[81]), .B(Key[80]), .S(prince_n202), .Z(
        prince_n260) );
  XOR2_X1 prince_U116 ( .A(prince_rounds_SR_Inv_Result_s1[33]), .B(prince_n259), .Z(output_s1[17]) );
  MUX2_X1 prince_U115 ( .A(Key[82]), .B(Key[81]), .S(prince_n202), .Z(
        prince_n259) );
  XOR2_X1 prince_U114 ( .A(prince_rounds_SR_Inv_Result_s1[34]), .B(prince_n258), .Z(output_s1[18]) );
  MUX2_X1 prince_U113 ( .A(Key[83]), .B(Key[82]), .S(prince_n202), .Z(
        prince_n258) );
  XOR2_X1 prince_U112 ( .A(prince_rounds_SR_Inv_Result_s1[35]), .B(prince_n257), .Z(output_s1[19]) );
  MUX2_X1 prince_U111 ( .A(Key[84]), .B(Key[83]), .S(prince_n202), .Z(
        prince_n257) );
  XOR2_X1 prince_U110 ( .A(prince_rounds_SR_Inv_Result_s1[17]), .B(prince_n256), .Z(output_s1[1]) );
  MUX2_X1 prince_U109 ( .A(Key[66]), .B(Key[65]), .S(prince_n202), .Z(
        prince_n256) );
  XOR2_X1 prince_U108 ( .A(prince_rounds_SR_Inv_Result_s1[52]), .B(prince_n255), .Z(output_s1[20]) );
  MUX2_X1 prince_U107 ( .A(Key[85]), .B(Key[84]), .S(prince_n202), .Z(
        prince_n255) );
  XOR2_X1 prince_U106 ( .A(prince_rounds_SR_Inv_Result_s1[53]), .B(prince_n254), .Z(output_s1[21]) );
  MUX2_X1 prince_U105 ( .A(Key[86]), .B(Key[85]), .S(prince_n202), .Z(
        prince_n254) );
  XOR2_X1 prince_U104 ( .A(prince_rounds_SR_Inv_Result_s1[54]), .B(prince_n253), .Z(output_s1[22]) );
  MUX2_X1 prince_U103 ( .A(Key[87]), .B(Key[86]), .S(prince_n202), .Z(
        prince_n253) );
  XOR2_X1 prince_U102 ( .A(prince_rounds_SR_Inv_Result_s1[55]), .B(prince_n252), .Z(output_s1[23]) );
  MUX2_X1 prince_U101 ( .A(Key[88]), .B(Key[87]), .S(prince_n202), .Z(
        prince_n252) );
  XOR2_X1 prince_U100 ( .A(prince_rounds_SR_Inv_Result_s1[8]), .B(prince_n251), 
        .Z(output_s1[24]) );
  MUX2_X1 prince_U99 ( .A(Key[89]), .B(Key[88]), .S(prince_n202), .Z(
        prince_n251) );
  XOR2_X1 prince_U98 ( .A(prince_rounds_SR_Inv_Result_s1[9]), .B(prince_n250), 
        .Z(output_s1[25]) );
  MUX2_X1 prince_U97 ( .A(Key[90]), .B(Key[89]), .S(prince_n201), .Z(
        prince_n250) );
  XOR2_X1 prince_U96 ( .A(prince_rounds_SR_Inv_Result_s1[10]), .B(prince_n249), 
        .Z(output_s1[26]) );
  MUX2_X1 prince_U95 ( .A(Key[91]), .B(Key[90]), .S(prince_n202), .Z(
        prince_n249) );
  XOR2_X1 prince_U94 ( .A(prince_rounds_SR_Inv_Result_s1[11]), .B(prince_n248), 
        .Z(output_s1[27]) );
  MUX2_X1 prince_U93 ( .A(Key[92]), .B(Key[91]), .S(prince_n203), .Z(
        prince_n248) );
  XOR2_X1 prince_U92 ( .A(prince_rounds_SR_Inv_Result_s1[28]), .B(prince_n247), 
        .Z(output_s1[28]) );
  MUX2_X1 prince_U91 ( .A(Key[93]), .B(Key[92]), .S(prince_n201), .Z(
        prince_n247) );
  XOR2_X1 prince_U90 ( .A(prince_rounds_SR_Inv_Result_s1[29]), .B(prince_n246), 
        .Z(output_s1[29]) );
  MUX2_X1 prince_U89 ( .A(Key[94]), .B(Key[93]), .S(prince_n202), .Z(
        prince_n246) );
  XOR2_X1 prince_U88 ( .A(prince_rounds_SR_Inv_Result_s1[18]), .B(prince_n245), 
        .Z(output_s1[2]) );
  MUX2_X1 prince_U87 ( .A(Key[67]), .B(Key[66]), .S(prince_n203), .Z(
        prince_n245) );
  XOR2_X1 prince_U86 ( .A(prince_rounds_SR_Inv_Result_s1[30]), .B(prince_n244), 
        .Z(output_s1[30]) );
  MUX2_X1 prince_U85 ( .A(Key[95]), .B(Key[94]), .S(prince_n201), .Z(
        prince_n244) );
  XOR2_X1 prince_U84 ( .A(prince_rounds_SR_Inv_Result_s1[31]), .B(prince_n243), 
        .Z(output_s1[31]) );
  MUX2_X1 prince_U83 ( .A(Key[96]), .B(Key[95]), .S(prince_n201), .Z(
        prince_n243) );
  XOR2_X1 prince_U82 ( .A(prince_rounds_SR_Inv_Result_s1[48]), .B(prince_n242), 
        .Z(output_s1[32]) );
  MUX2_X1 prince_U81 ( .A(Key[97]), .B(Key[96]), .S(prince_n201), .Z(
        prince_n242) );
  XOR2_X1 prince_U80 ( .A(prince_rounds_SR_Inv_Result_s1[49]), .B(prince_n241), 
        .Z(output_s1[33]) );
  MUX2_X1 prince_U79 ( .A(Key[98]), .B(Key[97]), .S(prince_n201), .Z(
        prince_n241) );
  XOR2_X1 prince_U78 ( .A(prince_rounds_SR_Inv_Result_s1[50]), .B(prince_n240), 
        .Z(output_s1[34]) );
  MUX2_X1 prince_U77 ( .A(Key[99]), .B(Key[98]), .S(prince_n201), .Z(
        prince_n240) );
  XOR2_X1 prince_U76 ( .A(prince_rounds_SR_Inv_Result_s1[51]), .B(prince_n239), 
        .Z(output_s1[35]) );
  MUX2_X1 prince_U75 ( .A(Key[100]), .B(Key[99]), .S(prince_n203), .Z(
        prince_n239) );
  XOR2_X1 prince_U74 ( .A(prince_rounds_SR_Inv_Result_s1[4]), .B(prince_n238), 
        .Z(output_s1[36]) );
  MUX2_X1 prince_U73 ( .A(Key[101]), .B(Key[100]), .S(prince_n203), .Z(
        prince_n238) );
  XOR2_X1 prince_U72 ( .A(prince_rounds_SR_Inv_Result_s1[5]), .B(prince_n237), 
        .Z(output_s1[37]) );
  MUX2_X1 prince_U71 ( .A(Key[102]), .B(Key[101]), .S(prince_n203), .Z(
        prince_n237) );
  XOR2_X1 prince_U70 ( .A(prince_rounds_SR_Inv_Result_s1[6]), .B(prince_n236), 
        .Z(output_s1[38]) );
  MUX2_X1 prince_U69 ( .A(Key[103]), .B(Key[102]), .S(prince_n203), .Z(
        prince_n236) );
  XOR2_X1 prince_U68 ( .A(prince_rounds_SR_Inv_Result_s1[7]), .B(prince_n235), 
        .Z(output_s1[39]) );
  MUX2_X1 prince_U67 ( .A(Key[104]), .B(Key[103]), .S(prince_n203), .Z(
        prince_n235) );
  XOR2_X1 prince_U66 ( .A(prince_rounds_SR_Inv_Result_s1[19]), .B(prince_n234), 
        .Z(output_s1[3]) );
  MUX2_X1 prince_U65 ( .A(Key[68]), .B(Key[67]), .S(prince_n203), .Z(
        prince_n234) );
  XOR2_X1 prince_U64 ( .A(prince_rounds_SR_Inv_Result_s1[24]), .B(prince_n233), 
        .Z(output_s1[40]) );
  MUX2_X1 prince_U63 ( .A(Key[105]), .B(Key[104]), .S(prince_n203), .Z(
        prince_n233) );
  XOR2_X1 prince_U62 ( .A(prince_rounds_SR_Inv_Result_s1[25]), .B(prince_n232), 
        .Z(output_s1[41]) );
  MUX2_X1 prince_U61 ( .A(Key[106]), .B(Key[105]), .S(prince_n203), .Z(
        prince_n232) );
  XOR2_X1 prince_U60 ( .A(prince_rounds_SR_Inv_Result_s1[26]), .B(prince_n231), 
        .Z(output_s1[42]) );
  MUX2_X1 prince_U59 ( .A(Key[107]), .B(Key[106]), .S(prince_n203), .Z(
        prince_n231) );
  XOR2_X1 prince_U58 ( .A(prince_rounds_SR_Inv_Result_s1[27]), .B(prince_n230), 
        .Z(output_s1[43]) );
  MUX2_X1 prince_U57 ( .A(Key[108]), .B(Key[107]), .S(prince_n202), .Z(
        prince_n230) );
  XOR2_X1 prince_U56 ( .A(prince_rounds_SR_Inv_Result_s1[44]), .B(prince_n229), 
        .Z(output_s1[44]) );
  MUX2_X1 prince_U55 ( .A(Key[109]), .B(Key[108]), .S(prince_n202), .Z(
        prince_n229) );
  XOR2_X1 prince_U54 ( .A(prince_rounds_SR_Inv_Result_s1[45]), .B(prince_n228), 
        .Z(output_s1[45]) );
  MUX2_X1 prince_U53 ( .A(Key[110]), .B(Key[109]), .S(prince_n201), .Z(
        prince_n228) );
  XOR2_X1 prince_U52 ( .A(prince_rounds_SR_Inv_Result_s1[46]), .B(prince_n227), 
        .Z(output_s1[46]) );
  MUX2_X1 prince_U51 ( .A(Key[111]), .B(Key[110]), .S(prince_n203), .Z(
        prince_n227) );
  XOR2_X1 prince_U50 ( .A(prince_rounds_SR_Inv_Result_s1[47]), .B(prince_n226), 
        .Z(output_s1[47]) );
  MUX2_X1 prince_U49 ( .A(Key[112]), .B(Key[111]), .S(prince_n202), .Z(
        prince_n226) );
  XOR2_X1 prince_U48 ( .A(prince_rounds_SR_Inv_Result_s1[0]), .B(prince_n225), 
        .Z(output_s1[48]) );
  MUX2_X1 prince_U47 ( .A(Key[113]), .B(Key[112]), .S(prince_n203), .Z(
        prince_n225) );
  XOR2_X1 prince_U46 ( .A(prince_rounds_SR_Inv_Result_s1[1]), .B(prince_n224), 
        .Z(output_s1[49]) );
  MUX2_X1 prince_U45 ( .A(Key[114]), .B(Key[113]), .S(prince_n201), .Z(
        prince_n224) );
  XOR2_X1 prince_U44 ( .A(prince_rounds_SR_Inv_Result_s1[36]), .B(prince_n223), 
        .Z(output_s1[4]) );
  MUX2_X1 prince_U43 ( .A(Key[69]), .B(Key[68]), .S(prince_n203), .Z(
        prince_n223) );
  XOR2_X1 prince_U42 ( .A(prince_rounds_SR_Inv_Result_s1[2]), .B(prince_n222), 
        .Z(output_s1[50]) );
  MUX2_X1 prince_U41 ( .A(Key[115]), .B(Key[114]), .S(prince_n202), .Z(
        prince_n222) );
  XOR2_X1 prince_U40 ( .A(prince_rounds_SR_Inv_Result_s1[3]), .B(prince_n221), 
        .Z(output_s1[51]) );
  MUX2_X1 prince_U39 ( .A(Key[116]), .B(Key[115]), .S(prince_n201), .Z(
        prince_n221) );
  XOR2_X1 prince_U38 ( .A(prince_rounds_SR_Inv_Result_s1[20]), .B(prince_n220), 
        .Z(output_s1[52]) );
  MUX2_X1 prince_U37 ( .A(Key[117]), .B(Key[116]), .S(prince_n201), .Z(
        prince_n220) );
  XOR2_X1 prince_U36 ( .A(prince_rounds_SR_Inv_Result_s1[21]), .B(prince_n219), 
        .Z(output_s1[53]) );
  MUX2_X1 prince_U35 ( .A(Key[118]), .B(Key[117]), .S(prince_n203), .Z(
        prince_n219) );
  XOR2_X1 prince_U34 ( .A(prince_rounds_SR_Inv_Result_s1[22]), .B(prince_n218), 
        .Z(output_s1[54]) );
  MUX2_X1 prince_U33 ( .A(Key[119]), .B(Key[118]), .S(prince_n202), .Z(
        prince_n218) );
  INV_X1 prince_U32 ( .A(prince_n200), .ZN(prince_n202) );
  XOR2_X1 prince_U31 ( .A(prince_rounds_SR_Inv_Result_s1[23]), .B(prince_n217), 
        .Z(output_s1[55]) );
  MUX2_X1 prince_U30 ( .A(Key[120]), .B(Key[119]), .S(prince_n203), .Z(
        prince_n217) );
  INV_X1 prince_U29 ( .A(prince_n200), .ZN(prince_n203) );
  XOR2_X1 prince_U28 ( .A(prince_rounds_SR_Inv_Result_s1[40]), .B(prince_n216), 
        .Z(output_s1[56]) );
  MUX2_X1 prince_U27 ( .A(Key[121]), .B(Key[120]), .S(prince_n201), .Z(
        prince_n216) );
  XOR2_X1 prince_U26 ( .A(prince_rounds_SR_Inv_Result_s1[41]), .B(prince_n215), 
        .Z(output_s1[57]) );
  MUX2_X1 prince_U25 ( .A(Key[122]), .B(Key[121]), .S(prince_n201), .Z(
        prince_n215) );
  XOR2_X1 prince_U24 ( .A(prince_rounds_SR_Inv_Result_s1[42]), .B(prince_n214), 
        .Z(output_s1[58]) );
  MUX2_X1 prince_U23 ( .A(Key[123]), .B(Key[122]), .S(prince_n201), .Z(
        prince_n214) );
  XOR2_X1 prince_U22 ( .A(prince_rounds_SR_Inv_Result_s1[43]), .B(prince_n213), 
        .Z(output_s1[59]) );
  MUX2_X1 prince_U21 ( .A(Key[124]), .B(Key[123]), .S(prince_n201), .Z(
        prince_n213) );
  XOR2_X1 prince_U20 ( .A(prince_rounds_SR_Inv_Result_s1[37]), .B(prince_n212), 
        .Z(output_s1[5]) );
  MUX2_X1 prince_U19 ( .A(Key[70]), .B(Key[69]), .S(prince_n201), .Z(
        prince_n212) );
  XOR2_X1 prince_U18 ( .A(prince_rounds_SR_Inv_Result_s1[60]), .B(prince_n211), 
        .Z(output_s1[60]) );
  MUX2_X1 prince_U17 ( .A(Key[125]), .B(Key[124]), .S(prince_n201), .Z(
        prince_n211) );
  XOR2_X1 prince_U16 ( .A(prince_rounds_SR_Inv_Result_s1[61]), .B(prince_n210), 
        .Z(output_s1[61]) );
  MUX2_X1 prince_U15 ( .A(Key[126]), .B(Key[125]), .S(prince_n201), .Z(
        prince_n210) );
  XOR2_X1 prince_U14 ( .A(prince_rounds_SR_Inv_Result_s1[62]), .B(prince_n209), 
        .Z(output_s1[62]) );
  MUX2_X1 prince_U13 ( .A(Key[127]), .B(Key[126]), .S(prince_n201), .Z(
        prince_n209) );
  XOR2_X1 prince_U12 ( .A(prince_rounds_SR_Inv_Result_s1[63]), .B(prince_n208), 
        .Z(output_s1[63]) );
  MUX2_X1 prince_U11 ( .A(Key[64]), .B(Key[127]), .S(prince_n201), .Z(
        prince_n208) );
  XOR2_X1 prince_U10 ( .A(prince_rounds_SR_Inv_Result_s1[38]), .B(prince_n207), 
        .Z(output_s1[6]) );
  MUX2_X1 prince_U9 ( .A(Key[71]), .B(Key[70]), .S(prince_n201), .Z(
        prince_n207) );
  XOR2_X1 prince_U8 ( .A(prince_rounds_SR_Inv_Result_s1[39]), .B(prince_n206), 
        .Z(output_s1[7]) );
  MUX2_X1 prince_U7 ( .A(Key[72]), .B(Key[71]), .S(prince_n201), .Z(
        prince_n206) );
  XOR2_X1 prince_U6 ( .A(prince_rounds_SR_Inv_Result_s1[56]), .B(prince_n205), 
        .Z(output_s1[8]) );
  MUX2_X1 prince_U5 ( .A(Key[73]), .B(Key[72]), .S(prince_n201), .Z(
        prince_n205) );
  XOR2_X1 prince_U4 ( .A(prince_rounds_SR_Inv_Result_s1[57]), .B(prince_n204), 
        .Z(output_s1[9]) );
  MUX2_X1 prince_U3 ( .A(Key[74]), .B(Key[73]), .S(prince_n201), .Z(
        prince_n204) );
  XNOR2_X1 prince_U2 ( .A(enc_dec), .B(rst), .ZN(prince_n200) );
  INV_X2 prince_U1 ( .A(prince_n200), .ZN(prince_n201) );
  XNOR2_X1 prince_rounds_U327 ( .A(prince_rounds_sub_Inv_Result_s1[63]), .B(
        prince_rounds_n402), .ZN(prince_rounds_SR_Inv_Result_s1[63]) );
  XNOR2_X1 prince_rounds_U326 ( .A(prince_rounds_SR_Result_s1[63]), .B(
        prince_rounds_n402), .ZN(prince_rounds_round_inputXORkeyRCON_s1[63])
         );
  XNOR2_X1 prince_rounds_U325 ( .A(Key[63]), .B(
        prince_rounds_round_Constant[63]), .ZN(prince_rounds_n402) );
  XNOR2_X1 prince_rounds_U324 ( .A(prince_rounds_sub_Inv_Result_s1[1]), .B(
        prince_rounds_n401), .ZN(prince_rounds_SR_Inv_Result_s1[17]) );
  XNOR2_X1 prince_rounds_U323 ( .A(prince_rounds_SR_Result_s1[1]), .B(
        prince_rounds_n401), .ZN(prince_rounds_round_inputXORkeyRCON_s1[1]) );
  XNOR2_X1 prince_rounds_U322 ( .A(Key[1]), .B(prince_rounds_round_Constant[1]), .ZN(prince_rounds_n401) );
  XNOR2_X1 prince_rounds_U321 ( .A(prince_rounds_sub_Inv_Result_s1[62]), .B(
        prince_rounds_n400), .ZN(prince_rounds_SR_Inv_Result_s1[62]) );
  XNOR2_X1 prince_rounds_U320 ( .A(prince_rounds_SR_Result_s1[62]), .B(
        prince_rounds_n400), .ZN(prince_rounds_round_inputXORkeyRCON_s1[62])
         );
  XNOR2_X1 prince_rounds_U319 ( .A(Key[62]), .B(
        prince_rounds_round_Constant[62]), .ZN(prince_rounds_n400) );
  XNOR2_X1 prince_rounds_U318 ( .A(prince_rounds_sub_Inv_Result_s1[60]), .B(
        prince_rounds_n399), .ZN(prince_rounds_SR_Inv_Result_s1[60]) );
  XNOR2_X1 prince_rounds_U317 ( .A(prince_rounds_SR_Result_s1[60]), .B(
        prince_rounds_n399), .ZN(prince_rounds_round_inputXORkeyRCON_s1[60])
         );
  XNOR2_X1 prince_rounds_U316 ( .A(Key[60]), .B(
        prince_rounds_round_Constant[60]), .ZN(prince_rounds_n399) );
  XNOR2_X1 prince_rounds_U315 ( .A(prince_rounds_sub_Inv_Result_s1[56]), .B(
        prince_rounds_n398), .ZN(prince_rounds_SR_Inv_Result_s1[40]) );
  XNOR2_X1 prince_rounds_U314 ( .A(prince_rounds_SR_Result_s1[56]), .B(
        prince_rounds_n398), .ZN(prince_rounds_round_inputXORkeyRCON_s1[56])
         );
  XNOR2_X1 prince_rounds_U313 ( .A(Key[56]), .B(
        prince_rounds_round_Constant[56]), .ZN(prince_rounds_n398) );
  XNOR2_X1 prince_rounds_U312 ( .A(prince_rounds_sub_Inv_Result_s1[48]), .B(
        prince_rounds_n397), .ZN(prince_rounds_SR_Inv_Result_s1[0]) );
  XNOR2_X1 prince_rounds_U311 ( .A(prince_rounds_SR_Result_s1[48]), .B(
        prince_rounds_n397), .ZN(prince_rounds_round_inputXORkeyRCON_s1[48])
         );
  XNOR2_X1 prince_rounds_U310 ( .A(Key[48]), .B(
        prince_rounds_round_Constant[48]), .ZN(prince_rounds_n397) );
  XNOR2_X1 prince_rounds_U309 ( .A(prince_rounds_sub_Inv_Result_s1[32]), .B(
        prince_rounds_n396), .ZN(prince_rounds_SR_Inv_Result_s1[48]) );
  XNOR2_X1 prince_rounds_U308 ( .A(prince_rounds_SR_Result_s1[32]), .B(
        prince_rounds_n396), .ZN(prince_rounds_round_inputXORkeyRCON_s1[32])
         );
  XNOR2_X1 prince_rounds_U307 ( .A(Key[32]), .B(
        prince_rounds_round_Constant[32]), .ZN(prince_rounds_n396) );
  XNOR2_X1 prince_rounds_U306 ( .A(prince_rounds_sub_Inv_Result_s1[31]), .B(
        prince_rounds_n395), .ZN(prince_rounds_SR_Inv_Result_s1[31]) );
  XNOR2_X1 prince_rounds_U305 ( .A(prince_rounds_SR_Result_s1[31]), .B(
        prince_rounds_n395), .ZN(prince_rounds_round_inputXORkeyRCON_s1[31])
         );
  XNOR2_X1 prince_rounds_U304 ( .A(Key[31]), .B(
        prince_rounds_round_Constant[36]), .ZN(prince_rounds_n395) );
  XNOR2_X1 prince_rounds_U303 ( .A(prince_rounds_sub_Inv_Result_s1[47]), .B(
        prince_rounds_n394), .ZN(prince_rounds_SR_Inv_Result_s1[47]) );
  XNOR2_X1 prince_rounds_U302 ( .A(prince_rounds_SR_Result_s1[47]), .B(
        prince_rounds_n394), .ZN(prince_rounds_round_inputXORkeyRCON_s1[47])
         );
  XNOR2_X1 prince_rounds_U301 ( .A(Key[47]), .B(
        prince_rounds_round_Constant[47]), .ZN(prince_rounds_n394) );
  XNOR2_X1 prince_rounds_U300 ( .A(prince_rounds_sub_Inv_Result_s1[30]), .B(
        prince_rounds_n393), .ZN(prince_rounds_SR_Inv_Result_s1[30]) );
  XNOR2_X1 prince_rounds_U299 ( .A(prince_rounds_SR_Result_s1[30]), .B(
        prince_rounds_n393), .ZN(prince_rounds_round_inputXORkeyRCON_s1[30])
         );
  XNOR2_X1 prince_rounds_U298 ( .A(Key[30]), .B(
        prince_rounds_round_Constant[36]), .ZN(prince_rounds_n393) );
  XNOR2_X1 prince_rounds_U297 ( .A(prince_rounds_sub_Inv_Result_s1[29]), .B(
        prince_rounds_n392), .ZN(prince_rounds_SR_Inv_Result_s1[29]) );
  XNOR2_X1 prince_rounds_U296 ( .A(prince_rounds_SR_Result_s1[29]), .B(
        prince_rounds_n392), .ZN(prince_rounds_round_inputXORkeyRCON_s1[29])
         );
  XNOR2_X1 prince_rounds_U295 ( .A(Key[29]), .B(
        prince_rounds_round_Constant[29]), .ZN(prince_rounds_n392) );
  XNOR2_X1 prince_rounds_U294 ( .A(prince_rounds_sub_Inv_Result_s1[55]), .B(
        prince_rounds_n391), .ZN(prince_rounds_SR_Inv_Result_s1[23]) );
  XNOR2_X1 prince_rounds_U293 ( .A(prince_rounds_SR_Result_s1[55]), .B(
        prince_rounds_n391), .ZN(prince_rounds_round_inputXORkeyRCON_s1[55])
         );
  XNOR2_X1 prince_rounds_U292 ( .A(Key[55]), .B(
        prince_rounds_round_Constant[55]), .ZN(prince_rounds_n391) );
  XNOR2_X1 prince_rounds_U291 ( .A(prince_rounds_sub_Inv_Result_s1[46]), .B(
        prince_rounds_n390), .ZN(prince_rounds_SR_Inv_Result_s1[46]) );
  XNOR2_X1 prince_rounds_U290 ( .A(prince_rounds_SR_Result_s1[46]), .B(
        prince_rounds_n390), .ZN(prince_rounds_round_inputXORkeyRCON_s1[46])
         );
  XNOR2_X1 prince_rounds_U289 ( .A(Key[46]), .B(
        prince_rounds_round_Constant[59]), .ZN(prince_rounds_n390) );
  XNOR2_X1 prince_rounds_U288 ( .A(prince_rounds_sub_Inv_Result_s1[28]), .B(
        prince_rounds_n389), .ZN(prince_rounds_SR_Inv_Result_s1[28]) );
  XNOR2_X1 prince_rounds_U287 ( .A(prince_rounds_SR_Result_s1[28]), .B(
        prince_rounds_n389), .ZN(prince_rounds_round_inputXORkeyRCON_s1[28])
         );
  XNOR2_X1 prince_rounds_U286 ( .A(Key[28]), .B(
        prince_rounds_round_Constant[38]), .ZN(prince_rounds_n389) );
  XNOR2_X1 prince_rounds_U285 ( .A(prince_rounds_sub_Inv_Result_s1[27]), .B(
        prince_rounds_n388), .ZN(prince_rounds_SR_Inv_Result_s1[11]) );
  XNOR2_X1 prince_rounds_U284 ( .A(prince_rounds_SR_Result_s1[27]), .B(
        prince_rounds_n388), .ZN(prince_rounds_round_inputXORkeyRCON_s1[27])
         );
  XNOR2_X1 prince_rounds_U283 ( .A(Key[27]), .B(
        prince_rounds_round_Constant[27]), .ZN(prince_rounds_n388) );
  XNOR2_X1 prince_rounds_U282 ( .A(prince_rounds_sub_Inv_Result_s1[45]), .B(
        prince_rounds_n387), .ZN(prince_rounds_SR_Inv_Result_s1[45]) );
  XNOR2_X1 prince_rounds_U281 ( .A(prince_rounds_SR_Result_s1[45]), .B(
        prince_rounds_n387), .ZN(prince_rounds_round_inputXORkeyRCON_s1[45])
         );
  XNOR2_X1 prince_rounds_U280 ( .A(Key[45]), .B(
        prince_rounds_round_Constant[45]), .ZN(prince_rounds_n387) );
  XNOR2_X1 prince_rounds_U279 ( .A(prince_rounds_sub_Inv_Result_s1[26]), .B(
        prince_rounds_n386), .ZN(prince_rounds_SR_Inv_Result_s1[10]) );
  XNOR2_X1 prince_rounds_U278 ( .A(prince_rounds_SR_Result_s1[26]), .B(
        prince_rounds_n386), .ZN(prince_rounds_round_inputXORkeyRCON_s1[26])
         );
  XNOR2_X1 prince_rounds_U277 ( .A(Key[26]), .B(
        prince_rounds_round_Constant[59]), .ZN(prince_rounds_n386) );
  XNOR2_X1 prince_rounds_U276 ( .A(prince_rounds_sub_Inv_Result_s1[25]), .B(
        prince_rounds_n385), .ZN(prince_rounds_SR_Inv_Result_s1[9]) );
  XNOR2_X1 prince_rounds_U275 ( .A(prince_rounds_SR_Result_s1[25]), .B(
        prince_rounds_n385), .ZN(prince_rounds_round_inputXORkeyRCON_s1[25])
         );
  XNOR2_X1 prince_rounds_U274 ( .A(Key[25]), .B(
        prince_rounds_round_Constant[25]), .ZN(prince_rounds_n385) );
  XNOR2_X1 prince_rounds_U273 ( .A(prince_rounds_sub_Inv_Result_s1[59]), .B(
        prince_rounds_n384), .ZN(prince_rounds_SR_Inv_Result_s1[43]) );
  XNOR2_X1 prince_rounds_U272 ( .A(prince_rounds_SR_Result_s1[59]), .B(
        prince_rounds_n384), .ZN(prince_rounds_round_inputXORkeyRCON_s1[59])
         );
  XNOR2_X1 prince_rounds_U271 ( .A(Key[59]), .B(
        prince_rounds_round_Constant[59]), .ZN(prince_rounds_n384) );
  XNOR2_X1 prince_rounds_U270 ( .A(prince_rounds_sub_Inv_Result_s1[54]), .B(
        prince_rounds_n383), .ZN(prince_rounds_SR_Inv_Result_s1[22]) );
  XNOR2_X1 prince_rounds_U269 ( .A(prince_rounds_SR_Result_s1[54]), .B(
        prince_rounds_n383), .ZN(prince_rounds_round_inputXORkeyRCON_s1[54])
         );
  XNOR2_X1 prince_rounds_U268 ( .A(Key[54]), .B(
        prince_rounds_round_Constant[54]), .ZN(prince_rounds_n383) );
  XNOR2_X1 prince_rounds_U267 ( .A(prince_rounds_sub_Inv_Result_s1[44]), .B(
        prince_rounds_n382), .ZN(prince_rounds_SR_Inv_Result_s1[44]) );
  XNOR2_X1 prince_rounds_U266 ( .A(prince_rounds_SR_Result_s1[44]), .B(
        prince_rounds_n382), .ZN(prince_rounds_round_inputXORkeyRCON_s1[44])
         );
  XNOR2_X1 prince_rounds_U265 ( .A(Key[44]), .B(
        prince_rounds_round_Constant[44]), .ZN(prince_rounds_n382) );
  XNOR2_X1 prince_rounds_U264 ( .A(prince_rounds_sub_Inv_Result_s1[24]), .B(
        prince_rounds_n381), .ZN(prince_rounds_SR_Inv_Result_s1[8]) );
  XNOR2_X1 prince_rounds_U263 ( .A(prince_rounds_SR_Result_s1[24]), .B(
        prince_rounds_n381), .ZN(prince_rounds_round_inputXORkeyRCON_s1[24])
         );
  XNOR2_X1 prince_rounds_U262 ( .A(Key[24]), .B(
        prince_rounds_round_Constant[24]), .ZN(prince_rounds_n381) );
  XNOR2_X1 prince_rounds_U261 ( .A(prince_rounds_sub_Inv_Result_s1[23]), .B(
        prince_rounds_n380), .ZN(prince_rounds_SR_Inv_Result_s1[55]) );
  XNOR2_X1 prince_rounds_U260 ( .A(prince_rounds_SR_Result_s1[23]), .B(
        prince_rounds_n380), .ZN(prince_rounds_round_inputXORkeyRCON_s1[23])
         );
  XNOR2_X1 prince_rounds_U259 ( .A(Key[23]), .B(
        prince_rounds_round_Constant[58]), .ZN(prince_rounds_n380) );
  XNOR2_X1 prince_rounds_U258 ( .A(prince_rounds_sub_Inv_Result_s1[43]), .B(
        prince_rounds_n379), .ZN(prince_rounds_SR_Inv_Result_s1[27]) );
  XNOR2_X1 prince_rounds_U257 ( .A(prince_rounds_SR_Result_s1[43]), .B(
        prince_rounds_n379), .ZN(prince_rounds_round_inputXORkeyRCON_s1[43])
         );
  XNOR2_X1 prince_rounds_U256 ( .A(Key[43]), .B(
        prince_rounds_round_Constant[43]), .ZN(prince_rounds_n379) );
  XNOR2_X1 prince_rounds_U255 ( .A(prince_rounds_sub_Inv_Result_s1[22]), .B(
        prince_rounds_n378), .ZN(prince_rounds_SR_Inv_Result_s1[54]) );
  XNOR2_X1 prince_rounds_U254 ( .A(prince_rounds_SR_Result_s1[22]), .B(
        prince_rounds_n378), .ZN(prince_rounds_round_inputXORkeyRCON_s1[22])
         );
  XNOR2_X1 prince_rounds_U253 ( .A(Key[22]), .B(
        prince_rounds_round_Constant[22]), .ZN(prince_rounds_n378) );
  XNOR2_X1 prince_rounds_U252 ( .A(prince_rounds_sub_Inv_Result_s1[21]), .B(
        prince_rounds_n377), .ZN(prince_rounds_SR_Inv_Result_s1[53]) );
  XNOR2_X1 prince_rounds_U251 ( .A(prince_rounds_SR_Result_s1[21]), .B(
        prince_rounds_n377), .ZN(prince_rounds_round_inputXORkeyRCON_s1[21])
         );
  XNOR2_X1 prince_rounds_U250 ( .A(Key[21]), .B(
        prince_rounds_round_Constant[21]), .ZN(prince_rounds_n377) );
  XNOR2_X1 prince_rounds_U249 ( .A(prince_rounds_sub_Inv_Result_s1[53]), .B(
        prince_rounds_n376), .ZN(prince_rounds_SR_Inv_Result_s1[21]) );
  XNOR2_X1 prince_rounds_U248 ( .A(prince_rounds_SR_Result_s1[53]), .B(
        prince_rounds_n376), .ZN(prince_rounds_round_inputXORkeyRCON_s1[53])
         );
  XNOR2_X1 prince_rounds_U247 ( .A(Key[53]), .B(
        prince_rounds_round_Constant[53]), .ZN(prince_rounds_n376) );
  XNOR2_X1 prince_rounds_U246 ( .A(prince_rounds_sub_Inv_Result_s1[42]), .B(
        prince_rounds_n375), .ZN(prince_rounds_SR_Inv_Result_s1[26]) );
  XNOR2_X1 prince_rounds_U245 ( .A(prince_rounds_SR_Result_s1[42]), .B(
        prince_rounds_n375), .ZN(prince_rounds_round_inputXORkeyRCON_s1[42])
         );
  XNOR2_X1 prince_rounds_U244 ( .A(Key[42]), .B(
        prince_rounds_round_Constant[54]), .ZN(prince_rounds_n375) );
  XNOR2_X1 prince_rounds_U243 ( .A(prince_rounds_sub_Inv_Result_s1[20]), .B(
        prince_rounds_n374), .ZN(prince_rounds_SR_Inv_Result_s1[52]) );
  XNOR2_X1 prince_rounds_U242 ( .A(prince_rounds_SR_Result_s1[20]), .B(
        prince_rounds_n374), .ZN(prince_rounds_round_inputXORkeyRCON_s1[20])
         );
  XNOR2_X1 prince_rounds_U241 ( .A(Key[20]), .B(
        prince_rounds_round_Constant[37]), .ZN(prince_rounds_n374) );
  XNOR2_X1 prince_rounds_U240 ( .A(prince_rounds_sub_Inv_Result_s1[19]), .B(
        prince_rounds_n373), .ZN(prince_rounds_SR_Inv_Result_s1[35]) );
  XNOR2_X1 prince_rounds_U239 ( .A(prince_rounds_SR_Result_s1[19]), .B(
        prince_rounds_n373), .ZN(prince_rounds_round_inputXORkeyRCON_s1[19])
         );
  XNOR2_X1 prince_rounds_U238 ( .A(Key[19]), .B(
        prince_rounds_round_Constant[19]), .ZN(prince_rounds_n373) );
  XNOR2_X1 prince_rounds_U237 ( .A(prince_rounds_sub_Inv_Result_s1[41]), .B(
        prince_rounds_n372), .ZN(prince_rounds_SR_Inv_Result_s1[25]) );
  XNOR2_X1 prince_rounds_U236 ( .A(prince_rounds_SR_Result_s1[41]), .B(
        prince_rounds_n372), .ZN(prince_rounds_round_inputXORkeyRCON_s1[41])
         );
  XNOR2_X1 prince_rounds_U235 ( .A(Key[41]), .B(
        prince_rounds_round_Constant[41]), .ZN(prince_rounds_n372) );
  XNOR2_X1 prince_rounds_U234 ( .A(prince_rounds_sub_Inv_Result_s1[18]), .B(
        prince_rounds_n371), .ZN(prince_rounds_SR_Inv_Result_s1[34]) );
  XNOR2_X1 prince_rounds_U233 ( .A(prince_rounds_SR_Result_s1[18]), .B(
        prince_rounds_n371), .ZN(prince_rounds_round_inputXORkeyRCON_s1[18])
         );
  XNOR2_X1 prince_rounds_U232 ( .A(Key[18]), .B(
        prince_rounds_round_Constant[18]), .ZN(prince_rounds_n371) );
  XNOR2_X1 prince_rounds_U231 ( .A(prince_rounds_sub_Inv_Result_s1[17]), .B(
        prince_rounds_n370), .ZN(prince_rounds_SR_Inv_Result_s1[33]) );
  XNOR2_X1 prince_rounds_U230 ( .A(prince_rounds_SR_Result_s1[17]), .B(
        prince_rounds_n370), .ZN(prince_rounds_round_inputXORkeyRCON_s1[17])
         );
  XNOR2_X1 prince_rounds_U229 ( .A(Key[17]), .B(
        prince_rounds_round_Constant[44]), .ZN(prince_rounds_n370) );
  XNOR2_X1 prince_rounds_U228 ( .A(prince_rounds_sub_Inv_Result_s1[61]), .B(
        prince_rounds_n369), .ZN(prince_rounds_SR_Inv_Result_s1[61]) );
  XNOR2_X1 prince_rounds_U227 ( .A(prince_rounds_SR_Result_s1[61]), .B(
        prince_rounds_n369), .ZN(prince_rounds_round_inputXORkeyRCON_s1[61])
         );
  XNOR2_X1 prince_rounds_U226 ( .A(Key[61]), .B(
        prince_rounds_round_Constant[61]), .ZN(prince_rounds_n369) );
  XNOR2_X1 prince_rounds_U225 ( .A(prince_rounds_sub_Inv_Result_s1[58]), .B(
        prince_rounds_n368), .ZN(prince_rounds_SR_Inv_Result_s1[42]) );
  XNOR2_X1 prince_rounds_U224 ( .A(prince_rounds_SR_Result_s1[58]), .B(
        prince_rounds_n368), .ZN(prince_rounds_round_inputXORkeyRCON_s1[58])
         );
  XNOR2_X1 prince_rounds_U223 ( .A(Key[58]), .B(
        prince_rounds_round_Constant[58]), .ZN(prince_rounds_n368) );
  XNOR2_X1 prince_rounds_U222 ( .A(prince_rounds_sub_Inv_Result_s1[52]), .B(
        prince_rounds_n367), .ZN(prince_rounds_SR_Inv_Result_s1[20]) );
  XNOR2_X1 prince_rounds_U221 ( .A(prince_rounds_SR_Result_s1[52]), .B(
        prince_rounds_n367), .ZN(prince_rounds_round_inputXORkeyRCON_s1[52])
         );
  XNOR2_X1 prince_rounds_U220 ( .A(Key[52]), .B(
        prince_rounds_round_Constant[60]), .ZN(prince_rounds_n367) );
  XNOR2_X1 prince_rounds_U219 ( .A(prince_rounds_sub_Inv_Result_s1[40]), .B(
        prince_rounds_n366), .ZN(prince_rounds_SR_Inv_Result_s1[24]) );
  XNOR2_X1 prince_rounds_U218 ( .A(prince_rounds_SR_Result_s1[40]), .B(
        prince_rounds_n366), .ZN(prince_rounds_round_inputXORkeyRCON_s1[40])
         );
  XNOR2_X1 prince_rounds_U217 ( .A(Key[40]), .B(
        prince_rounds_round_Constant[62]), .ZN(prince_rounds_n366) );
  XNOR2_X1 prince_rounds_U216 ( .A(prince_rounds_sub_Inv_Result_s1[16]), .B(
        prince_rounds_n365), .ZN(prince_rounds_SR_Inv_Result_s1[32]) );
  XNOR2_X1 prince_rounds_U215 ( .A(prince_rounds_SR_Result_s1[16]), .B(
        prince_rounds_n365), .ZN(prince_rounds_round_inputXORkeyRCON_s1[16])
         );
  XNOR2_X1 prince_rounds_U214 ( .A(Key[16]), .B(
        prince_rounds_round_Constant[61]), .ZN(prince_rounds_n365) );
  XNOR2_X1 prince_rounds_U213 ( .A(prince_rounds_sub_Inv_Result_s1[0]), .B(
        prince_rounds_n364), .ZN(prince_rounds_SR_Inv_Result_s1[16]) );
  XNOR2_X1 prince_rounds_U212 ( .A(prince_rounds_SR_Result_s1[0]), .B(
        prince_rounds_n364), .ZN(prince_rounds_round_inputXORkeyRCON_s1[0]) );
  XNOR2_X1 prince_rounds_U211 ( .A(Key[0]), .B(
        prince_rounds_round_Constant[53]), .ZN(prince_rounds_n364) );
  XNOR2_X1 prince_rounds_U210 ( .A(prince_rounds_sub_Inv_Result_s1[39]), .B(
        prince_rounds_n363), .ZN(prince_rounds_SR_Inv_Result_s1[7]) );
  XNOR2_X1 prince_rounds_U209 ( .A(prince_rounds_SR_Result_s1[39]), .B(
        prince_rounds_n363), .ZN(prince_rounds_round_inputXORkeyRCON_s1[39])
         );
  XNOR2_X1 prince_rounds_U208 ( .A(Key[39]), .B(
        prince_rounds_round_Constant[39]), .ZN(prince_rounds_n363) );
  XNOR2_X1 prince_rounds_U207 ( .A(prince_rounds_sub_Inv_Result_s1[14]), .B(
        prince_rounds_n362), .ZN(prince_rounds_SR_Inv_Result_s1[14]) );
  XNOR2_X1 prince_rounds_U206 ( .A(prince_rounds_SR_Result_s1[14]), .B(
        prince_rounds_n362), .ZN(prince_rounds_round_inputXORkeyRCON_s1[14])
         );
  XNOR2_X1 prince_rounds_U205 ( .A(Key[14]), .B(
        prince_rounds_round_Constant[14]), .ZN(prince_rounds_n362) );
  XNOR2_X1 prince_rounds_U204 ( .A(prince_rounds_sub_Inv_Result_s1[13]), .B(
        prince_rounds_n361), .ZN(prince_rounds_SR_Inv_Result_s1[13]) );
  XNOR2_X1 prince_rounds_U203 ( .A(prince_rounds_SR_Result_s1[13]), .B(
        prince_rounds_n361), .ZN(prince_rounds_round_inputXORkeyRCON_s1[13])
         );
  XNOR2_X1 prince_rounds_U202 ( .A(Key[13]), .B(
        prince_rounds_round_Constant[13]), .ZN(prince_rounds_n361) );
  XNOR2_X1 prince_rounds_U201 ( .A(prince_rounds_sub_Inv_Result_s1[51]), .B(
        prince_rounds_n360), .ZN(prince_rounds_SR_Inv_Result_s1[3]) );
  XNOR2_X1 prince_rounds_U200 ( .A(prince_rounds_SR_Result_s1[51]), .B(
        prince_rounds_n360), .ZN(prince_rounds_round_inputXORkeyRCON_s1[51])
         );
  XNOR2_X1 prince_rounds_U199 ( .A(Key[51]), .B(
        prince_rounds_round_Constant[51]), .ZN(prince_rounds_n360) );
  XNOR2_X1 prince_rounds_U198 ( .A(prince_rounds_sub_Inv_Result_s1[38]), .B(
        prince_rounds_n359), .ZN(prince_rounds_SR_Inv_Result_s1[6]) );
  XNOR2_X1 prince_rounds_U197 ( .A(prince_rounds_SR_Result_s1[38]), .B(
        prince_rounds_n359), .ZN(prince_rounds_round_inputXORkeyRCON_s1[38])
         );
  XNOR2_X1 prince_rounds_U196 ( .A(Key[38]), .B(
        prince_rounds_round_Constant[38]), .ZN(prince_rounds_n359) );
  XNOR2_X1 prince_rounds_U195 ( .A(prince_rounds_sub_Inv_Result_s1[12]), .B(
        prince_rounds_n358), .ZN(prince_rounds_SR_Inv_Result_s1[12]) );
  XNOR2_X1 prince_rounds_U194 ( .A(prince_rounds_SR_Result_s1[12]), .B(
        prince_rounds_n358), .ZN(prince_rounds_round_inputXORkeyRCON_s1[12])
         );
  XNOR2_X1 prince_rounds_U193 ( .A(Key[12]), .B(
        prince_rounds_round_Constant[37]), .ZN(prince_rounds_n358) );
  XNOR2_X1 prince_rounds_U192 ( .A(prince_rounds_sub_Inv_Result_s1[11]), .B(
        prince_rounds_n357), .ZN(prince_rounds_SR_Inv_Result_s1[59]) );
  XNOR2_X1 prince_rounds_U191 ( .A(prince_rounds_SR_Result_s1[11]), .B(
        prince_rounds_n357), .ZN(prince_rounds_round_inputXORkeyRCON_s1[11])
         );
  XNOR2_X1 prince_rounds_U190 ( .A(Key[11]), .B(
        prince_rounds_round_Constant[59]), .ZN(prince_rounds_n357) );
  XNOR2_X1 prince_rounds_U189 ( .A(prince_rounds_sub_Inv_Result_s1[37]), .B(
        prince_rounds_n356), .ZN(prince_rounds_SR_Inv_Result_s1[5]) );
  XNOR2_X1 prince_rounds_U188 ( .A(prince_rounds_SR_Result_s1[37]), .B(
        prince_rounds_n356), .ZN(prince_rounds_round_inputXORkeyRCON_s1[37])
         );
  XNOR2_X1 prince_rounds_U187 ( .A(Key[37]), .B(
        prince_rounds_round_Constant[37]), .ZN(prince_rounds_n356) );
  XNOR2_X1 prince_rounds_U186 ( .A(prince_rounds_sub_Inv_Result_s1[10]), .B(
        prince_rounds_n355), .ZN(prince_rounds_SR_Inv_Result_s1[58]) );
  XNOR2_X1 prince_rounds_U185 ( .A(prince_rounds_SR_Result_s1[10]), .B(
        prince_rounds_n355), .ZN(prince_rounds_round_inputXORkeyRCON_s1[10])
         );
  XNOR2_X1 prince_rounds_U184 ( .A(Key[10]), .B(
        prince_rounds_round_Constant[59]), .ZN(prince_rounds_n355) );
  XNOR2_X1 prince_rounds_U183 ( .A(prince_rounds_sub_Inv_Result_s1[9]), .B(
        prince_rounds_n354), .ZN(prince_rounds_SR_Inv_Result_s1[57]) );
  XNOR2_X1 prince_rounds_U182 ( .A(prince_rounds_SR_Result_s1[9]), .B(
        prince_rounds_n354), .ZN(prince_rounds_round_inputXORkeyRCON_s1[9]) );
  XNOR2_X1 prince_rounds_U181 ( .A(Key[9]), .B(
        prince_rounds_round_Constant[56]), .ZN(prince_rounds_n354) );
  XNOR2_X1 prince_rounds_U180 ( .A(prince_rounds_sub_Inv_Result_s1[57]), .B(
        prince_rounds_n353), .ZN(prince_rounds_SR_Inv_Result_s1[41]) );
  XNOR2_X1 prince_rounds_U179 ( .A(prince_rounds_SR_Result_s1[57]), .B(
        prince_rounds_n353), .ZN(prince_rounds_round_inputXORkeyRCON_s1[57])
         );
  XNOR2_X1 prince_rounds_U178 ( .A(Key[57]), .B(
        prince_rounds_round_Constant[60]), .ZN(prince_rounds_n353) );
  XNOR2_X1 prince_rounds_U177 ( .A(prince_rounds_sub_Inv_Result_s1[50]), .B(
        prince_rounds_n352), .ZN(prince_rounds_SR_Inv_Result_s1[2]) );
  XNOR2_X1 prince_rounds_U176 ( .A(prince_rounds_SR_Result_s1[50]), .B(
        prince_rounds_n352), .ZN(prince_rounds_round_inputXORkeyRCON_s1[50])
         );
  XNOR2_X1 prince_rounds_U175 ( .A(Key[50]), .B(
        prince_rounds_round_Constant[50]), .ZN(prince_rounds_n352) );
  XNOR2_X1 prince_rounds_U174 ( .A(prince_rounds_sub_Inv_Result_s1[36]), .B(
        prince_rounds_n351), .ZN(prince_rounds_SR_Inv_Result_s1[4]) );
  XNOR2_X1 prince_rounds_U173 ( .A(prince_rounds_SR_Result_s1[36]), .B(
        prince_rounds_n351), .ZN(prince_rounds_round_inputXORkeyRCON_s1[36])
         );
  XNOR2_X1 prince_rounds_U172 ( .A(Key[36]), .B(
        prince_rounds_round_Constant[36]), .ZN(prince_rounds_n351) );
  XNOR2_X1 prince_rounds_U171 ( .A(prince_rounds_sub_Inv_Result_s1[8]), .B(
        prince_rounds_n350), .ZN(prince_rounds_SR_Inv_Result_s1[56]) );
  XNOR2_X1 prince_rounds_U170 ( .A(prince_rounds_SR_Result_s1[8]), .B(
        prince_rounds_n350), .ZN(prince_rounds_round_inputXORkeyRCON_s1[8]) );
  XNOR2_X1 prince_rounds_U169 ( .A(Key[8]), .B(prince_rounds_round_Constant[8]), .ZN(prince_rounds_n350) );
  XNOR2_X1 prince_rounds_U168 ( .A(prince_rounds_sub_Inv_Result_s1[7]), .B(
        prince_rounds_n349), .ZN(prince_rounds_SR_Inv_Result_s1[39]) );
  XNOR2_X1 prince_rounds_U167 ( .A(prince_rounds_SR_Result_s1[7]), .B(
        prince_rounds_n349), .ZN(prince_rounds_round_inputXORkeyRCON_s1[7]) );
  XNOR2_X1 prince_rounds_U166 ( .A(Key[7]), .B(
        prince_rounds_round_Constant[18]), .ZN(prince_rounds_n349) );
  XNOR2_X1 prince_rounds_U165 ( .A(prince_rounds_sub_Inv_Result_s1[35]), .B(
        prince_rounds_n348), .ZN(prince_rounds_SR_Inv_Result_s1[51]) );
  XNOR2_X1 prince_rounds_U164 ( .A(prince_rounds_SR_Result_s1[35]), .B(
        prince_rounds_n348), .ZN(prince_rounds_round_inputXORkeyRCON_s1[35])
         );
  XNOR2_X1 prince_rounds_U163 ( .A(Key[35]), .B(
        prince_rounds_round_Constant[41]), .ZN(prince_rounds_n348) );
  XNOR2_X1 prince_rounds_U162 ( .A(prince_rounds_sub_Inv_Result_s1[6]), .B(
        prince_rounds_n347), .ZN(prince_rounds_SR_Inv_Result_s1[38]) );
  XNOR2_X1 prince_rounds_U161 ( .A(prince_rounds_SR_Result_s1[6]), .B(
        prince_rounds_n347), .ZN(prince_rounds_round_inputXORkeyRCON_s1[6]) );
  XNOR2_X1 prince_rounds_U160 ( .A(Key[6]), .B(
        prince_rounds_round_Constant[33]), .ZN(prince_rounds_n347) );
  XNOR2_X1 prince_rounds_U159 ( .A(prince_rounds_sub_Inv_Result_s1[5]), .B(
        prince_rounds_n346), .ZN(prince_rounds_SR_Inv_Result_s1[37]) );
  XNOR2_X1 prince_rounds_U158 ( .A(prince_rounds_SR_Result_s1[5]), .B(
        prince_rounds_n346), .ZN(prince_rounds_round_inputXORkeyRCON_s1[5]) );
  XNOR2_X1 prince_rounds_U157 ( .A(Key[5]), .B(
        prince_rounds_round_Constant[38]), .ZN(prince_rounds_n346) );
  XNOR2_X1 prince_rounds_U156 ( .A(prince_rounds_sub_Inv_Result_s1[49]), .B(
        prince_rounds_n345), .ZN(prince_rounds_SR_Inv_Result_s1[1]) );
  XNOR2_X1 prince_rounds_U155 ( .A(prince_rounds_SR_Result_s1[49]), .B(
        prince_rounds_n345), .ZN(prince_rounds_round_inputXORkeyRCON_s1[49])
         );
  XNOR2_X1 prince_rounds_U154 ( .A(Key[49]), .B(
        prince_rounds_round_Constant[49]), .ZN(prince_rounds_n345) );
  XNOR2_X1 prince_rounds_U153 ( .A(prince_rounds_sub_Inv_Result_s1[34]), .B(
        prince_rounds_n344), .ZN(prince_rounds_SR_Inv_Result_s1[50]) );
  XNOR2_X1 prince_rounds_U152 ( .A(prince_rounds_SR_Result_s1[34]), .B(
        prince_rounds_n344), .ZN(prince_rounds_round_inputXORkeyRCON_s1[34])
         );
  XNOR2_X1 prince_rounds_U151 ( .A(Key[34]), .B(
        prince_rounds_round_Constant[34]), .ZN(prince_rounds_n344) );
  XNOR2_X1 prince_rounds_U150 ( .A(prince_rounds_sub_Inv_Result_s1[4]), .B(
        prince_rounds_n343), .ZN(prince_rounds_SR_Inv_Result_s1[36]) );
  XNOR2_X1 prince_rounds_U149 ( .A(prince_rounds_SR_Result_s1[4]), .B(
        prince_rounds_n343), .ZN(prince_rounds_round_inputXORkeyRCON_s1[4]) );
  XNOR2_X1 prince_rounds_U148 ( .A(Key[4]), .B(prince_rounds_round_Constant[4]), .ZN(prince_rounds_n343) );
  XNOR2_X1 prince_rounds_U147 ( .A(prince_rounds_sub_Inv_Result_s1[3]), .B(
        prince_rounds_n342), .ZN(prince_rounds_SR_Inv_Result_s1[19]) );
  XNOR2_X1 prince_rounds_U146 ( .A(prince_rounds_SR_Result_s1[3]), .B(
        prince_rounds_n342), .ZN(prince_rounds_round_inputXORkeyRCON_s1[3]) );
  XNOR2_X1 prince_rounds_U145 ( .A(Key[3]), .B(
        prince_rounds_round_Constant[50]), .ZN(prince_rounds_n342) );
  XNOR2_X1 prince_rounds_U144 ( .A(prince_rounds_sub_Inv_Result_s1[33]), .B(
        prince_rounds_n341), .ZN(prince_rounds_SR_Inv_Result_s1[49]) );
  XNOR2_X1 prince_rounds_U143 ( .A(prince_rounds_SR_Result_s1[33]), .B(
        prince_rounds_n341), .ZN(prince_rounds_round_inputXORkeyRCON_s1[33])
         );
  XNOR2_X1 prince_rounds_U142 ( .A(Key[33]), .B(
        prince_rounds_round_Constant[33]), .ZN(prince_rounds_n341) );
  XNOR2_X1 prince_rounds_U141 ( .A(prince_rounds_sub_Inv_Result_s1[2]), .B(
        prince_rounds_n340), .ZN(prince_rounds_SR_Inv_Result_s1[18]) );
  XNOR2_X1 prince_rounds_U140 ( .A(prince_rounds_SR_Result_s1[2]), .B(
        prince_rounds_n340), .ZN(prince_rounds_round_inputXORkeyRCON_s1[2]) );
  XNOR2_X1 prince_rounds_U139 ( .A(Key[2]), .B(
        prince_rounds_round_Constant[34]), .ZN(prince_rounds_n340) );
  XOR2_X1 prince_rounds_U138 ( .A(Key[15]), .B(prince_rounds_SR_Result_s1[15]), 
        .Z(prince_rounds_round_inputXORkeyRCON_s1[15]) );
  MUX2_X1 prince_rounds_U137 ( .A(prince_rounds_sub_Inv_Result_s1[15]), .B(
        prince_rounds_SR_Inv_Result_s1[15]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[15]) );
  MUX2_X1 prince_rounds_U136 ( .A(output_s2[55]), .B(output_s2[23]), .S(
        prince_rounds_n339), .Z(prince_rounds_mul_input_s2[55]) );
  MUX2_X1 prince_rounds_U135 ( .A(output_s2[50]), .B(output_s2[34]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[50]) );
  MUX2_X1 prince_rounds_U134 ( .A(output_s2[57]), .B(output_s2[9]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[57]) );
  MUX2_X1 prince_rounds_U133 ( .A(output_s2[52]), .B(output_s2[20]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[52]) );
  MUX2_X1 prince_rounds_U132 ( .A(output_s2[54]), .B(output_s2[22]), .S(
        prince_rounds_n336), .Z(prince_rounds_mul_input_s2[54]) );
  MUX2_X1 prince_rounds_U131 ( .A(output_s2[49]), .B(output_s2[33]), .S(
        prince_rounds_n335), .Z(prince_rounds_mul_input_s2[49]) );
  MUX2_X1 prince_rounds_U130 ( .A(output_s2[48]), .B(output_s2[32]), .S(
        prince_rounds_n334), .Z(prince_rounds_mul_input_s2[48]) );
  MUX2_X1 prince_rounds_U129 ( .A(output_s2[51]), .B(output_s2[35]), .S(
        roundEnd_Select_Signal), .Z(prince_rounds_mul_input_s2[51]) );
  MUX2_X1 prince_rounds_U128 ( .A(output_s2[39]), .B(output_s2[7]), .S(
        prince_rounds_n336), .Z(prince_rounds_mul_input_s2[39]) );
  MUX2_X1 prince_rounds_U127 ( .A(output_s2[34]), .B(output_s2[18]), .S(
        roundEnd_Select_Signal), .Z(prince_rounds_mul_input_s2[34]) );
  MUX2_X1 prince_rounds_U126 ( .A(output_s2[37]), .B(output_s2[5]), .S(
        prince_rounds_n339), .Z(prince_rounds_mul_input_s2[37]) );
  MUX2_X1 prince_rounds_U125 ( .A(output_s2[40]), .B(output_s2[56]), .S(
        roundEnd_Select_Signal), .Z(prince_rounds_mul_input_s2[40]) );
  MUX2_X1 prince_rounds_U124 ( .A(output_s2[35]), .B(output_s2[19]), .S(
        prince_rounds_n334), .Z(prince_rounds_mul_input_s2[35]) );
  MUX2_X1 prince_rounds_U123 ( .A(output_s2[38]), .B(output_s2[6]), .S(
        prince_rounds_n336), .Z(prince_rounds_mul_input_s2[38]) );
  MUX2_X1 prince_rounds_U122 ( .A(output_s2[33]), .B(output_s2[17]), .S(
        prince_rounds_n339), .Z(prince_rounds_mul_input_s2[33]) );
  MUX2_X1 prince_rounds_U121 ( .A(output_s2[32]), .B(output_s2[16]), .S(
        prince_rounds_n335), .Z(prince_rounds_mul_input_s2[32]) );
  MUX2_X1 prince_rounds_U120 ( .A(output_s2[23]), .B(output_s2[55]), .S(
        prince_rounds_n334), .Z(prince_rounds_mul_input_s2[23]) );
  MUX2_X1 prince_rounds_U119 ( .A(output_s2[18]), .B(output_s2[2]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[18]) );
  MUX2_X1 prince_rounds_U118 ( .A(output_s2[17]), .B(output_s2[1]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[17]) );
  MUX2_X1 prince_rounds_U117 ( .A(output_s2[16]), .B(output_s2[0]), .S(
        prince_rounds_n335), .Z(prince_rounds_mul_input_s2[16]) );
  MUX2_X1 prince_rounds_U116 ( .A(output_s2[19]), .B(output_s2[3]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[19]) );
  MUX2_X1 prince_rounds_U115 ( .A(output_s2[26]), .B(output_s2[42]), .S(
        prince_rounds_n334), .Z(prince_rounds_mul_input_s2[26]) );
  MUX2_X1 prince_rounds_U114 ( .A(output_s2[25]), .B(output_s2[41]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[25]) );
  MUX2_X1 prince_rounds_U113 ( .A(output_s2[20]), .B(output_s2[52]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[20]) );
  MUX2_X1 prince_rounds_U112 ( .A(output_s2[11]), .B(output_s2[27]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[11]) );
  MUX2_X1 prince_rounds_U111 ( .A(output_s2[14]), .B(output_s2[14]), .S(
        prince_rounds_n339), .Z(prince_rounds_mul_input_s2[14]) );
  MUX2_X1 prince_rounds_U110 ( .A(output_s2[13]), .B(output_s2[13]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[13]) );
  MUX2_X1 prince_rounds_U109 ( .A(output_s2[12]), .B(output_s2[12]), .S(
        prince_rounds_n339), .Z(prince_rounds_mul_input_s2[12]) );
  MUX2_X1 prince_rounds_U108 ( .A(output_s2[10]), .B(output_s2[26]), .S(
        prince_rounds_n334), .Z(prince_rounds_mul_input_s2[10]) );
  MUX2_X1 prince_rounds_U107 ( .A(output_s2[1]), .B(output_s2[49]), .S(
        prince_rounds_n336), .Z(prince_rounds_mul_input_s2[1]) );
  MUX2_X1 prince_rounds_U106 ( .A(output_s2[15]), .B(output_s2[15]), .S(
        prince_rounds_n335), .Z(prince_rounds_mul_input_s2[15]) );
  MUX2_X1 prince_rounds_U105 ( .A(output_s2[0]), .B(output_s2[48]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[0]) );
  MUX2_X1 prince_rounds_U104 ( .A(output_s2[9]), .B(output_s2[25]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[9]) );
  MUX2_X1 prince_rounds_U103 ( .A(output_s2[59]), .B(output_s2[11]), .S(
        prince_rounds_n339), .Z(prince_rounds_mul_input_s2[59]) );
  MUX2_X1 prince_rounds_U102 ( .A(output_s2[62]), .B(output_s2[62]), .S(
        prince_rounds_n336), .Z(prince_rounds_mul_input_s2[62]) );
  MUX2_X1 prince_rounds_U101 ( .A(output_s2[61]), .B(output_s2[61]), .S(
        prince_rounds_n335), .Z(prince_rounds_mul_input_s2[61]) );
  MUX2_X1 prince_rounds_U100 ( .A(output_s2[60]), .B(output_s2[60]), .S(
        prince_rounds_n334), .Z(prince_rounds_mul_input_s2[60]) );
  MUX2_X1 prince_rounds_U99 ( .A(output_s2[58]), .B(output_s2[10]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[58]) );
  MUX2_X1 prince_rounds_U98 ( .A(output_s2[53]), .B(output_s2[21]), .S(
        prince_rounds_n339), .Z(prince_rounds_mul_input_s2[53]) );
  MUX2_X1 prince_rounds_U97 ( .A(output_s2[56]), .B(output_s2[8]), .S(
        prince_rounds_n336), .Z(prince_rounds_mul_input_s2[56]) );
  MUX2_X1 prince_rounds_U96 ( .A(output_s2[63]), .B(output_s2[63]), .S(
        prince_rounds_n335), .Z(prince_rounds_mul_input_s2[63]) );
  MUX2_X1 prince_rounds_U95 ( .A(output_s2[43]), .B(output_s2[59]), .S(
        prince_rounds_n334), .Z(prince_rounds_mul_input_s2[43]) );
  MUX2_X1 prince_rounds_U94 ( .A(output_s2[42]), .B(output_s2[58]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[42]) );
  MUX2_X1 prince_rounds_U93 ( .A(output_s2[45]), .B(output_s2[45]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[45]) );
  MUX2_X1 prince_rounds_U92 ( .A(output_s2[44]), .B(output_s2[44]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[44]) );
  MUX2_X1 prince_rounds_U91 ( .A(output_s2[47]), .B(output_s2[47]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[47]) );
  MUX2_X1 prince_rounds_U90 ( .A(output_s2[46]), .B(output_s2[46]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[46]) );
  MUX2_X1 prince_rounds_U89 ( .A(output_s2[41]), .B(output_s2[57]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[41]) );
  MUX2_X1 prince_rounds_U88 ( .A(output_s2[36]), .B(output_s2[4]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[36]) );
  MUX2_X1 prince_rounds_U87 ( .A(output_s2[27]), .B(output_s2[43]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[27]) );
  MUX2_X1 prince_rounds_U86 ( .A(output_s2[22]), .B(output_s2[54]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[22]) );
  MUX2_X1 prince_rounds_U85 ( .A(output_s2[21]), .B(output_s2[53]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[21]) );
  MUX2_X1 prince_rounds_U84 ( .A(output_s2[28]), .B(output_s2[28]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[28]) );
  MUX2_X1 prince_rounds_U83 ( .A(output_s2[31]), .B(output_s2[31]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[31]) );
  MUX2_X1 prince_rounds_U82 ( .A(output_s2[30]), .B(output_s2[30]), .S(
        prince_rounds_n337), .Z(prince_rounds_mul_input_s2[30]) );
  INV_X1 prince_rounds_U81 ( .A(prince_rounds_n333), .ZN(prince_rounds_n337)
         );
  MUX2_X1 prince_rounds_U80 ( .A(output_s2[29]), .B(output_s2[29]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[29]) );
  MUX2_X1 prince_rounds_U79 ( .A(output_s2[24]), .B(output_s2[40]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[24]) );
  MUX2_X1 prince_rounds_U78 ( .A(output_s2[7]), .B(output_s2[39]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[7]) );
  MUX2_X1 prince_rounds_U77 ( .A(output_s2[6]), .B(output_s2[38]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[6]) );
  MUX2_X1 prince_rounds_U76 ( .A(output_s2[8]), .B(output_s2[24]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[8]) );
  MUX2_X1 prince_rounds_U75 ( .A(output_s2[2]), .B(output_s2[50]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[2]) );
  MUX2_X1 prince_rounds_U74 ( .A(output_s2[5]), .B(output_s2[37]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[5]) );
  MUX2_X1 prince_rounds_U73 ( .A(output_s2[3]), .B(output_s2[51]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[3]) );
  MUX2_X1 prince_rounds_U72 ( .A(output_s2[4]), .B(output_s2[36]), .S(
        prince_rounds_n338), .Z(prince_rounds_mul_input_s2[4]) );
  XOR2_X1 prince_rounds_U71 ( .A(prince_rounds_sub_Inv_Result_s1[15]), .B(
        Key[15]), .Z(prince_rounds_SR_Inv_Result_s1[15]) );
  MUX2_X1 prince_rounds_U70 ( .A(prince_rounds_sub_Inv_Result_s1[0]), .B(
        prince_rounds_SR_Inv_Result_s1[0]), .S(prince_rounds_n338), .Z(
        prince_rounds_mul_input_s1[0]) );
  MUX2_X1 prince_rounds_U69 ( .A(prince_rounds_sub_Inv_Result_s1[55]), .B(
        prince_rounds_SR_Inv_Result_s1[55]), .S(prince_rounds_n338), .Z(
        prince_rounds_mul_input_s1[55]) );
  MUX2_X1 prince_rounds_U68 ( .A(prince_rounds_sub_Inv_Result_s1[50]), .B(
        prince_rounds_SR_Inv_Result_s1[50]), .S(prince_rounds_n338), .Z(
        prince_rounds_mul_input_s1[50]) );
  INV_X1 prince_rounds_U67 ( .A(prince_rounds_n333), .ZN(prince_rounds_n338)
         );
  MUX2_X1 prince_rounds_U66 ( .A(prince_rounds_sub_Inv_Result_s1[57]), .B(
        prince_rounds_SR_Inv_Result_s1[57]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[57]) );
  MUX2_X1 prince_rounds_U65 ( .A(prince_rounds_sub_Inv_Result_s1[52]), .B(
        prince_rounds_SR_Inv_Result_s1[52]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[52]) );
  MUX2_X1 prince_rounds_U64 ( .A(prince_rounds_sub_Inv_Result_s1[54]), .B(
        prince_rounds_SR_Inv_Result_s1[54]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[54]) );
  MUX2_X1 prince_rounds_U63 ( .A(prince_rounds_sub_Inv_Result_s1[49]), .B(
        prince_rounds_SR_Inv_Result_s1[49]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[49]) );
  MUX2_X1 prince_rounds_U62 ( .A(prince_rounds_sub_Inv_Result_s1[48]), .B(
        prince_rounds_SR_Inv_Result_s1[48]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[48]) );
  MUX2_X1 prince_rounds_U61 ( .A(prince_rounds_sub_Inv_Result_s1[51]), .B(
        prince_rounds_SR_Inv_Result_s1[51]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[51]) );
  MUX2_X1 prince_rounds_U60 ( .A(prince_rounds_sub_Inv_Result_s1[39]), .B(
        prince_rounds_SR_Inv_Result_s1[39]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[39]) );
  MUX2_X1 prince_rounds_U59 ( .A(prince_rounds_sub_Inv_Result_s1[34]), .B(
        prince_rounds_SR_Inv_Result_s1[34]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[34]) );
  MUX2_X1 prince_rounds_U58 ( .A(prince_rounds_sub_Inv_Result_s1[37]), .B(
        prince_rounds_SR_Inv_Result_s1[37]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[37]) );
  MUX2_X1 prince_rounds_U57 ( .A(prince_rounds_sub_Inv_Result_s1[40]), .B(
        prince_rounds_SR_Inv_Result_s1[40]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[40]) );
  MUX2_X1 prince_rounds_U56 ( .A(prince_rounds_sub_Inv_Result_s1[35]), .B(
        prince_rounds_SR_Inv_Result_s1[35]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[35]) );
  MUX2_X1 prince_rounds_U55 ( .A(prince_rounds_sub_Inv_Result_s1[38]), .B(
        prince_rounds_SR_Inv_Result_s1[38]), .S(prince_rounds_n334), .Z(
        prince_rounds_mul_input_s1[38]) );
  INV_X1 prince_rounds_U54 ( .A(prince_rounds_n333), .ZN(prince_rounds_n334)
         );
  MUX2_X1 prince_rounds_U53 ( .A(prince_rounds_sub_Inv_Result_s1[33]), .B(
        prince_rounds_SR_Inv_Result_s1[33]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[33]) );
  MUX2_X1 prince_rounds_U52 ( .A(prince_rounds_sub_Inv_Result_s1[32]), .B(
        prince_rounds_SR_Inv_Result_s1[32]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[32]) );
  MUX2_X1 prince_rounds_U51 ( .A(prince_rounds_sub_Inv_Result_s1[23]), .B(
        prince_rounds_SR_Inv_Result_s1[23]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[23]) );
  MUX2_X1 prince_rounds_U50 ( .A(prince_rounds_sub_Inv_Result_s1[18]), .B(
        prince_rounds_SR_Inv_Result_s1[18]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[18]) );
  MUX2_X1 prince_rounds_U49 ( .A(prince_rounds_sub_Inv_Result_s1[17]), .B(
        prince_rounds_SR_Inv_Result_s1[17]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[17]) );
  MUX2_X1 prince_rounds_U48 ( .A(prince_rounds_sub_Inv_Result_s1[16]), .B(
        prince_rounds_SR_Inv_Result_s1[16]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[16]) );
  MUX2_X1 prince_rounds_U47 ( .A(prince_rounds_sub_Inv_Result_s1[19]), .B(
        prince_rounds_SR_Inv_Result_s1[19]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[19]) );
  MUX2_X1 prince_rounds_U46 ( .A(prince_rounds_sub_Inv_Result_s1[26]), .B(
        prince_rounds_SR_Inv_Result_s1[26]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[26]) );
  MUX2_X1 prince_rounds_U45 ( .A(prince_rounds_sub_Inv_Result_s1[25]), .B(
        prince_rounds_SR_Inv_Result_s1[25]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[25]) );
  MUX2_X1 prince_rounds_U44 ( .A(prince_rounds_sub_Inv_Result_s1[20]), .B(
        prince_rounds_SR_Inv_Result_s1[20]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[20]) );
  MUX2_X1 prince_rounds_U43 ( .A(prince_rounds_sub_Inv_Result_s1[11]), .B(
        prince_rounds_SR_Inv_Result_s1[11]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[11]) );
  MUX2_X1 prince_rounds_U42 ( .A(prince_rounds_sub_Inv_Result_s1[14]), .B(
        prince_rounds_SR_Inv_Result_s1[14]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[14]) );
  MUX2_X1 prince_rounds_U41 ( .A(prince_rounds_sub_Inv_Result_s1[13]), .B(
        prince_rounds_SR_Inv_Result_s1[13]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[13]) );
  MUX2_X1 prince_rounds_U40 ( .A(prince_rounds_sub_Inv_Result_s1[12]), .B(
        prince_rounds_SR_Inv_Result_s1[12]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[12]) );
  MUX2_X1 prince_rounds_U39 ( .A(prince_rounds_sub_Inv_Result_s1[1]), .B(
        prince_rounds_SR_Inv_Result_s1[1]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[1]) );
  MUX2_X1 prince_rounds_U38 ( .A(prince_rounds_sub_Inv_Result_s1[10]), .B(
        prince_rounds_SR_Inv_Result_s1[10]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[10]) );
  MUX2_X1 prince_rounds_U37 ( .A(prince_rounds_sub_Inv_Result_s1[4]), .B(
        prince_rounds_SR_Inv_Result_s1[4]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[4]) );
  MUX2_X1 prince_rounds_U36 ( .A(prince_rounds_sub_Inv_Result_s1[62]), .B(
        prince_rounds_SR_Inv_Result_s1[62]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[62]) );
  MUX2_X1 prince_rounds_U35 ( .A(prince_rounds_sub_Inv_Result_s1[61]), .B(
        prince_rounds_SR_Inv_Result_s1[61]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[61]) );
  MUX2_X1 prince_rounds_U34 ( .A(prince_rounds_sub_Inv_Result_s1[60]), .B(
        prince_rounds_SR_Inv_Result_s1[60]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[60]) );
  MUX2_X1 prince_rounds_U33 ( .A(prince_rounds_sub_Inv_Result_s1[53]), .B(
        prince_rounds_SR_Inv_Result_s1[53]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[53]) );
  MUX2_X1 prince_rounds_U32 ( .A(prince_rounds_sub_Inv_Result_s1[56]), .B(
        prince_rounds_SR_Inv_Result_s1[56]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[56]) );
  MUX2_X1 prince_rounds_U31 ( .A(prince_rounds_sub_Inv_Result_s1[63]), .B(
        prince_rounds_SR_Inv_Result_s1[63]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[63]) );
  MUX2_X1 prince_rounds_U30 ( .A(prince_rounds_sub_Inv_Result_s1[42]), .B(
        prince_rounds_SR_Inv_Result_s1[42]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[42]) );
  MUX2_X1 prince_rounds_U29 ( .A(prince_rounds_sub_Inv_Result_s1[45]), .B(
        prince_rounds_SR_Inv_Result_s1[45]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[45]) );
  MUX2_X1 prince_rounds_U28 ( .A(prince_rounds_sub_Inv_Result_s1[44]), .B(
        prince_rounds_SR_Inv_Result_s1[44]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[44]) );
  MUX2_X1 prince_rounds_U27 ( .A(prince_rounds_sub_Inv_Result_s1[47]), .B(
        prince_rounds_SR_Inv_Result_s1[47]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[47]) );
  MUX2_X1 prince_rounds_U26 ( .A(prince_rounds_sub_Inv_Result_s1[41]), .B(
        prince_rounds_SR_Inv_Result_s1[41]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[41]) );
  MUX2_X1 prince_rounds_U25 ( .A(prince_rounds_sub_Inv_Result_s1[36]), .B(
        prince_rounds_SR_Inv_Result_s1[36]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[36]) );
  MUX2_X1 prince_rounds_U24 ( .A(prince_rounds_sub_Inv_Result_s1[27]), .B(
        prince_rounds_SR_Inv_Result_s1[27]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[27]) );
  MUX2_X1 prince_rounds_U23 ( .A(prince_rounds_sub_Inv_Result_s1[22]), .B(
        prince_rounds_SR_Inv_Result_s1[22]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[22]) );
  MUX2_X1 prince_rounds_U22 ( .A(prince_rounds_sub_Inv_Result_s1[21]), .B(
        prince_rounds_SR_Inv_Result_s1[21]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[21]) );
  MUX2_X1 prince_rounds_U21 ( .A(prince_rounds_sub_Inv_Result_s1[28]), .B(
        prince_rounds_SR_Inv_Result_s1[28]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[28]) );
  MUX2_X1 prince_rounds_U20 ( .A(prince_rounds_sub_Inv_Result_s1[31]), .B(
        prince_rounds_SR_Inv_Result_s1[31]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[31]) );
  MUX2_X1 prince_rounds_U19 ( .A(prince_rounds_sub_Inv_Result_s1[30]), .B(
        prince_rounds_SR_Inv_Result_s1[30]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[30]) );
  MUX2_X1 prince_rounds_U18 ( .A(prince_rounds_sub_Inv_Result_s1[29]), .B(
        prince_rounds_SR_Inv_Result_s1[29]), .S(prince_rounds_n339), .Z(
        prince_rounds_mul_input_s1[29]) );
  INV_X1 prince_rounds_U17 ( .A(prince_rounds_n333), .ZN(prince_rounds_n339)
         );
  MUX2_X1 prince_rounds_U16 ( .A(prince_rounds_sub_Inv_Result_s1[24]), .B(
        prince_rounds_SR_Inv_Result_s1[24]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[24]) );
  MUX2_X1 prince_rounds_U15 ( .A(prince_rounds_sub_Inv_Result_s1[7]), .B(
        prince_rounds_SR_Inv_Result_s1[7]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[7]) );
  MUX2_X1 prince_rounds_U14 ( .A(prince_rounds_sub_Inv_Result_s1[6]), .B(
        prince_rounds_SR_Inv_Result_s1[6]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[6]) );
  MUX2_X1 prince_rounds_U13 ( .A(prince_rounds_sub_Inv_Result_s1[9]), .B(
        prince_rounds_SR_Inv_Result_s1[9]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[9]) );
  MUX2_X1 prince_rounds_U12 ( .A(prince_rounds_sub_Inv_Result_s1[8]), .B(
        prince_rounds_SR_Inv_Result_s1[8]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[8]) );
  MUX2_X1 prince_rounds_U11 ( .A(prince_rounds_sub_Inv_Result_s1[2]), .B(
        prince_rounds_SR_Inv_Result_s1[2]), .S(prince_rounds_n335), .Z(
        prince_rounds_mul_input_s1[2]) );
  INV_X1 prince_rounds_U10 ( .A(prince_rounds_n333), .ZN(prince_rounds_n335)
         );
  MUX2_X1 prince_rounds_U9 ( .A(prince_rounds_sub_Inv_Result_s1[5]), .B(
        prince_rounds_SR_Inv_Result_s1[5]), .S(prince_rounds_n336), .Z(
        prince_rounds_mul_input_s1[5]) );
  INV_X1 prince_rounds_U8 ( .A(prince_rounds_n333), .ZN(prince_rounds_n336) );
  MUX2_X1 prince_rounds_U7 ( .A(prince_rounds_sub_Inv_Result_s1[3]), .B(
        prince_rounds_SR_Inv_Result_s1[3]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[3]) );
  MUX2_X1 prince_rounds_U6 ( .A(prince_rounds_sub_Inv_Result_s1[59]), .B(
        prince_rounds_SR_Inv_Result_s1[59]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[59]) );
  MUX2_X1 prince_rounds_U5 ( .A(prince_rounds_sub_Inv_Result_s1[58]), .B(
        prince_rounds_SR_Inv_Result_s1[58]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[58]) );
  MUX2_X1 prince_rounds_U4 ( .A(prince_rounds_sub_Inv_Result_s1[43]), .B(
        prince_rounds_SR_Inv_Result_s1[43]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[43]) );
  MUX2_X1 prince_rounds_U3 ( .A(prince_rounds_sub_Inv_Result_s1[46]), .B(
        prince_rounds_SR_Inv_Result_s1[46]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s1[46]) );
  INV_X1 prince_rounds_U2 ( .A(roundEnd_Select_Signal), .ZN(prince_rounds_n333) );
  NAND2_X1 prince_rounds_constant_MUX_U90 ( .A1(prince_rounds_constant_MUX_n56), .A2(prince_rounds_constant_MUX_n55), .ZN(prince_rounds_round_Constant[63])
         );
  NAND2_X1 prince_rounds_constant_MUX_U89 ( .A1(prince_rounds_constant_MUX_n54), .A2(prince_rounds_constant_MUX_n53), .ZN(prince_rounds_round_Constant[55])
         );
  NAND2_X1 prince_rounds_constant_MUX_U88 ( .A1(prince_rounds_constant_MUX_n52), .A2(prince_rounds_constant_MUX_n51), .ZN(prince_rounds_round_Constant[51])
         );
  NAND2_X1 prince_rounds_constant_MUX_U87 ( .A1(prince_rounds_constant_MUX_n50), .A2(prince_rounds_constant_MUX_n49), .ZN(prince_rounds_round_Constant[45])
         );
  NAND2_X1 prince_rounds_constant_MUX_U86 ( .A1(prince_rounds_constant_MUX_n48), .A2(prince_rounds_constant_MUX_n51), .ZN(prince_rounds_round_Constant[43])
         );
  NAND2_X1 prince_rounds_constant_MUX_U85 ( .A1(prince_rounds_constant_MUX_n47), .A2(prince_rounds_constant_MUX_n49), .ZN(prince_rounds_round_Constant[39])
         );
  NAND2_X1 prince_rounds_constant_MUX_U84 ( .A1(prince_rounds_constant_MUX_n46), .A2(prince_rounds_constant_MUX_n45), .ZN(prince_rounds_round_Constant[58])
         );
  NAND2_X1 prince_rounds_constant_MUX_U83 ( .A1(prince_rounds_constant_MUX_n44), .A2(prince_rounds_constant_MUX_n45), .ZN(prince_rounds_round_Constant[29])
         );
  INV_X1 prince_rounds_constant_MUX_U82 ( .A(prince_rounds_round_Constant[38]), 
        .ZN(prince_rounds_constant_MUX_n45) );
  NAND2_X1 prince_rounds_constant_MUX_U81 ( .A1(prince_rounds_constant_MUX_n43), .A2(prince_rounds_constant_MUX_n50), .ZN(prince_rounds_round_Constant[27])
         );
  NAND2_X1 prince_rounds_constant_MUX_U80 ( .A1(prince_rounds_constant_MUX_n56), .A2(prince_rounds_constant_MUX_n42), .ZN(prince_rounds_round_Constant[21])
         );
  NAND2_X1 prince_rounds_constant_MUX_U79 ( .A1(prince_rounds_constant_MUX_n56), .A2(prince_rounds_constant_MUX_n50), .ZN(prince_rounds_round_Constant[19])
         );
  NAND2_X1 prince_rounds_constant_MUX_U78 ( .A1(prince_rounds_constant_MUX_n41), .A2(prince_rounds_constant_MUX_n46), .ZN(prince_rounds_round_Constant[48])
         );
  NAND2_X1 prince_rounds_constant_MUX_U77 ( .A1(prince_rounds_constant_MUX_n41), .A2(prince_rounds_constant_MUX_n44), .ZN(prince_rounds_round_Constant[13])
         );
  NAND2_X1 prince_rounds_constant_MUX_U76 ( .A1(prince_rounds_constant_MUX_n40), .A2(prince_rounds_constant_MUX_n49), .ZN(prince_rounds_round_Constant[22])
         );
  NAND2_X1 prince_rounds_constant_MUX_U75 ( .A1(prince_rounds_constant_MUX_n40), .A2(prince_rounds_constant_MUX_n53), .ZN(prince_rounds_round_Constant[14])
         );
  NOR2_X1 prince_rounds_constant_MUX_U74 ( .A1(prince_rounds_constant_MUX_n39), 
        .A2(prince_rounds_constant_MUX_n38), .ZN(
        prince_rounds_constant_MUX_n40) );
  NAND2_X1 prince_rounds_constant_MUX_U73 ( .A1(prince_rounds_constant_MUX_n56), .A2(prince_rounds_constant_MUX_n37), .ZN(prince_rounds_round_Constant[32])
         );
  NAND2_X1 prince_rounds_constant_MUX_U72 ( .A1(prince_rounds_constant_MUX_n48), .A2(prince_rounds_constant_MUX_n36), .ZN(prince_rounds_round_Constant[24])
         );
  NOR2_X1 prince_rounds_constant_MUX_U71 ( .A1(prince_rounds_constant_MUX_n35), 
        .A2(prince_rounds_constant_MUX_n34), .ZN(
        prince_rounds_constant_MUX_n48) );
  NAND2_X1 prince_rounds_constant_MUX_U70 ( .A1(prince_rounds_constant_MUX_n33), .A2(prince_rounds_constant_MUX_n46), .ZN(prince_rounds_round_Constant[8]) );
  NAND2_X1 prince_rounds_constant_MUX_U69 ( .A1(prince_rounds_constant_MUX_n43), .A2(prince_rounds_constant_MUX_n55), .ZN(prince_rounds_round_Constant[4]) );
  NOR2_X1 prince_rounds_constant_MUX_U68 ( .A1(prince_rounds_constant_MUX_n32), 
        .A2(prince_rounds_constant_MUX_n31), .ZN(
        prince_rounds_constant_MUX_n55) );
  NAND2_X1 prince_rounds_constant_MUX_U67 ( .A1(prince_rounds_constant_MUX_n36), .A2(prince_rounds_constant_MUX_n30), .ZN(prince_rounds_constant_MUX_n31) );
  NAND2_X1 prince_rounds_constant_MUX_U66 ( .A1(prince_rounds_constant_MUX_n52), .A2(prince_rounds_constant_MUX_n36), .ZN(prince_rounds_round_Constant[37])
         );
  NOR2_X1 prince_rounds_constant_MUX_U65 ( .A1(prince_rounds_constant_MUX_n34), 
        .A2(prince_rounds_constant_MUX_n29), .ZN(
        prince_rounds_constant_MUX_n52) );
  NAND2_X1 prince_rounds_constant_MUX_U64 ( .A1(prince_rounds_constant_MUX_n28), .A2(prince_rounds_constant_MUX_n41), .ZN(prince_rounds_round_Constant[60])
         );
  NAND2_X1 prince_rounds_constant_MUX_U63 ( .A1(prince_rounds_constant_MUX_n27), .A2(prince_rounds_constant_MUX_n36), .ZN(prince_rounds_round_Constant[33])
         );
  NOR2_X1 prince_rounds_constant_MUX_U62 ( .A1(prince_rounds_constant_MUX_n26), 
        .A2(prince_rounds_constant_MUX_n34), .ZN(
        prince_rounds_constant_MUX_n27) );
  NAND2_X1 prince_rounds_constant_MUX_U61 ( .A1(prince_rounds_constant_MUX_n25), .A2(prince_rounds_constant_MUX_n30), .ZN(prince_rounds_constant_MUX_n34) );
  NAND2_X1 prince_rounds_constant_MUX_U60 ( .A1(prince_rounds_constant_MUX_n42), .A2(prince_rounds_constant_MUX_n49), .ZN(prince_rounds_round_Constant[34])
         );
  NOR2_X1 prince_rounds_constant_MUX_U59 ( .A1(prince_rounds_constant_MUX_n24), 
        .A2(prince_rounds_constant_MUX_n39), .ZN(
        prince_rounds_constant_MUX_n42) );
  INV_X1 prince_rounds_constant_MUX_U58 ( .A(prince_rounds_constant_MUX_n25), 
        .ZN(prince_rounds_constant_MUX_n39) );
  NAND2_X1 prince_rounds_constant_MUX_U57 ( .A1(prince_rounds_constant_MUX_n23), .A2(prince_rounds_constant_MUX_n22), .ZN(prince_rounds_constant_MUX_n25) );
  XNOR2_X1 prince_rounds_constant_MUX_U56 ( .A(roundEnd_Select_Signal), .B(
        round_Signal[2]), .ZN(prince_rounds_constant_MUX_n23) );
  NAND2_X1 prince_rounds_constant_MUX_U55 ( .A1(prince_rounds_constant_MUX_n50), .A2(prince_rounds_constant_MUX_n53), .ZN(prince_rounds_round_Constant[18])
         );
  NOR2_X1 prince_rounds_constant_MUX_U54 ( .A1(prince_rounds_constant_MUX_n21), 
        .A2(prince_rounds_constant_MUX_n32), .ZN(
        prince_rounds_constant_MUX_n50) );
  NAND2_X1 prince_rounds_constant_MUX_U53 ( .A1(prince_rounds_constant_MUX_n43), .A2(prince_rounds_constant_MUX_n37), .ZN(prince_rounds_round_Constant[62])
         );
  NAND2_X1 prince_rounds_constant_MUX_U52 ( .A1(prince_rounds_constant_MUX_n20), .A2(prince_rounds_constant_MUX_n53), .ZN(prince_rounds_constant_MUX_n37) );
  NAND2_X1 prince_rounds_constant_MUX_U51 ( .A1(prince_rounds_constant_MUX_n43), .A2(prince_rounds_constant_MUX_n47), .ZN(prince_rounds_round_Constant[53])
         );
  INV_X1 prince_rounds_constant_MUX_U50 ( .A(prince_rounds_constant_MUX_n29), 
        .ZN(prince_rounds_constant_MUX_n43) );
  NAND2_X1 prince_rounds_constant_MUX_U49 ( .A1(prince_rounds_constant_MUX_n19), .A2(prince_rounds_constant_MUX_n18), .ZN(prince_rounds_constant_MUX_n29) );
  NAND2_X1 prince_rounds_constant_MUX_U48 ( .A1(prince_rounds_constant_MUX_n47), .A2(prince_rounds_constant_MUX_n56), .ZN(prince_rounds_round_Constant[50])
         );
  AND2_X1 prince_rounds_constant_MUX_U47 ( .A1(prince_rounds_constant_MUX_n17), 
        .A2(prince_rounds_constant_MUX_n16), .ZN(
        prince_rounds_constant_MUX_n56) );
  NAND2_X1 prince_rounds_constant_MUX_U46 ( .A1(prince_rounds_constant_MUX_n47), .A2(prince_rounds_constant_MUX_n53), .ZN(prince_rounds_round_Constant[36])
         );
  NOR2_X1 prince_rounds_constant_MUX_U45 ( .A1(prince_rounds_constant_MUX_n32), 
        .A2(prince_rounds_constant_MUX_n38), .ZN(
        prince_rounds_constant_MUX_n47) );
  NAND2_X1 prince_rounds_constant_MUX_U44 ( .A1(prince_rounds_constant_MUX_n51), .A2(prince_rounds_constant_MUX_n15), .ZN(prince_rounds_constant_MUX_n38) );
  NAND2_X1 prince_rounds_constant_MUX_U43 ( .A1(prince_rounds_constant_MUX_n28), .A2(prince_rounds_constant_MUX_n46), .ZN(prince_rounds_round_Constant[61])
         );
  AND2_X1 prince_rounds_constant_MUX_U42 ( .A1(prince_rounds_constant_MUX_n30), 
        .A2(prince_rounds_constant_MUX_n15), .ZN(
        prince_rounds_constant_MUX_n46) );
  NAND2_X1 prince_rounds_constant_MUX_U41 ( .A1(prince_rounds_constant_MUX_n22), .A2(prince_rounds_constant_MUX_n24), .ZN(prince_rounds_constant_MUX_n15) );
  NAND2_X1 prince_rounds_constant_MUX_U40 ( .A1(prince_rounds_constant_MUX_n21), .A2(prince_rounds_constant_MUX_n14), .ZN(prince_rounds_constant_MUX_n30) );
  NAND2_X1 prince_rounds_constant_MUX_U39 ( .A1(prince_rounds_constant_MUX_n28), .A2(prince_rounds_constant_MUX_n13), .ZN(prince_rounds_round_Constant[59])
         );
  INV_X1 prince_rounds_constant_MUX_U38 ( .A(prince_rounds_round_Constant[54]), 
        .ZN(prince_rounds_constant_MUX_n28) );
  OR2_X1 prince_rounds_constant_MUX_U37 ( .A1(prince_rounds_round_Constant[54]), .A2(prince_rounds_round_Constant[47]), .ZN(prince_rounds_round_Constant[41])
         );
  NAND2_X1 prince_rounds_constant_MUX_U36 ( .A1(prince_rounds_constant_MUX_n41), .A2(prince_rounds_constant_MUX_n13), .ZN(prince_rounds_round_Constant[47])
         );
  INV_X1 prince_rounds_constant_MUX_U35 ( .A(prince_rounds_round_Constant[49]), 
        .ZN(prince_rounds_constant_MUX_n13) );
  INV_X1 prince_rounds_constant_MUX_U34 ( .A(prince_rounds_round_Constant[25]), 
        .ZN(prince_rounds_constant_MUX_n41) );
  NAND2_X1 prince_rounds_constant_MUX_U33 ( .A1(prince_rounds_constant_MUX_n36), .A2(prince_rounds_constant_MUX_n51), .ZN(prince_rounds_round_Constant[49])
         );
  NAND2_X1 prince_rounds_constant_MUX_U32 ( .A1(prince_rounds_constant_MUX_n22), .A2(prince_rounds_constant_MUX_n21), .ZN(prince_rounds_constant_MUX_n51) );
  NAND2_X1 prince_rounds_constant_MUX_U31 ( .A1(prince_rounds_constant_MUX_n24), .A2(prince_rounds_constant_MUX_n14), .ZN(prince_rounds_constant_MUX_n36) );
  NAND2_X1 prince_rounds_constant_MUX_U30 ( .A1(prince_rounds_constant_MUX_n18), .A2(prince_rounds_constant_MUX_n16), .ZN(prince_rounds_round_Constant[54])
         );
  NAND2_X1 prince_rounds_constant_MUX_U29 ( .A1(prince_rounds_constant_MUX_n22), .A2(prince_rounds_constant_MUX_n26), .ZN(prince_rounds_constant_MUX_n16) );
  NAND2_X1 prince_rounds_constant_MUX_U28 ( .A1(prince_rounds_constant_MUX_n35), .A2(prince_rounds_constant_MUX_n14), .ZN(prince_rounds_constant_MUX_n18) );
  INV_X1 prince_rounds_constant_MUX_U27 ( .A(prince_rounds_constant_MUX_n33), 
        .ZN(prince_rounds_round_Constant[56]) );
  NOR2_X1 prince_rounds_constant_MUX_U26 ( .A1(
        prince_rounds_round_Constant[25]), .A2(prince_rounds_round_Constant[1]), .ZN(prince_rounds_constant_MUX_n33) );
  NAND2_X1 prince_rounds_constant_MUX_U25 ( .A1(prince_rounds_constant_MUX_n19), .A2(prince_rounds_constant_MUX_n17), .ZN(prince_rounds_round_Constant[1]) );
  NAND2_X1 prince_rounds_constant_MUX_U24 ( .A1(prince_rounds_constant_MUX_n22), .A2(prince_rounds_constant_MUX_n35), .ZN(prince_rounds_constant_MUX_n17) );
  NAND2_X1 prince_rounds_constant_MUX_U23 ( .A1(prince_rounds_constant_MUX_n26), .A2(prince_rounds_constant_MUX_n14), .ZN(prince_rounds_constant_MUX_n19) );
  MUX2_X1 prince_rounds_constant_MUX_U22 ( .A(prince_rounds_constant_MUX_n12), 
        .B(prince_rounds_constant_MUX_n32), .S(prince_rounds_constant_MUX_n14), 
        .Z(prince_rounds_round_Constant[25]) );
  INV_X1 prince_rounds_constant_MUX_U21 ( .A(prince_rounds_constant_MUX_n22), 
        .ZN(prince_rounds_constant_MUX_n14) );
  XOR2_X1 prince_rounds_constant_MUX_U20 ( .A(round_Signal[0]), .B(enc_dec), 
        .Z(prince_rounds_constant_MUX_n22) );
  NOR2_X1 prince_rounds_constant_MUX_U19 ( .A1(prince_rounds_constant_MUX_n54), 
        .A2(prince_rounds_constant_MUX_n11), .ZN(
        prince_rounds_constant_MUX_n32) );
  NOR2_X1 prince_rounds_constant_MUX_U18 ( .A1(prince_rounds_constant_MUX_n20), 
        .A2(prince_rounds_constant_MUX_n10), .ZN(
        prince_rounds_constant_MUX_n12) );
  NAND2_X1 prince_rounds_constant_MUX_U17 ( .A1(prince_rounds_constant_MUX_n49), .A2(prince_rounds_constant_MUX_n53), .ZN(prince_rounds_round_Constant[38])
         );
  INV_X1 prince_rounds_constant_MUX_U16 ( .A(prince_rounds_constant_MUX_n35), 
        .ZN(prince_rounds_constant_MUX_n53) );
  NOR2_X1 prince_rounds_constant_MUX_U15 ( .A1(prince_rounds_constant_MUX_n9), 
        .A2(prince_rounds_constant_MUX_n10), .ZN(
        prince_rounds_constant_MUX_n35) );
  INV_X1 prince_rounds_constant_MUX_U14 ( .A(prince_rounds_constant_MUX_n11), 
        .ZN(prince_rounds_constant_MUX_n10) );
  INV_X1 prince_rounds_constant_MUX_U13 ( .A(prince_rounds_constant_MUX_n26), 
        .ZN(prince_rounds_constant_MUX_n49) );
  NOR2_X1 prince_rounds_constant_MUX_U12 ( .A1(prince_rounds_constant_MUX_n8), 
        .A2(prince_rounds_constant_MUX_n11), .ZN(
        prince_rounds_constant_MUX_n26) );
  INV_X1 prince_rounds_constant_MUX_U11 ( .A(prince_rounds_constant_MUX_n44), 
        .ZN(prince_rounds_round_Constant[44]) );
  NOR2_X1 prince_rounds_constant_MUX_U10 ( .A1(prince_rounds_constant_MUX_n24), 
        .A2(prince_rounds_constant_MUX_n21), .ZN(
        prince_rounds_constant_MUX_n44) );
  NOR2_X1 prince_rounds_constant_MUX_U9 ( .A1(prince_rounds_constant_MUX_n9), 
        .A2(prince_rounds_constant_MUX_n20), .ZN(
        prince_rounds_constant_MUX_n21) );
  NOR2_X1 prince_rounds_constant_MUX_U8 ( .A1(prince_rounds_constant_MUX_n8), 
        .A2(prince_rounds_constant_MUX_n54), .ZN(
        prince_rounds_constant_MUX_n24) );
  INV_X1 prince_rounds_constant_MUX_U7 ( .A(prince_rounds_constant_MUX_n20), 
        .ZN(prince_rounds_constant_MUX_n54) );
  XOR2_X1 prince_rounds_constant_MUX_U6 ( .A(enc_dec), .B(
        roundEnd_Select_Signal), .Z(prince_rounds_constant_MUX_n20) );
  INV_X1 prince_rounds_constant_MUX_U5 ( .A(prince_rounds_constant_MUX_n9), 
        .ZN(prince_rounds_constant_MUX_n8) );
  XNOR2_X1 prince_rounds_constant_MUX_U4 ( .A(enc_dec), .B(round_Signal[2]), 
        .ZN(prince_rounds_constant_MUX_n11) );
  XOR2_X1 prince_rounds_constant_MUX_U3 ( .A(enc_dec), .B(round_Signal[1]), 
        .Z(prince_rounds_constant_MUX_n9) );
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_0_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[0]), .B(prince_SR_Inv_Result_s1[0]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_0_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_0_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_0_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[48]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_1_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[1]), .B(prince_SR_Inv_Result_s1[1]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_1_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_1_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_1_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[49]), .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_2_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[2]), .B(prince_SR_Inv_Result_s1[2]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_2_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_2_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_2_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[50]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_3_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[3]), .B(prince_SR_Inv_Result_s1[3]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_3_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_3_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_3_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[51]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_4_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[4]), .B(prince_SR_Inv_Result_s1[4]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_4_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_4_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_4_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[36]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_5_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[5]), .B(prince_SR_Inv_Result_s1[5]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_5_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_5_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_5_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[37]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_6_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[6]), .B(prince_SR_Inv_Result_s1[6]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_6_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_6_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_6_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[38]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_7_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[7]), .B(prince_SR_Inv_Result_s1[7]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_7_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_7_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_7_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[39]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_8_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[8]), .B(prince_SR_Inv_Result_s1[8]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_8_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_8_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_8_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[24]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_9_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[9]), .B(prince_SR_Inv_Result_s1[9]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_9_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_9_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_9_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[25]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_10_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[10]), .B(prince_SR_Inv_Result_s1[10]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_10_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_10_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_10_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[26]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_11_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[11]), .B(prince_SR_Inv_Result_s1[11]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_11_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_11_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_11_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[27]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_12_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[12]), .B(prince_SR_Inv_Result_s1[12]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_12_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_12_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_12_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[12]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_13_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[13]), .B(prince_SR_Inv_Result_s1[13]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_13_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_13_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_13_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[13]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_14_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[14]), .B(prince_SR_Inv_Result_s1[14]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_14_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_14_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_14_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[14]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_15_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[15]), .B(prince_SR_Inv_Result_s1[15]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_15_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_15_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_15_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[15]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_16_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[16]), .B(prince_SR_Inv_Result_s1[16]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_16_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_16_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_16_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[0]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_17_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[17]), .B(prince_SR_Inv_Result_s1[17]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_17_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_17_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_17_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[1]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_18_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[18]), .B(prince_SR_Inv_Result_s1[18]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_18_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_18_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_18_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[2]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_19_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[19]), .B(prince_SR_Inv_Result_s1[19]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_19_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_19_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_19_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[3]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_20_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[20]), .B(prince_SR_Inv_Result_s1[20]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_20_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_20_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_20_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[52]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_21_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[21]), .B(prince_SR_Inv_Result_s1[21]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_21_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_21_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_21_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[53]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_22_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[22]), .B(prince_SR_Inv_Result_s1[22]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_22_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_22_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_22_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[54]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_23_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[23]), .B(prince_SR_Inv_Result_s1[23]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_23_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_23_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_23_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[55]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_24_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[24]), .B(prince_SR_Inv_Result_s1[24]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_24_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_24_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_24_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[40]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_25_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[25]), .B(prince_SR_Inv_Result_s1[25]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_25_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_25_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_25_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[41]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_26_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[26]), .B(prince_SR_Inv_Result_s1[26]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_26_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_26_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_26_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[42]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_27_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[27]), .B(prince_SR_Inv_Result_s1[27]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_27_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_27_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_27_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[43]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_28_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[28]), .B(prince_SR_Inv_Result_s1[28]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_28_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_28_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_28_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[28]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_29_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[29]), .B(prince_SR_Inv_Result_s1[29]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_29_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_29_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_29_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[29]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_30_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[30]), .B(prince_SR_Inv_Result_s1[30]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_30_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_30_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_30_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[30]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_31_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[31]), .B(prince_SR_Inv_Result_s1[31]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_31_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_31_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_31_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[31]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_32_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[32]), .B(prince_SR_Inv_Result_s1[32]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_32_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_32_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_32_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[16]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_33_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[33]), .B(prince_SR_Inv_Result_s1[33]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_33_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_33_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_33_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[17]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_34_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[34]), .B(prince_SR_Inv_Result_s1[34]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_34_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_34_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_34_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[18]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_35_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[35]), .B(prince_SR_Inv_Result_s1[35]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_35_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_35_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_35_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[19]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_36_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[36]), .B(prince_SR_Inv_Result_s1[36]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_36_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_36_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_36_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[4]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_37_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[37]), .B(prince_SR_Inv_Result_s1[37]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_37_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_37_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_37_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[5]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_38_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[38]), .B(prince_SR_Inv_Result_s1[38]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_38_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_38_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_38_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[6]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_39_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[39]), .B(prince_SR_Inv_Result_s1[39]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_39_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_39_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_39_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[7]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_40_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[40]), .B(prince_SR_Inv_Result_s1[40]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_40_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_40_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_40_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[56]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_41_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[41]), .B(prince_SR_Inv_Result_s1[41]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_41_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_41_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_41_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[57]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_42_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[42]), .B(prince_SR_Inv_Result_s1[42]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_42_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_42_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_42_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[58]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_43_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[43]), .B(prince_SR_Inv_Result_s1[43]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_43_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_43_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_43_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[59]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_44_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[44]), .B(prince_SR_Inv_Result_s1[44]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_44_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_44_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_44_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[44]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_45_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[45]), .B(prince_SR_Inv_Result_s1[45]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_45_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_45_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_45_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[45]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_46_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[46]), .B(prince_SR_Inv_Result_s1[46]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_46_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_46_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_46_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[46]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_47_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[47]), .B(prince_SR_Inv_Result_s1[47]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_47_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_47_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_47_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[47]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_48_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[48]), .B(prince_SR_Inv_Result_s1[48]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_48_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_48_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_48_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[32]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_49_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[49]), .B(prince_SR_Inv_Result_s1[49]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_49_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_49_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_49_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[33]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_50_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[50]), .B(prince_SR_Inv_Result_s1[50]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_50_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_50_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_50_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[34]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_51_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[51]), .B(prince_SR_Inv_Result_s1[51]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_51_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_51_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_51_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[35]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_52_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[52]), .B(prince_SR_Inv_Result_s1[52]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_52_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_52_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_52_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[20]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_53_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[53]), .B(prince_SR_Inv_Result_s1[53]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_53_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_53_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_53_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[21]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_54_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[54]), .B(prince_SR_Inv_Result_s1[54]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_54_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_54_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_54_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[22]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_55_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[55]), .B(prince_SR_Inv_Result_s1[55]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_55_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_55_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_55_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[23]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_56_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[56]), .B(prince_SR_Inv_Result_s1[56]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_56_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_56_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_56_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[8]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_57_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[57]), .B(prince_SR_Inv_Result_s1[57]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_57_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_57_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_57_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[9]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_58_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[58]), .B(prince_SR_Inv_Result_s1[58]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_58_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_58_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_58_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[10]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_59_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[59]), .B(prince_SR_Inv_Result_s1[59]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_59_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_59_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_59_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[11]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_60_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[60]), .B(prince_SR_Inv_Result_s1[60]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_60_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_60_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_60_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[60]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_61_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[61]), .B(prince_SR_Inv_Result_s1[61]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_61_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_61_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_61_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[61]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_62_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[62]), .B(prince_SR_Inv_Result_s1[62]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_62_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_62_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_62_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[62]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s1_SFF_63_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s1[63]), .B(prince_SR_Inv_Result_s1[63]), .S(
        rst), .Z(prince_rounds_roundResult_Reg_s1_SFF_63_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s1_SFF_63_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s1_SFF_63_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s1[63]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_0_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[0]), .B(input_s2[48]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_0_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_0_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_0_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[48]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_1_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[1]), .B(input_s2[49]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_1_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_1_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_1_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[49]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_2_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[2]), .B(input_s2[50]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_2_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_2_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_2_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[50]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_3_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[3]), .B(input_s2[51]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_3_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_3_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_3_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[51]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_4_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[4]), .B(input_s2[36]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_4_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_4_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_4_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[36]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_5_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[5]), .B(input_s2[37]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_5_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_5_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_5_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[37]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_6_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[6]), .B(input_s2[38]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_6_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_6_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_6_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[38]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_7_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[7]), .B(input_s2[39]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_7_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_7_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_7_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[39]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_8_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[8]), .B(input_s2[24]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_8_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_8_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_8_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[24]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_9_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[9]), .B(input_s2[25]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_9_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_9_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_9_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[25]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_10_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[10]), .B(input_s2[26]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_10_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_10_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_10_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[26]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_11_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[11]), .B(input_s2[27]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_11_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_11_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_11_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[27]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_12_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[12]), .B(input_s2[12]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_12_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_12_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_12_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[12]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_13_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[13]), .B(input_s2[13]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_13_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_13_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_13_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[13]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_14_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[14]), .B(input_s2[14]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_14_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_14_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_14_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[14]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_15_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[15]), .B(input_s2[15]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_15_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_15_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_15_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[15]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_16_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[16]), .B(input_s2[0]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_16_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_16_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_16_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[0]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_17_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[17]), .B(input_s2[1]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_17_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_17_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_17_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[1]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_18_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[18]), .B(input_s2[2]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_18_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_18_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_18_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[2]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_19_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[19]), .B(input_s2[3]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_19_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_19_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_19_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[3]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_20_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[20]), .B(input_s2[52]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_20_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_20_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_20_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[52]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_21_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[21]), .B(input_s2[53]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_21_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_21_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_21_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[53]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_22_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[22]), .B(input_s2[54]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_22_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_22_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_22_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[54]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_23_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[23]), .B(input_s2[55]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_23_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_23_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_23_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[55]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_24_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[24]), .B(input_s2[40]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_24_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_24_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_24_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[40]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_25_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[25]), .B(input_s2[41]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_25_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_25_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_25_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[41]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_26_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[26]), .B(input_s2[42]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_26_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_26_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_26_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[42]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_27_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[27]), .B(input_s2[43]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_27_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_27_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_27_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[43]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_28_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[28]), .B(input_s2[28]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_28_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_28_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_28_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[28]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_29_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[29]), .B(input_s2[29]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_29_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_29_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_29_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[29]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_30_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[30]), .B(input_s2[30]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_30_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_30_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_30_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[30]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_31_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[31]), .B(input_s2[31]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_31_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_31_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_31_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[31]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_32_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[32]), .B(input_s2[16]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_32_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_32_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_32_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[16]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_33_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[33]), .B(input_s2[17]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_33_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_33_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_33_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[17]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_34_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[34]), .B(input_s2[18]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_34_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_34_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_34_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[18]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_35_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[35]), .B(input_s2[19]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_35_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_35_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_35_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[19]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_36_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[36]), .B(input_s2[4]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_36_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_36_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_36_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[4]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_37_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[37]), .B(input_s2[5]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_37_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_37_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_37_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[5]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_38_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[38]), .B(input_s2[6]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_38_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_38_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_38_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[6]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_39_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[39]), .B(input_s2[7]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_39_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_39_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_39_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[7]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_40_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[40]), .B(input_s2[56]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_40_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_40_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_40_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[56]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_41_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[41]), .B(input_s2[57]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_41_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_41_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_41_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[57]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_42_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[42]), .B(input_s2[58]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_42_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_42_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_42_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[58]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_43_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[43]), .B(input_s2[59]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_43_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_43_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_43_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[59]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_44_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[44]), .B(input_s2[44]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_44_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_44_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_44_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[44]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_45_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[45]), .B(input_s2[45]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_45_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_45_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_45_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[45]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_46_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[46]), .B(input_s2[46]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_46_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_46_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_46_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[46]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_47_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[47]), .B(input_s2[47]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_47_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_47_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_47_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[47]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_48_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[48]), .B(input_s2[32]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_48_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_48_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_48_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[32]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_49_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[49]), .B(input_s2[33]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_49_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_49_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_49_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[33]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_50_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[50]), .B(input_s2[34]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_50_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_50_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_50_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[34]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_51_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[51]), .B(input_s2[35]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_51_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_51_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_51_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[35]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_52_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[52]), .B(input_s2[20]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_52_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_52_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_52_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[20]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_53_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[53]), .B(input_s2[21]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_53_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_53_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_53_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[21]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_54_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[54]), .B(input_s2[22]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_54_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_54_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_54_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[22]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_55_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[55]), .B(input_s2[23]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_55_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_55_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_55_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[23]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_56_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[56]), .B(input_s2[8]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_56_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_56_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_56_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[8]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_57_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[57]), .B(input_s2[9]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_57_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_57_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_57_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[9]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_58_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[58]), .B(input_s2[10]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_58_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_58_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_58_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[10]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_59_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[59]), .B(input_s2[11]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_59_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_59_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_59_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[11]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_60_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[60]), .B(input_s2[60]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_60_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_60_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_60_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[60]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_61_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[61]), .B(input_s2[61]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_61_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_61_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_61_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[61]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_62_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[62]), .B(input_s2[62]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_62_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_62_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_62_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[62]) , .QN());
  MUX2_X1 prince_rounds_roundResult_Reg_s2_SFF_63_SFFInst_U3 ( .A(
        prince_rounds_mul_result_s2[63]), .B(input_s2[63]), .S(rst), .Z(
        prince_rounds_roundResult_Reg_s2_SFF_63_SFFInst_N3) );
  DFF_X1 prince_rounds_roundResult_Reg_s2_SFF_63_SFFInst_Q_reg ( .D(
        prince_rounds_roundResult_Reg_s2_SFF_63_SFFInst_N3), .CK(clk), .Q(
        prince_rounds_SR_Result_s2[63]) , .QN());
  INV_X1 prince_rounds_MUX_inst0_U4 ( .A(roundHalf_Select_Signal), .ZN(
        prince_rounds_MUX_inst0_n11) );
  INV_X1 prince_rounds_MUX_inst0_U3 ( .A(prince_rounds_MUX_inst0_n11), .ZN(
        prince_rounds_MUX_inst0_n8) );
  INV_X1 prince_rounds_MUX_inst0_U2 ( .A(prince_rounds_MUX_inst0_n11), .ZN(
        prince_rounds_MUX_inst0_n9) );
  INV_X2 prince_rounds_MUX_inst0_U1 ( .A(prince_rounds_MUX_inst0_n11), .ZN(
        prince_rounds_MUX_inst0_n10) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_0_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[0]), .B(
        prince_rounds_SR_Result_s1[48]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[0]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[1]), .B(
        prince_rounds_SR_Result_s1[49]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[1]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[2]), .B(
        prince_rounds_SR_Result_s1[50]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[2]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[3]), .B(
        prince_rounds_SR_Result_s1[51]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[3]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_4_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[4]), .B(
        prince_rounds_SR_Result_s1[36]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[4]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_5_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[5]), .B(
        prince_rounds_SR_Result_s1[37]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[5]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_6_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[6]), .B(
        prince_rounds_SR_Result_s1[38]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[6]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_7_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[7]), .B(
        prince_rounds_SR_Result_s1[39]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[7]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_8_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[8]), .B(
        prince_rounds_SR_Result_s1[24]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[8]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_9_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[9]), .B(
        prince_rounds_SR_Result_s1[25]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[9]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_10_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[10]), .B(
        prince_rounds_SR_Result_s1[26]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[10]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_11_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[11]), .B(
        prince_rounds_SR_Result_s1[27]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[11]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_12_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[12]), .B(
        prince_rounds_SR_Result_s1[12]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[12]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_13_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[13]), .B(
        prince_rounds_SR_Result_s1[13]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[13]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_14_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[14]), .B(
        prince_rounds_SR_Result_s1[14]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[14]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_15_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[15]), .B(
        prince_rounds_SR_Result_s1[15]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[15]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_16_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[16]), .B(
        prince_rounds_SR_Result_s1[0]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[16]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_17_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[17]), .B(
        prince_rounds_SR_Result_s1[1]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[17]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_18_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[18]), .B(
        prince_rounds_SR_Result_s1[2]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[18]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_19_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[19]), .B(
        prince_rounds_SR_Result_s1[3]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[19]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_20_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[20]), .B(
        prince_rounds_SR_Result_s1[52]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[20]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_21_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[21]), .B(
        prince_rounds_SR_Result_s1[53]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[21]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_22_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[22]), .B(
        prince_rounds_SR_Result_s1[54]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[22]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_23_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[23]), .B(
        prince_rounds_SR_Result_s1[55]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[23]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_24_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[24]), .B(
        prince_rounds_SR_Result_s1[40]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[24]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_25_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[25]), .B(
        prince_rounds_SR_Result_s1[41]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[25]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_26_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[26]), .B(
        prince_rounds_SR_Result_s1[42]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[26]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_27_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[27]), .B(
        prince_rounds_SR_Result_s1[43]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[27]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_28_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[28]), .B(
        prince_rounds_SR_Result_s1[28]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[28]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_29_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[29]), .B(
        prince_rounds_SR_Result_s1[29]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[29]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_30_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[30]), .B(
        prince_rounds_SR_Result_s1[30]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[30]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_31_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[31]), .B(
        prince_rounds_SR_Result_s1[31]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[31]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_32_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[32]), .B(
        prince_rounds_SR_Result_s1[16]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[32]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_33_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[33]), .B(
        prince_rounds_SR_Result_s1[17]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[33]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_34_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[34]), .B(
        prince_rounds_SR_Result_s1[18]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[34]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_35_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[35]), .B(
        prince_rounds_SR_Result_s1[19]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[35]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_36_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[36]), .B(
        prince_rounds_SR_Result_s1[4]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[36]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_37_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[37]), .B(
        prince_rounds_SR_Result_s1[5]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[37]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_38_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[38]), .B(
        prince_rounds_SR_Result_s1[6]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[38]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_39_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[39]), .B(
        prince_rounds_SR_Result_s1[7]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[39]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_40_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[40]), .B(
        prince_rounds_SR_Result_s1[56]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[40]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_41_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[41]), .B(
        prince_rounds_SR_Result_s1[57]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[41]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_42_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[42]), .B(
        prince_rounds_SR_Result_s1[58]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[42]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_43_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[43]), .B(
        prince_rounds_SR_Result_s1[59]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[43]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_44_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[44]), .B(
        prince_rounds_SR_Result_s1[44]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[44]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_45_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[45]), .B(
        prince_rounds_SR_Result_s1[45]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[45]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_46_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[46]), .B(
        prince_rounds_SR_Result_s1[46]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[46]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_47_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[47]), .B(
        prince_rounds_SR_Result_s1[47]), .S(prince_rounds_MUX_inst0_n9), .Z(
        prince_rounds_Sbox_Input_s1[47]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_48_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[48]), .B(
        prince_rounds_SR_Result_s1[32]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[48]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_49_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[49]), .B(
        prince_rounds_SR_Result_s1[33]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[49]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_50_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[50]), .B(
        prince_rounds_SR_Result_s1[34]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[50]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_51_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[51]), .B(
        prince_rounds_SR_Result_s1[35]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[51]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_52_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[52]), .B(
        prince_rounds_SR_Result_s1[20]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[52]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_53_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[53]), .B(
        prince_rounds_SR_Result_s1[21]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[53]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_54_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[54]), .B(
        prince_rounds_SR_Result_s1[22]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[54]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_55_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[55]), .B(
        prince_rounds_SR_Result_s1[23]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[55]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_56_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[56]), .B(
        prince_rounds_SR_Result_s1[8]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[56]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_57_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[57]), .B(
        prince_rounds_SR_Result_s1[9]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[57]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_58_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[58]), .B(
        prince_rounds_SR_Result_s1[10]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[58]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_59_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[59]), .B(
        prince_rounds_SR_Result_s1[11]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[59]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_60_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[60]), .B(
        prince_rounds_SR_Result_s1[60]), .S(prince_rounds_MUX_inst0_n8), .Z(
        prince_rounds_Sbox_Input_s1[60]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_61_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[61]), .B(
        prince_rounds_SR_Result_s1[61]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[61]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_62_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[62]), .B(
        prince_rounds_SR_Result_s1[62]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[62]) );
  MUX2_X1 prince_rounds_MUX_inst0_MUXInst_63_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[63]), .B(
        prince_rounds_SR_Result_s1[63]), .S(prince_rounds_MUX_inst0_n10), .Z(
        prince_rounds_Sbox_Input_s1[63]) );
  INV_X1 prince_rounds_MUX_inst1_U5 ( .A(roundHalf_Select_Signal), .ZN(
        prince_rounds_MUX_inst1_n12) );
  INV_X1 prince_rounds_MUX_inst1_U4 ( .A(prince_rounds_MUX_inst1_n12), .ZN(
        prince_rounds_MUX_inst1_n9) );
  INV_X1 prince_rounds_MUX_inst1_U3 ( .A(prince_rounds_MUX_inst1_n12), .ZN(
        prince_rounds_MUX_inst1_n10) );
  INV_X1 prince_rounds_MUX_inst1_U2 ( .A(prince_rounds_MUX_inst1_n12), .ZN(
        prince_rounds_MUX_inst1_n11) );
  INV_X1 prince_rounds_MUX_inst1_U1 ( .A(prince_rounds_MUX_inst1_n12), .ZN(
        prince_rounds_MUX_inst1_n8) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_0_U1 ( .A(
        prince_rounds_SR_Result_s2[0]), .B(prince_rounds_SR_Result_s2[48]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[0]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_1_U1 ( .A(
        prince_rounds_SR_Result_s2[1]), .B(prince_rounds_SR_Result_s2[49]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[1]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_2_U1 ( .A(
        prince_rounds_SR_Result_s2[2]), .B(prince_rounds_SR_Result_s2[50]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[2]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_3_U1 ( .A(
        prince_rounds_SR_Result_s2[3]), .B(prince_rounds_SR_Result_s2[51]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[3]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_4_U1 ( .A(
        prince_rounds_SR_Result_s2[4]), .B(prince_rounds_SR_Result_s2[36]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[4]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_5_U1 ( .A(
        prince_rounds_SR_Result_s2[5]), .B(prince_rounds_SR_Result_s2[37]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[5]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_6_U1 ( .A(
        prince_rounds_SR_Result_s2[6]), .B(prince_rounds_SR_Result_s2[38]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[6]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_7_U1 ( .A(
        prince_rounds_SR_Result_s2[7]), .B(prince_rounds_SR_Result_s2[39]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[7]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_8_U1 ( .A(
        prince_rounds_SR_Result_s2[8]), .B(prince_rounds_SR_Result_s2[24]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[8]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_9_U1 ( .A(
        prince_rounds_SR_Result_s2[9]), .B(prince_rounds_SR_Result_s2[25]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[9]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_10_U1 ( .A(
        prince_rounds_SR_Result_s2[10]), .B(prince_rounds_SR_Result_s2[26]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[10]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_11_U1 ( .A(
        prince_rounds_SR_Result_s2[11]), .B(prince_rounds_SR_Result_s2[27]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[11]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_12_U1 ( .A(
        prince_rounds_SR_Result_s2[12]), .B(prince_rounds_SR_Result_s2[12]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[12]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_13_U1 ( .A(
        prince_rounds_SR_Result_s2[13]), .B(prince_rounds_SR_Result_s2[13]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[13]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_14_U1 ( .A(
        prince_rounds_SR_Result_s2[14]), .B(prince_rounds_SR_Result_s2[14]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[14]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_15_U1 ( .A(
        prince_rounds_SR_Result_s2[15]), .B(prince_rounds_SR_Result_s2[15]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[15]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_16_U1 ( .A(
        prince_rounds_SR_Result_s2[16]), .B(prince_rounds_SR_Result_s2[0]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[16]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_17_U1 ( .A(
        prince_rounds_SR_Result_s2[17]), .B(prince_rounds_SR_Result_s2[1]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[17]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_18_U1 ( .A(
        prince_rounds_SR_Result_s2[18]), .B(prince_rounds_SR_Result_s2[2]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[18]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_19_U1 ( .A(
        prince_rounds_SR_Result_s2[19]), .B(prince_rounds_SR_Result_s2[3]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[19]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_20_U1 ( .A(
        prince_rounds_SR_Result_s2[20]), .B(prince_rounds_SR_Result_s2[52]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[20]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_21_U1 ( .A(
        prince_rounds_SR_Result_s2[21]), .B(prince_rounds_SR_Result_s2[53]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[21]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_22_U1 ( .A(
        prince_rounds_SR_Result_s2[22]), .B(prince_rounds_SR_Result_s2[54]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[22]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_23_U1 ( .A(
        prince_rounds_SR_Result_s2[23]), .B(prince_rounds_SR_Result_s2[55]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[23]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_24_U1 ( .A(
        prince_rounds_SR_Result_s2[24]), .B(prince_rounds_SR_Result_s2[40]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[24])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_25_U1 ( .A(
        prince_rounds_SR_Result_s2[25]), .B(prince_rounds_SR_Result_s2[41]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[25])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_26_U1 ( .A(
        prince_rounds_SR_Result_s2[26]), .B(prince_rounds_SR_Result_s2[42]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[26])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_27_U1 ( .A(
        prince_rounds_SR_Result_s2[27]), .B(prince_rounds_SR_Result_s2[43]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[27])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_28_U1 ( .A(
        prince_rounds_SR_Result_s2[28]), .B(prince_rounds_SR_Result_s2[28]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[28])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_29_U1 ( .A(
        prince_rounds_SR_Result_s2[29]), .B(prince_rounds_SR_Result_s2[29]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[29])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_30_U1 ( .A(
        prince_rounds_SR_Result_s2[30]), .B(prince_rounds_SR_Result_s2[30]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[30])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_31_U1 ( .A(
        prince_rounds_SR_Result_s2[31]), .B(prince_rounds_SR_Result_s2[31]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[31])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_32_U1 ( .A(
        prince_rounds_SR_Result_s2[32]), .B(prince_rounds_SR_Result_s2[16]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[32])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_33_U1 ( .A(
        prince_rounds_SR_Result_s2[33]), .B(prince_rounds_SR_Result_s2[17]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[33])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_34_U1 ( .A(
        prince_rounds_SR_Result_s2[34]), .B(prince_rounds_SR_Result_s2[18]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[34])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_35_U1 ( .A(
        prince_rounds_SR_Result_s2[35]), .B(prince_rounds_SR_Result_s2[19]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[35])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_36_U1 ( .A(
        prince_rounds_SR_Result_s2[36]), .B(prince_rounds_SR_Result_s2[4]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[36]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_37_U1 ( .A(
        prince_rounds_SR_Result_s2[37]), .B(prince_rounds_SR_Result_s2[5]), 
        .S(prince_rounds_MUX_inst1_n8), .Z(prince_rounds_Sbox_Input_s2[37]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_38_U1 ( .A(
        prince_rounds_SR_Result_s2[38]), .B(prince_rounds_SR_Result_s2[6]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[38]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_39_U1 ( .A(
        prince_rounds_SR_Result_s2[39]), .B(prince_rounds_SR_Result_s2[7]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[39]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_40_U1 ( .A(
        prince_rounds_SR_Result_s2[40]), .B(prince_rounds_SR_Result_s2[56]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[40])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_41_U1 ( .A(
        prince_rounds_SR_Result_s2[41]), .B(prince_rounds_SR_Result_s2[57]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[41])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_42_U1 ( .A(
        prince_rounds_SR_Result_s2[42]), .B(prince_rounds_SR_Result_s2[58]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[42])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_43_U1 ( .A(
        prince_rounds_SR_Result_s2[43]), .B(prince_rounds_SR_Result_s2[59]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[43])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_44_U1 ( .A(
        prince_rounds_SR_Result_s2[44]), .B(prince_rounds_SR_Result_s2[44]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[44])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_45_U1 ( .A(
        prince_rounds_SR_Result_s2[45]), .B(prince_rounds_SR_Result_s2[45]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[45]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_46_U1 ( .A(
        prince_rounds_SR_Result_s2[46]), .B(prince_rounds_SR_Result_s2[46]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[46])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_47_U1 ( .A(
        prince_rounds_SR_Result_s2[47]), .B(prince_rounds_SR_Result_s2[47]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[47]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_48_U1 ( .A(
        prince_rounds_SR_Result_s2[48]), .B(prince_rounds_SR_Result_s2[32]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[48])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_49_U1 ( .A(
        prince_rounds_SR_Result_s2[49]), .B(prince_rounds_SR_Result_s2[33]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[49])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_50_U1 ( .A(
        prince_rounds_SR_Result_s2[50]), .B(prince_rounds_SR_Result_s2[34]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[50])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_51_U1 ( .A(
        prince_rounds_SR_Result_s2[51]), .B(prince_rounds_SR_Result_s2[35]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[51])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_52_U1 ( .A(
        prince_rounds_SR_Result_s2[52]), .B(prince_rounds_SR_Result_s2[20]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[52])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_53_U1 ( .A(
        prince_rounds_SR_Result_s2[53]), .B(prince_rounds_SR_Result_s2[21]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[53])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_54_U1 ( .A(
        prince_rounds_SR_Result_s2[54]), .B(prince_rounds_SR_Result_s2[22]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[54])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_55_U1 ( .A(
        prince_rounds_SR_Result_s2[55]), .B(prince_rounds_SR_Result_s2[23]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[55])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_56_U1 ( .A(
        prince_rounds_SR_Result_s2[56]), .B(prince_rounds_SR_Result_s2[8]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[56])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_57_U1 ( .A(
        prince_rounds_SR_Result_s2[57]), .B(prince_rounds_SR_Result_s2[9]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[57])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_58_U1 ( .A(
        prince_rounds_SR_Result_s2[58]), .B(prince_rounds_SR_Result_s2[10]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[58])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_59_U1 ( .A(
        prince_rounds_SR_Result_s2[59]), .B(prince_rounds_SR_Result_s2[11]), 
        .S(prince_rounds_MUX_inst1_n11), .Z(prince_rounds_Sbox_Input_s2[59])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_60_U1 ( .A(
        prince_rounds_SR_Result_s2[60]), .B(prince_rounds_SR_Result_s2[60]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[60]) );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_61_U1 ( .A(
        prince_rounds_SR_Result_s2[61]), .B(prince_rounds_SR_Result_s2[61]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[61])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_62_U1 ( .A(
        prince_rounds_SR_Result_s2[62]), .B(prince_rounds_SR_Result_s2[62]), 
        .S(prince_rounds_MUX_inst1_n10), .Z(prince_rounds_Sbox_Input_s2[62])
         );
  MUX2_X1 prince_rounds_MUX_inst1_MUXInst_63_U1 ( .A(
        prince_rounds_SR_Result_s2[63]), .B(prince_rounds_SR_Result_s2[63]), 
        .S(prince_rounds_MUX_inst1_n9), .Z(prince_rounds_Sbox_Input_s2[63]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n53), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n52), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n53) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U30 ( .A(
        prince_rounds_Sbox_Input_s1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n52) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n49), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n48), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n47), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n46), .S(
        prince_rounds_Sbox_Input_s1[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n49) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n45), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n46) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n44), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n45) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n43), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n42), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n41), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n43) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U23 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n41) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n40), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n42) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n39), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n38), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n37), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n44), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n38) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n47), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n51), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n39) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n36), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n35), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U17 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n34), .B(
        prince_rounds_Sbox_Input_s1[0]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n44), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n35) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n47), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n36) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n37), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n47) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n33), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n37), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n40), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n33) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n44), .A2(
        prince_rounds_Sbox_Input_s1[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n40) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n32), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n31), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n34), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n31) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n37), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n48), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n32) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n30), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n48), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n44), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n48) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U6 ( .A(
        prince_rounds_Sbox_Input_s1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n44) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n34), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n50) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s2[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n34) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n37), .B(
        prince_rounds_Sbox_Input_s1[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n30) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n51) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F1_n37) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n28), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n27), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n26), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n27) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(prince_rounds_Sbox_Input_s1[3]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n26) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n24), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n28) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n23), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n22), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n22) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n21), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n20), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n23) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(prince_rounds_Sbox_Input_s1[1]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n20) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n18), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n19) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n17) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n14), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n18) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n14) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n13), .S(
        prince_rounds_Sbox_Input_s1[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n13) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n12), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n11), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n21), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n10), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n11) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(prince_rounds_Sbox_Input_s1[1]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n12) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n9), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n8), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n8) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n7), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n9) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n10), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n5), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n5) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n16), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n10) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n4), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n7), .A2(
        prince_rounds_Sbox_Input_s1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n3) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n7) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n24), .A2(
        prince_rounds_Sbox_Input_s1[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n21) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n15), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n25), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n4) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n16), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n25) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n16) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n24), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n15) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F2_n24) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n29), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n28), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n27), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n26), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n29) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n25), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n24), .S(
        prince_rounds_Sbox_Input_s1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n23), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n22), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n24) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n28), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n22) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n25) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n20), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n28), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n19) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n28) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n18), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n27), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n20) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n26), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n18) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n26) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n14), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n13), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n15) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n27), .B(
        prince_rounds_Sbox_Input_s1[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n14) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n12), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n11), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n10), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n11) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n27), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n16), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n10) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n12) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(prince_rounds_Sbox_Input_s1[3]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[0]), .B(prince_rounds_Sbox_Input_s1[3]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n9), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(prince_rounds_Sbox_Input_s1[2]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n9) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n8), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n7), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n27), .A2(
        prince_rounds_Sbox_Input_s1[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n7) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n27) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n23), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n8) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(prince_rounds_Sbox_Input_s1[0]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n21) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(prince_rounds_Sbox_Input_s1[0]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n23) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n13), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n16), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n16) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n13) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(prince_rounds_Sbox_Input_s1[2]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F3_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U37 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n32), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n31), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U36 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n31) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U35 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n29), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n32) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n28), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n27), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n26), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n25), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n27) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n24), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n23), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n28) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n22), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n29), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n21) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n26), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n20), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n22) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n24), .B(
        prince_rounds_Sbox_Input_s2[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n23), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n20) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(prince_rounds_Sbox_Input_s2[2]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n23) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n24) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n18), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n26) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n14), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n15) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n14) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n13), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n29), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n16) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n12), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n11), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n18), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n11) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U18 ( .A(
        prince_rounds_Sbox_Input_s2[3]), .B(prince_rounds_Sbox_Input_s2[2]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n12) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n10), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n9), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n13), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n10) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n8), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n13) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n18), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n7), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n7) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n17), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n9), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U11 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n5), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n9) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U10 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n17) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n18) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n8), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n4), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n29), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n4) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n30) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n19) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n25), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n29) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n25) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n5), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n8) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F4_n5) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[3]), .B(prince_rounds_Sbox_Input_s2[0]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n32), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n31), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n32) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n29), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n28), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n27), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n29) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n26), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n31), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n28) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n24), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n23), .B(
        prince_rounds_Sbox_Input_s2[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n25) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n22), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n26), .A2(
        prince_rounds_Sbox_Input_s1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n23), .B(
        prince_rounds_Sbox_Input_s1[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n22) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n20), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n19), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n20) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n30), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n18) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n14), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n27), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n13), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n24), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n23), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n16) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n31), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n24) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n19), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n12), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n13) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n11), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n10), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n14), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n9), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n11) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n23), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n8), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n9) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n7), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n8) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n26), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n27), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n7) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n14) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n12), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n23), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n5), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n10), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n26), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n10) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n31), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n27), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n19) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n27) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n31) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n23) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n30) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n17), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n26), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n12) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n26) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(prince_rounds_Sbox_Input_s1[3]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F5_n17) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n31), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n30), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n29), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n28), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n30) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n27), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n26), .S(
        prince_rounds_Sbox_Input_s2[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n31) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n25), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n27) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n24), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n23), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n29), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n22), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n23) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n22) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n20), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n19), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n18), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n24), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n17), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n19) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n16), .A2(
        prince_rounds_Sbox_Input_s2[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n20) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n15), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n14), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n13), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n14) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n12), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n11), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n15) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n11) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n10), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n16), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n12), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n9), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n10) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n8), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n9) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n26), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n12) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[0]), .A2(prince_rounds_Sbox_Input_s2[3]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n26) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n7), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n8), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n7) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[0]), .A2(prince_rounds_Sbox_Input_s2[3]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n25) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n6), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n5), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n28), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n5) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n4), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n16), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n24), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n8), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n4) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n29), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n8) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(prince_rounds_Sbox_Input_s1[1]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n29) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n16) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n3), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n21) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n17) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n2), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n1), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n28), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n13), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n1) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n24), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n13) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n28) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n24), .A2(
        prince_rounds_Sbox_Input_s2[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n18) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n24) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n2) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F6_n3) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n57), .A2(
        prince_rounds_Sbox_Input_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n55), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n54), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n53), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n52), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n54) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n52) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n55), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n50), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n49), .A2(
        prince_rounds_Sbox_Input_s2[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n50) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n48), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n47), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n49) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n46), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n48) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n45), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n55) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n44), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n45) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(prince_rounds_Sbox_Input_s2[3]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n44) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n47), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n43), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n57), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n42), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n43) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(prince_rounds_Sbox_Input_s1[2]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n42) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n41), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n47) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n40), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n39), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n39) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n41), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n40) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n57) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(prince_rounds_Sbox_Input_s1[2]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n41) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n38), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n37), .A2(
        prince_rounds_Sbox_Input_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n38) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[2]), .B(prince_rounds_Sbox_Input_s2[3]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n37) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n36), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n53), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n46), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n53) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n46) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51), .B(
        prince_rounds_Sbox_Input_s1[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n36) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n51) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n35), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n56), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n35) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(prince_rounds_Sbox_Input_s2[0]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F7_n56) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n30), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n29), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n28), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n29) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n27), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n26), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n30) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n25), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n24), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n27) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n23), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n22), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n21), .A2(
        prince_rounds_Sbox_Input_s2[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n22) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20), .B(
        prince_rounds_Sbox_Input_s1[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n23) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n19), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n18), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n19) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n17) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n21), .A2(
        prince_rounds_Sbox_Input_s2[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n15) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n14), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n18) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n24), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n13), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n28), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n26), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n13) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[0]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n12), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n26) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n28) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n12), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n11), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n24), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n25), .S(
        prince_rounds_Sbox_Input_s2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n11) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n16), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n25) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n14), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n24) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n12) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n10), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n9), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n16), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n9) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n14), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n16) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n14) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n8), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n7), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n10) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n7), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[2]), .B(prince_rounds_Sbox_Input_s1[3]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n7) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n5), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n4), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[3]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n4) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n2), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n3) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20), .A2(
        prince_rounds_Sbox_Input_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n2) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n8), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n1), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n5) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[1]), .A2(prince_rounds_Sbox_Input_s2[2]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n1) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n21), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n8) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n21) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_N_F8_n20) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_n2), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_n1), .ZN(
        prince_rounds_sub_Inv_Result_s1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_n1) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst1_n2) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_n5), .ZN(
        output_s2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_n5), .ZN(
        output_s2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_n5), .ZN(
        output_s2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_n5), .ZN(
        output_s2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n79) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U30 ( .A(
        prince_rounds_Sbox_Input_s1[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U23 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n77), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U17 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n66), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n57) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U6 ( .A(
        prince_rounds_Sbox_Input_s1[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n70) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s2[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n60) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(prince_rounds_Sbox_Input_s1[7]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(prince_rounds_Sbox_Input_s1[5]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(prince_rounds_Sbox_Input_s1[5]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(prince_rounds_Sbox_Input_s1[7]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[4]), .B(prince_rounds_Sbox_Input_s1[7]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(prince_rounds_Sbox_Input_s1[6]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(prince_rounds_Sbox_Input_s1[4]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(prince_rounds_Sbox_Input_s1[4]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(prince_rounds_Sbox_Input_s1[6]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U37 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U36 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U35 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n74) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n76), .B(
        prince_rounds_Sbox_Input_s2[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n75), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(prince_rounds_Sbox_Input_s2[6]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U18 ( .A(
        prince_rounds_Sbox_Input_s2[7]), .B(prince_rounds_Sbox_Input_s2[6]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U11 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U10 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[7]), .B(prince_rounds_Sbox_Input_s2[4]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(prince_rounds_Sbox_Input_s1[7]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[4]), .A2(prince_rounds_Sbox_Input_s2[7]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[4]), .A2(prince_rounds_Sbox_Input_s2[7]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(prince_rounds_Sbox_Input_s1[5]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(prince_rounds_Sbox_Input_s2[7]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(prince_rounds_Sbox_Input_s1[6]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(prince_rounds_Sbox_Input_s1[6]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[6]), .B(prince_rounds_Sbox_Input_s2[7]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(prince_rounds_Sbox_Input_s2[4]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n88) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86), .B(
        prince_rounds_Sbox_Input_s1[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[4]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[6]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[6]), .B(prince_rounds_Sbox_Input_s1[7]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[7]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[6]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86), .A2(
        prince_rounds_Sbox_Input_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[5]), .A2(prince_rounds_Sbox_Input_s2[6]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n87) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_N_F8_n86) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[4]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_n5), .ZN(
        output_s2[4]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_n5), .ZN(
        output_s2[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[6]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_n5), .ZN(
        output_s2[6]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[7]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_n5), .ZN(
        output_s2[7]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[8]), .B(prince_rounds_Sbox_Input_s2[11]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(prince_rounds_Sbox_Input_s1[11]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(prince_rounds_Sbox_Input_s1[9]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(prince_rounds_Sbox_Input_s1[9]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[10]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[10]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(prince_rounds_Sbox_Input_s1[11]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[8]), .B(prince_rounds_Sbox_Input_s1[11]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(prince_rounds_Sbox_Input_s1[10]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(prince_rounds_Sbox_Input_s1[8]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(prince_rounds_Sbox_Input_s1[8]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[11]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(prince_rounds_Sbox_Input_s1[10]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[9]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[11]), .B(prince_rounds_Sbox_Input_s2[8]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(prince_rounds_Sbox_Input_s1[11]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[8]), .A2(prince_rounds_Sbox_Input_s2[11]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[8]), .A2(prince_rounds_Sbox_Input_s2[11]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(prince_rounds_Sbox_Input_s1[9]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(prince_rounds_Sbox_Input_s2[11]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(prince_rounds_Sbox_Input_s1[10]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(prince_rounds_Sbox_Input_s1[10]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[10]), .B(prince_rounds_Sbox_Input_s2[11]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[11]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(prince_rounds_Sbox_Input_s2[8]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[8]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[10]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[10]), .B(prince_rounds_Sbox_Input_s1[11]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[11]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[10]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[9]), .A2(prince_rounds_Sbox_Input_s2[10]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[8]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_n5), .ZN(
        output_s2[8]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[9]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_n5), .ZN(
        output_s2[9]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[10]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_n5), .ZN(
        output_s2[10]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[11]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_n5), .ZN(
        output_s2[11]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[12]), .B(prince_rounds_Sbox_Input_s2[15]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[12]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(prince_rounds_Sbox_Input_s1[15]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(prince_rounds_Sbox_Input_s1[13]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[12]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(prince_rounds_Sbox_Input_s1[13]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[14]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[14]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(prince_rounds_Sbox_Input_s1[15]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[12]), .B(prince_rounds_Sbox_Input_s1[15]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(prince_rounds_Sbox_Input_s1[14]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(prince_rounds_Sbox_Input_s1[12]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(prince_rounds_Sbox_Input_s1[12]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[15]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(prince_rounds_Sbox_Input_s1[14]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[13]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[15]), .B(prince_rounds_Sbox_Input_s2[12]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(prince_rounds_Sbox_Input_s1[15]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[12]), .A2(prince_rounds_Sbox_Input_s2[15]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[12]), .A2(prince_rounds_Sbox_Input_s2[15]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(prince_rounds_Sbox_Input_s1[13]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(prince_rounds_Sbox_Input_s2[15]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(prince_rounds_Sbox_Input_s1[14]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(prince_rounds_Sbox_Input_s1[14]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[14]), .B(prince_rounds_Sbox_Input_s2[15]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[15]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(prince_rounds_Sbox_Input_s2[12]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[12]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[14]), .B(prince_rounds_Sbox_Input_s1[15]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[15]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[14]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[13]), .A2(prince_rounds_Sbox_Input_s2[14]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[12]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_n5), .ZN(
        output_s2[12]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[13]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_n5), .ZN(
        output_s2[13]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[14]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_n5), .ZN(
        output_s2[14]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[15]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_n5), .ZN(
        output_s2[15]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[16]), .B(prince_rounds_Sbox_Input_s2[19]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[16]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(prince_rounds_Sbox_Input_s1[19]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(prince_rounds_Sbox_Input_s1[17]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[16]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(prince_rounds_Sbox_Input_s1[17]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[18]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[18]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(prince_rounds_Sbox_Input_s1[19]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[16]), .B(prince_rounds_Sbox_Input_s1[19]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(prince_rounds_Sbox_Input_s1[18]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(prince_rounds_Sbox_Input_s1[16]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(prince_rounds_Sbox_Input_s1[16]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[19]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(prince_rounds_Sbox_Input_s1[18]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[17]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[19]), .B(prince_rounds_Sbox_Input_s2[16]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(prince_rounds_Sbox_Input_s1[19]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[16]), .A2(prince_rounds_Sbox_Input_s2[19]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[16]), .A2(prince_rounds_Sbox_Input_s2[19]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(prince_rounds_Sbox_Input_s1[17]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(prince_rounds_Sbox_Input_s2[19]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(prince_rounds_Sbox_Input_s1[18]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(prince_rounds_Sbox_Input_s1[18]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[18]), .B(prince_rounds_Sbox_Input_s2[19]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[19]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(prince_rounds_Sbox_Input_s2[16]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n88) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86), .B(
        prince_rounds_Sbox_Input_s1[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[16]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n94) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n73) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U17 ( .A(
        prince_rounds_Sbox_Input_s2[18]), .B(prince_rounds_Sbox_Input_s1[19]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n72) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U14 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U11 ( .A(
        prince_rounds_Sbox_Input_s1[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[18]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n78) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[19]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[18]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86), .A2(
        prince_rounds_Sbox_Input_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[17]), .A2(prince_rounds_Sbox_Input_s2[18]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n75) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n87) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_N_F8_n86) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[16]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_n5), .ZN(
        output_s2[16]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[17]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_n5), .ZN(
        output_s2[17]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[18]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_n5), .ZN(
        output_s2[18]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[19]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_n5), .ZN(
        output_s2[19]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[20]), .B(prince_rounds_Sbox_Input_s2[23]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[20]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(prince_rounds_Sbox_Input_s1[23]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(prince_rounds_Sbox_Input_s1[21]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[20]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(prince_rounds_Sbox_Input_s1[21]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[22]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[22]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(prince_rounds_Sbox_Input_s1[23]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[20]), .B(prince_rounds_Sbox_Input_s1[23]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(prince_rounds_Sbox_Input_s1[22]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(prince_rounds_Sbox_Input_s1[20]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(prince_rounds_Sbox_Input_s1[20]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[23]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(prince_rounds_Sbox_Input_s1[22]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[21]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[23]), .B(prince_rounds_Sbox_Input_s2[20]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(prince_rounds_Sbox_Input_s1[23]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[20]), .A2(prince_rounds_Sbox_Input_s2[23]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[20]), .A2(prince_rounds_Sbox_Input_s2[23]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(prince_rounds_Sbox_Input_s1[21]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(prince_rounds_Sbox_Input_s2[23]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(prince_rounds_Sbox_Input_s1[22]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(prince_rounds_Sbox_Input_s1[22]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[22]), .B(prince_rounds_Sbox_Input_s2[23]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[23]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(prince_rounds_Sbox_Input_s2[20]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[20]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[22]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[22]), .B(prince_rounds_Sbox_Input_s1[23]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[23]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[22]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[21]), .A2(prince_rounds_Sbox_Input_s2[22]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[20]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_n5), .ZN(
        output_s2[20]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[21]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_n5), .ZN(
        output_s2[21]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[22]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_n5), .ZN(
        output_s2[22]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[23]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_n5), .ZN(
        output_s2[23]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[24]), .B(prince_rounds_Sbox_Input_s2[27]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[24]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(prince_rounds_Sbox_Input_s1[27]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(prince_rounds_Sbox_Input_s1[25]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[24]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(prince_rounds_Sbox_Input_s1[25]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[26]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[26]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(prince_rounds_Sbox_Input_s1[27]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[24]), .B(prince_rounds_Sbox_Input_s1[27]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(prince_rounds_Sbox_Input_s1[26]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(prince_rounds_Sbox_Input_s1[24]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(prince_rounds_Sbox_Input_s1[24]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[27]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(prince_rounds_Sbox_Input_s1[26]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[25]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[27]), .B(prince_rounds_Sbox_Input_s2[24]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(prince_rounds_Sbox_Input_s1[27]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[24]), .A2(prince_rounds_Sbox_Input_s2[27]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[24]), .A2(prince_rounds_Sbox_Input_s2[27]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(prince_rounds_Sbox_Input_s1[25]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(prince_rounds_Sbox_Input_s2[27]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(prince_rounds_Sbox_Input_s1[26]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(prince_rounds_Sbox_Input_s1[26]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[26]), .B(prince_rounds_Sbox_Input_s2[27]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[27]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(prince_rounds_Sbox_Input_s2[24]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n88) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86), .B(
        prince_rounds_Sbox_Input_s1[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[24]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n94) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n73) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U17 ( .A(
        prince_rounds_Sbox_Input_s2[26]), .B(prince_rounds_Sbox_Input_s1[27]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n72) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U14 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U11 ( .A(
        prince_rounds_Sbox_Input_s1[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[26]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n78) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[27]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[26]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86), .A2(
        prince_rounds_Sbox_Input_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[25]), .A2(prince_rounds_Sbox_Input_s2[26]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n75) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n87) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_N_F8_n86) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[24]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_n5), .ZN(
        output_s2[24]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[25]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_n5), .ZN(
        output_s2[25]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[26]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_n5), .ZN(
        output_s2[26]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[27]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_n5), .ZN(
        output_s2[27]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[28]), .B(prince_rounds_Sbox_Input_s2[31]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[28]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(prince_rounds_Sbox_Input_s1[31]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(prince_rounds_Sbox_Input_s1[29]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[28]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(prince_rounds_Sbox_Input_s1[29]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[30]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[30]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(prince_rounds_Sbox_Input_s1[31]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[28]), .B(prince_rounds_Sbox_Input_s1[31]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(prince_rounds_Sbox_Input_s1[30]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(prince_rounds_Sbox_Input_s1[28]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(prince_rounds_Sbox_Input_s1[28]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[31]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(prince_rounds_Sbox_Input_s1[30]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[29]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[31]), .B(prince_rounds_Sbox_Input_s2[28]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(prince_rounds_Sbox_Input_s1[31]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[28]), .A2(prince_rounds_Sbox_Input_s2[31]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[28]), .A2(prince_rounds_Sbox_Input_s2[31]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(prince_rounds_Sbox_Input_s1[29]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(prince_rounds_Sbox_Input_s2[31]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(prince_rounds_Sbox_Input_s1[30]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(prince_rounds_Sbox_Input_s1[30]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[30]), .B(prince_rounds_Sbox_Input_s2[31]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[31]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(prince_rounds_Sbox_Input_s2[28]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n88) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86), .B(
        prince_rounds_Sbox_Input_s1[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[28]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[30]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[30]), .B(prince_rounds_Sbox_Input_s1[31]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[31]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[30]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86), .A2(
        prince_rounds_Sbox_Input_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[29]), .A2(prince_rounds_Sbox_Input_s2[30]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n87) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_N_F8_n86) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[28]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_n5), .ZN(
        output_s2[28]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[29]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_n5), .ZN(
        output_s2[29]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[30]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_n5), .ZN(
        output_s2[30]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[31]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_n5), .ZN(
        output_s2[31]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[32]), .B(prince_rounds_Sbox_Input_s2[35]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[32]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(prince_rounds_Sbox_Input_s1[35]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(prince_rounds_Sbox_Input_s1[33]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[32]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(prince_rounds_Sbox_Input_s1[33]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[34]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[34]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(prince_rounds_Sbox_Input_s1[35]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[32]), .B(prince_rounds_Sbox_Input_s1[35]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(prince_rounds_Sbox_Input_s1[34]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(prince_rounds_Sbox_Input_s1[32]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(prince_rounds_Sbox_Input_s1[32]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[35]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(prince_rounds_Sbox_Input_s1[34]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[33]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[35]), .B(prince_rounds_Sbox_Input_s2[32]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(prince_rounds_Sbox_Input_s1[35]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[32]), .A2(prince_rounds_Sbox_Input_s2[35]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[32]), .A2(prince_rounds_Sbox_Input_s2[35]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(prince_rounds_Sbox_Input_s1[33]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(prince_rounds_Sbox_Input_s2[35]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(prince_rounds_Sbox_Input_s1[34]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(prince_rounds_Sbox_Input_s1[34]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[34]), .B(prince_rounds_Sbox_Input_s2[35]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[35]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(prince_rounds_Sbox_Input_s2[32]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n88) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86), .B(
        prince_rounds_Sbox_Input_s1[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[32]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[34]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[34]), .B(prince_rounds_Sbox_Input_s1[35]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[35]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[34]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86), .A2(
        prince_rounds_Sbox_Input_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[33]), .A2(prince_rounds_Sbox_Input_s2[34]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n87) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_N_F8_n86) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[32]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_n5), .ZN(
        output_s2[32]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[33]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_n5), .ZN(
        output_s2[33]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[34]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_n5), .ZN(
        output_s2[34]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[35]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_n5), .ZN(
        output_s2[35]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n70) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n69) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n65), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n73), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U17 ( .A(
        prince_rounds_Sbox_Input_s1[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n62), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n62) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n68) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n64), .A2(
        prince_rounds_Sbox_Input_s1[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n63), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n64), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n75), .A2(
        prince_rounds_Sbox_Input_s1[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n63) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U5 ( .A(
        prince_rounds_Sbox_Input_s1[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n75) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n64) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U3 ( .A(
        prince_rounds_Sbox_Input_s2[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n80), .B(
        prince_rounds_Sbox_Input_s1[38]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F1_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(prince_rounds_Sbox_Input_s1[39]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(prince_rounds_Sbox_Input_s1[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[36]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[37]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(prince_rounds_Sbox_Input_s1[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[38]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[39]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[38]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[38]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(prince_rounds_Sbox_Input_s1[39]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[36]), .B(prince_rounds_Sbox_Input_s1[39]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(prince_rounds_Sbox_Input_s1[38]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(prince_rounds_Sbox_Input_s1[36]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(prince_rounds_Sbox_Input_s1[36]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[39]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(prince_rounds_Sbox_Input_s1[38]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U37 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U36 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U35 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n74) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n76), .B(
        prince_rounds_Sbox_Input_s2[37]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n75), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(prince_rounds_Sbox_Input_s2[38]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U18 ( .A(
        prince_rounds_Sbox_Input_s2[39]), .B(prince_rounds_Sbox_Input_s2[38]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U11 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U10 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[39]), .B(prince_rounds_Sbox_Input_s2[36]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(prince_rounds_Sbox_Input_s1[39]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[38]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[36]), .A2(prince_rounds_Sbox_Input_s2[39]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[36]), .A2(prince_rounds_Sbox_Input_s2[39]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(prince_rounds_Sbox_Input_s1[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(prince_rounds_Sbox_Input_s2[39]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(prince_rounds_Sbox_Input_s1[38]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(prince_rounds_Sbox_Input_s1[38]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[38]), .B(prince_rounds_Sbox_Input_s2[39]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[39]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(prince_rounds_Sbox_Input_s2[36]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[36]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[36]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[38]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[38]), .B(prince_rounds_Sbox_Input_s1[39]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[39]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[38]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[37]), .A2(prince_rounds_Sbox_Input_s2[38]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_0_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_1_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_2_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_3_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_4_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_5_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_6_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_7_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_8_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_9_SFFInst_N3), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[36]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_n5), .ZN(
        output_s2[36]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[37]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_n5), .ZN(
        output_s2[37]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[38]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_n5), .ZN(
        output_s2[38]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[39]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_n5), .ZN(
        output_s2[39]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n79) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U30 ( .A(
        prince_rounds_Sbox_Input_s1[40]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[42]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U23 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n77), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U17 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[40]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n66), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n57) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U6 ( .A(
        prince_rounds_Sbox_Input_s1[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n70) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s2[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n60) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[42]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(prince_rounds_Sbox_Input_s1[43]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(prince_rounds_Sbox_Input_s1[41]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[40]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[41]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(prince_rounds_Sbox_Input_s1[41]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[42]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[43]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[42]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[42]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(prince_rounds_Sbox_Input_s1[43]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[40]), .B(prince_rounds_Sbox_Input_s1[43]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(prince_rounds_Sbox_Input_s1[42]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(prince_rounds_Sbox_Input_s1[40]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(prince_rounds_Sbox_Input_s1[40]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[43]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(prince_rounds_Sbox_Input_s1[42]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U37 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U36 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U35 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n74) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n76), .B(
        prince_rounds_Sbox_Input_s2[41]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n75), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(prince_rounds_Sbox_Input_s2[42]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U18 ( .A(
        prince_rounds_Sbox_Input_s2[43]), .B(prince_rounds_Sbox_Input_s2[42]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U11 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U10 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[43]), .B(prince_rounds_Sbox_Input_s2[40]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(prince_rounds_Sbox_Input_s1[43]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[42]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[40]), .A2(prince_rounds_Sbox_Input_s2[43]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[40]), .A2(prince_rounds_Sbox_Input_s2[43]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(prince_rounds_Sbox_Input_s1[41]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(prince_rounds_Sbox_Input_s2[43]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(prince_rounds_Sbox_Input_s1[42]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(prince_rounds_Sbox_Input_s1[42]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[42]), .B(prince_rounds_Sbox_Input_s2[43]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[43]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(prince_rounds_Sbox_Input_s2[40]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[40]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[40]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[42]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[42]), .B(prince_rounds_Sbox_Input_s1[43]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[43]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[42]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[41]), .A2(prince_rounds_Sbox_Input_s2[42]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_0_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_1_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_2_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_3_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_4_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_5_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_6_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_7_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_8_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_9_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[40]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_n5), .ZN(
        output_s2[40]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[41]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_n5), .ZN(
        output_s2[41]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[42]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_n5), .ZN(
        output_s2[42]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[43]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_n5), .ZN(
        output_s2[43]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n79) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U30 ( .A(
        prince_rounds_Sbox_Input_s1[44]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[46]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U23 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n77), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U17 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[44]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n66), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n57) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U6 ( .A(
        prince_rounds_Sbox_Input_s1[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n70) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s2[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n60) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[46]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(prince_rounds_Sbox_Input_s1[47]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(prince_rounds_Sbox_Input_s1[45]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[44]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[45]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(prince_rounds_Sbox_Input_s1[45]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[46]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[47]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[46]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[46]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(prince_rounds_Sbox_Input_s1[47]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[44]), .B(prince_rounds_Sbox_Input_s1[47]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(prince_rounds_Sbox_Input_s1[46]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(prince_rounds_Sbox_Input_s1[44]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(prince_rounds_Sbox_Input_s1[44]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[47]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(prince_rounds_Sbox_Input_s1[46]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U37 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U36 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U35 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n74) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n76), .B(
        prince_rounds_Sbox_Input_s2[45]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n75), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(prince_rounds_Sbox_Input_s2[46]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U18 ( .A(
        prince_rounds_Sbox_Input_s2[47]), .B(prince_rounds_Sbox_Input_s2[46]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U11 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U10 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[47]), .B(prince_rounds_Sbox_Input_s2[44]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(prince_rounds_Sbox_Input_s1[47]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[46]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[44]), .A2(prince_rounds_Sbox_Input_s2[47]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[44]), .A2(prince_rounds_Sbox_Input_s2[47]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(prince_rounds_Sbox_Input_s1[45]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(prince_rounds_Sbox_Input_s2[47]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(prince_rounds_Sbox_Input_s1[46]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(prince_rounds_Sbox_Input_s1[46]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[46]), .B(prince_rounds_Sbox_Input_s2[47]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[47]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(prince_rounds_Sbox_Input_s2[44]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[44]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[44]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[46]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[46]), .B(prince_rounds_Sbox_Input_s1[47]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[47]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[46]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[45]), .A2(prince_rounds_Sbox_Input_s2[46]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_0_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_1_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_2_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_3_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_4_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_5_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_6_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_7_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_8_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_9_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[44]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_n5), .ZN(
        output_s2[44]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[45]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_n5), .ZN(
        output_s2[45]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[46]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_n5), .ZN(
        output_s2[46]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[47]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_n5), .ZN(
        output_s2[47]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[48]), .B(prince_rounds_Sbox_Input_s2[51]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[50]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[48]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[51]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[50]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(prince_rounds_Sbox_Input_s1[51]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(prince_rounds_Sbox_Input_s1[49]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[48]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[49]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(prince_rounds_Sbox_Input_s1[49]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[50]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[51]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[50]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[50]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(prince_rounds_Sbox_Input_s1[51]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[48]), .B(prince_rounds_Sbox_Input_s1[51]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(prince_rounds_Sbox_Input_s1[50]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(prince_rounds_Sbox_Input_s1[48]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(prince_rounds_Sbox_Input_s1[48]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[51]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(prince_rounds_Sbox_Input_s1[50]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[49]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[51]), .B(prince_rounds_Sbox_Input_s2[48]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(prince_rounds_Sbox_Input_s1[51]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[50]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[48]), .A2(prince_rounds_Sbox_Input_s2[51]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[48]), .A2(prince_rounds_Sbox_Input_s2[51]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(prince_rounds_Sbox_Input_s1[49]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(prince_rounds_Sbox_Input_s2[51]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(prince_rounds_Sbox_Input_s1[50]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(prince_rounds_Sbox_Input_s1[50]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[50]), .B(prince_rounds_Sbox_Input_s2[51]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[51]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(prince_rounds_Sbox_Input_s2[48]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[48]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[48]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[50]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[50]), .B(prince_rounds_Sbox_Input_s1[51]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[51]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[50]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[49]), .A2(prince_rounds_Sbox_Input_s2[50]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_0_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_1_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_2_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_3_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_4_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_5_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_6_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_7_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_8_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_9_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[48]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_n5), .ZN(
        output_s2[48]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[49]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_n5), .ZN(
        output_s2[49]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[50]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_n5), .ZN(
        output_s2[50]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[51]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_n5), .ZN(
        output_s2[51]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n79) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U30 ( .A(
        prince_rounds_Sbox_Input_s1[52]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[54]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U23 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n77), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U17 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[52]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n66), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n57) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U6 ( .A(
        prince_rounds_Sbox_Input_s1[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n70) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s2[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n60) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[54]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(prince_rounds_Sbox_Input_s1[55]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(prince_rounds_Sbox_Input_s1[53]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[52]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[53]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(prince_rounds_Sbox_Input_s1[53]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[54]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[55]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[54]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[54]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(prince_rounds_Sbox_Input_s1[55]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[52]), .B(prince_rounds_Sbox_Input_s1[55]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(prince_rounds_Sbox_Input_s1[54]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(prince_rounds_Sbox_Input_s1[52]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(prince_rounds_Sbox_Input_s1[52]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[55]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(prince_rounds_Sbox_Input_s1[54]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U37 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U36 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U35 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n74) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n76), .B(
        prince_rounds_Sbox_Input_s2[53]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n75), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(prince_rounds_Sbox_Input_s2[54]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U18 ( .A(
        prince_rounds_Sbox_Input_s2[55]), .B(prince_rounds_Sbox_Input_s2[54]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U11 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U10 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[55]), .B(prince_rounds_Sbox_Input_s2[52]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(prince_rounds_Sbox_Input_s1[55]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[54]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[52]), .A2(prince_rounds_Sbox_Input_s2[55]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[52]), .A2(prince_rounds_Sbox_Input_s2[55]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(prince_rounds_Sbox_Input_s1[53]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(prince_rounds_Sbox_Input_s2[55]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(prince_rounds_Sbox_Input_s1[54]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(prince_rounds_Sbox_Input_s1[54]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[54]), .B(prince_rounds_Sbox_Input_s2[55]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[55]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(prince_rounds_Sbox_Input_s2[52]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n88) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86), .B(
        prince_rounds_Sbox_Input_s1[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n87), .A2(
        prince_rounds_Sbox_Input_s2[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[52]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[52]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[54]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[54]), .B(prince_rounds_Sbox_Input_s1[55]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[55]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[54]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86), .A2(
        prince_rounds_Sbox_Input_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[53]), .A2(prince_rounds_Sbox_Input_s2[54]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n87) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_N_F8_n86) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_0_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_1_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_2_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_3_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_4_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_5_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_6_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_7_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_8_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_9_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[52]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_n5), .ZN(
        output_s2[52]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[53]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_n5), .ZN(
        output_s2[53]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[54]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_n5), .ZN(
        output_s2[54]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[55]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_n5), .ZN(
        output_s2[55]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U31 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n78) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U29 ( .A(
        prince_rounds_Sbox_Input_s1[56]), .B(prince_rounds_Sbox_Input_s2[59]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n77) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n72), .S(
        prince_rounds_Sbox_Input_s1[58]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U24 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n73), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[56]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n73) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U12 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[59]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n70), .A2(
        prince_rounds_Sbox_Input_s1[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U8 ( .A(
        prince_rounds_Sbox_Input_s2[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U5 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U4 ( .A(
        prince_rounds_Sbox_Input_s1[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n63), .B(
        prince_rounds_Sbox_Input_s1[58]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n76) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(prince_rounds_Sbox_Input_s1[59]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U29 ( .A1(
        prince_rounds_Sbox_Input_s1[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(prince_rounds_Sbox_Input_s1[57]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U26 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n71) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U22 ( .A(
        prince_rounds_Sbox_Input_s1[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n67) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U21 ( .A(
        prince_rounds_Sbox_Input_s1[56]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n66), .S(
        prince_rounds_Sbox_Input_s1[57]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[2]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n66) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(prince_rounds_Sbox_Input_s1[57]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n59) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U12 ( .A(
        prince_rounds_Sbox_Input_s1[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n56) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n60) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n77), .A2(
        prince_rounds_Sbox_Input_s1[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U4 ( .A(
        prince_rounds_Sbox_Input_s1[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n69) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F2_n77) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n101), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[58]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n99), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n98), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n97), .S(
        prince_rounds_Sbox_Input_s1[59]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n97) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U23 ( .A(
        prince_rounds_Sbox_Input_s1[58]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n91), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n93) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n91) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n88) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U18 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n100), .B(
        prince_rounds_Sbox_Input_s1[58]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s1[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U14 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U13 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(prince_rounds_Sbox_Input_s1[59]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n90) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[56]), .B(prince_rounds_Sbox_Input_s1[59]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(prince_rounds_Sbox_Input_s1[58]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[3]) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n100), .A2(
        prince_rounds_Sbox_Input_s1[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(prince_rounds_Sbox_Input_s1[56]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n94) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(prince_rounds_Sbox_Input_s1[56]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[59]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(prince_rounds_Sbox_Input_s1[58]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[57]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[59]), .B(prince_rounds_Sbox_Input_s2[56]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(prince_rounds_Sbox_Input_s1[59]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[58]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[56]), .A2(prince_rounds_Sbox_Input_s2[59]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[56]), .A2(prince_rounds_Sbox_Input_s2[59]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(prince_rounds_Sbox_Input_s1[57]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F6_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n89), .A2(
        prince_rounds_Sbox_Input_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U31 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U28 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U21 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(prince_rounds_Sbox_Input_s2[59]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n89), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(prince_rounds_Sbox_Input_s1[58]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n89) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(prince_rounds_Sbox_Input_s1[58]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n69), .A2(
        prince_rounds_Sbox_Input_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U9 ( .A(
        prince_rounds_Sbox_Input_s1[58]), .B(prince_rounds_Sbox_Input_s2[59]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n78) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83), .B(
        prince_rounds_Sbox_Input_s1[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U3 ( .A1(
        prince_rounds_Sbox_Input_s1[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U2 ( .A(
        prince_rounds_Sbox_Input_s2[59]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n88), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(prince_rounds_Sbox_Input_s2[56]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F7_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[56]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[56]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n91) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U19 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U18 ( .A(
        prince_rounds_Sbox_Input_s2[58]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n85) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U14 ( .A(
        prince_rounds_Sbox_Input_s1[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n72) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[58]), .B(prince_rounds_Sbox_Input_s1[59]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n73) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[59]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[58]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[57]), .A2(prince_rounds_Sbox_Input_s2[58]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_0_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_1_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_2_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_3_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_4_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_5_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_6_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_7_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_8_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_9_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[56]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_n5), .ZN(
        output_s2[56]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[57]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_n5), .ZN(
        output_s2[57]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[58]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_n5), .ZN(
        output_s2[58]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[59]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_n5), .ZN(
        output_s2[59]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Inst_L_XORInst8_n6) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n79) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U30 ( .A(
        prince_rounds_Sbox_Input_s1[60]), .B(prince_rounds_Sbox_Input_s2[63]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U28 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n74), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n73), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n72), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U23 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n66), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[1]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n64) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n74), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n77), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n65) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U17 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n60), .B(
        prince_rounds_Sbox_Input_s1[60]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n70), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n61) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U15 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n59), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n66), .B(
        prince_rounds_Sbox_Input_s2[63]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n58), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n57) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U9 ( .A(
        prince_rounds_Sbox_Input_s2[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n58) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n56), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n75) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U5 ( .A(
        prince_rounds_Sbox_Input_s1[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n63), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n72), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n72) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U2 ( .A(
        prince_rounds_Sbox_Input_s1[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n77) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_U1 ( .A(
        prince_rounds_Sbox_Input_s1[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F1_n63) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U35 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n82) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U34 ( .A1(
        prince_rounds_Sbox_Input_s1[60]), .A2(prince_rounds_Sbox_Input_s2[62]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n76), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U30 ( .A1(
        prince_rounds_Sbox_Input_s1[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n76) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n73), .A2(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U27 ( .A1(
        prince_rounds_Sbox_Input_s1[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(prince_rounds_Sbox_Input_s1[60]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U23 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n68), .B(
        prince_rounds_Sbox_Input_s1[60]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n75), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n65), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[2]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n64), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n65) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n70) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U18 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(prince_rounds_Sbox_Input_s1[60]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n63), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n62), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n61), .A2(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n62) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n63) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n59) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n57), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n56) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n75), .A2(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n79) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U8 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n74), .A2(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U6 ( .A(
        prince_rounds_Sbox_Input_s1[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n60), .A2(
        prince_rounds_Sbox_Input_s1[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n57) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n60) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U3 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n67) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U2 ( .A(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n58) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_U1 ( .A(
        prince_rounds_Sbox_Input_s1[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F2_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U32 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n102), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n101), .S(
        prince_rounds_Sbox_Input_s2[61]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U31 ( .A(
        prince_rounds_Sbox_Input_s1[62]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n101) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n99), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n98), .S(
        prince_rounds_Sbox_Input_s1[63]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n97), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n99) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U25 ( .A1(
        prince_rounds_Sbox_Input_s1[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n93) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U24 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n102) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U23 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n92), .B(
        prince_rounds_Sbox_Input_s1[62]), .S(prince_rounds_Sbox_Input_s2[61]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n94) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U22 ( .A1(
        prince_rounds_Sbox_Input_s1[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n91), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n89) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U19 ( .A(
        prince_rounds_Sbox_Input_s2[61]), .B(prince_rounds_Sbox_Input_s1[62]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U17 ( .A1(
        prince_rounds_Sbox_Input_s1[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n85) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U16 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(prince_rounds_Sbox_Input_s1[60]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n84) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n86) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U14 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n91), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n91) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U12 ( .A(
        prince_rounds_Sbox_Input_s1[60]), .B(prince_rounds_Sbox_Input_s1[63]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n82), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U11 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(prince_rounds_Sbox_Input_s1[62]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n82) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[3]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U9 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U8 ( .A(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n83) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U6 ( .A1(
        prince_rounds_Sbox_Input_s1[62]), .A2(prince_rounds_Sbox_Input_s1[60]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[62]), .A2(prince_rounds_Sbox_Input_s1[60]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n96) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[3]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U3 ( .A(
        prince_rounds_Sbox_Input_s1[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U2 ( .A(
        prince_rounds_Sbox_Input_s1[63]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_U1 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(prince_rounds_Sbox_Input_s1[62]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F3_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U37 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U36 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n75) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U29 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n77), .B(
        prince_rounds_Sbox_Input_s2[61]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n76), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n72) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n73), .A2(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U27 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n66), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n66) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n64), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n63), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n63) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U19 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n73), .B(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n64) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n62), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n65), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n62) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U16 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n60), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n65) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n59), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n58), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n59) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n61), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n58) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U12 ( .A1(
        prince_rounds_Sbox_Input_s1[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n61) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n69) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U10 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n73) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U9 ( .A(
        prince_rounds_Sbox_Input_s2[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n60), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n56), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[4]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n56) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U5 ( .A(
        prince_rounds_Sbox_Input_s1[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U4 ( .A1(
        prince_rounds_Sbox_Input_s1[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U3 ( .A(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U2 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n57), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n60) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_U1 ( .A(
        prince_rounds_Sbox_Input_s2[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F4_n57) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U36 ( .A(
        prince_rounds_Sbox_Input_s1[63]), .B(prince_rounds_Sbox_Input_s2[60]), 
        .S(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n101), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n101) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n98), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U33 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n97), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n98) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n97) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[5]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U30 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s2[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n94) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n95), .A2(
        prince_rounds_Sbox_Input_s1[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n90) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n92), .B(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U26 ( .A1(
        prince_rounds_Sbox_Input_s2[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n99), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n84) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U21 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n82), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n93), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n92), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U20 ( .A1(
        prince_rounds_Sbox_Input_s1[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[5]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n83), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n80) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n78) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U15 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n95), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n76) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n75) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n74) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U9 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n96), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U7 ( .A(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n96) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U6 ( .A(
        prince_rounds_Sbox_Input_s1[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n100) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n92) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U4 ( .A(
        prince_rounds_Sbox_Input_s1[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n81) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U2 ( .A(
        prince_rounds_Sbox_Input_s2[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n95) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_U1 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(prince_rounds_Sbox_Input_s1[63]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F5_n86) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U39 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n107), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n106), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n104), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n106) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U37 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n103), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n102), .S(
        prince_rounds_Sbox_Input_s2[62]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n107) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U36 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n101), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n103) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n100), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n99), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n105), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n98), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n99) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U33 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n98) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[6]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U31 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n94), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n100), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n93), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n95) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n92), .A2(
        prince_rounds_Sbox_Input_s2[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U28 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n87), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n86), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U23 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n85) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n102), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n88) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U21 ( .A1(
        prince_rounds_Sbox_Input_s2[60]), .A2(prince_rounds_Sbox_Input_s2[63]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n102) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n101), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n83) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U18 ( .A1(
        prince_rounds_Sbox_Input_s2[60]), .A2(prince_rounds_Sbox_Input_s2[63]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n101) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n82), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n81), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n81) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n80), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n92), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n100), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U14 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n92), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n80) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U13 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n105), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(prince_rounds_Sbox_Input_s1[61]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n105) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U11 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n97), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U10 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n93), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n97) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U9 ( .A(
        prince_rounds_Sbox_Input_s1[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U8 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[6]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U7 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n104), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U6 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n100), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n89) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n104) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U4 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n100), .A2(
        prince_rounds_Sbox_Input_s2[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n94) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U3 ( .A(
        prince_rounds_Sbox_Input_s2[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n100) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U2 ( .A1(
        prince_rounds_Sbox_Input_s1[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n78) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_U1 ( .A(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F6_n79) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[7]) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n92) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U33 ( .A1(
        prince_rounds_Sbox_Input_s1[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n90) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U32 ( .A1(
        prince_rounds_Sbox_Input_s1[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n88) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U30 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U29 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n87) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U27 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n81), .A2(
        prince_rounds_Sbox_Input_s2[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n82) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n80), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n81) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U25 ( .A1(
        prince_rounds_Sbox_Input_s2[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n80) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U24 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n77), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n77) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U22 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(prince_rounds_Sbox_Input_s1[62]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n79), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n75), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[7]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U20 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n85), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n74), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n75) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84), .A2(
        prince_rounds_Sbox_Input_s1[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n74) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U17 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n72), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n71), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U16 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n71) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U15 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n73), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n72) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U14 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n85) );
  AND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U13 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84), .A2(
        prince_rounds_Sbox_Input_s1[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n73) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U12 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n70), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[7]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U11 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n69), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n70) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U10 ( .A(
        prince_rounds_Sbox_Input_s2[63]), .B(prince_rounds_Sbox_Input_s1[62]), 
        .Z(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n68), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n91), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U8 ( .A1(
        prince_rounds_Sbox_Input_s2[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n91) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U7 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89), .B(
        prince_rounds_Sbox_Input_s1[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n68) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U6 ( .A(
        prince_rounds_Sbox_Input_s2[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U5 ( .A1(
        prince_rounds_Sbox_Input_s1[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U4 ( .A(
        prince_rounds_Sbox_Input_s2[63]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n83), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n67) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84), .A2(
        prince_rounds_Sbox_Input_s2[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n84) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_U1 ( .A(
        prince_rounds_Sbox_Input_s2[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F7_n78) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U38 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n96), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n95), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U37 ( .A1(
        prince_rounds_Sbox_Input_s1[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n94), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n95) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U36 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n93), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n96) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U35 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n91), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n90), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n93) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U34 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n89), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U33 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n87), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n86), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n89) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U32 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n84), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n86) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U31 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n84) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U30 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n87) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U29 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n81), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n80), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U28 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n83), .A2(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n80) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U27 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88), .B(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n81) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U26 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n90), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n79), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U25 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n94), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n92), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n79) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U24 ( .A1(
        prince_rounds_Sbox_Input_s2[60]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n78), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n92) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U23 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n94) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U22 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n77), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n76), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U21 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n85), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n76) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U20 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n74), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n77) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U19 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n73), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U18 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n74), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n73) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U17 ( .A(
        prince_rounds_Sbox_Input_s2[62]), .B(prince_rounds_Sbox_Input_s1[63]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n74) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U16 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n78), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n72), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[8]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U15 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n90), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n91), .S(
        prince_rounds_Sbox_Input_s2[60]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n72) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U14 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n85), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n91) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U13 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n85) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U12 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n82), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n90) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U11 ( .A(
        prince_rounds_Sbox_Input_s1[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n82) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U10 ( .A(
        prince_rounds_Sbox_Input_s2[62]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n78) );
  OR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U9 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n71), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n70), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[8]) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U8 ( .A1(
        prince_rounds_Sbox_Input_s1[63]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n69), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n70) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U7 ( .A1(
        prince_rounds_Sbox_Input_s2[62]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n68), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n69) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U6 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88), .A2(
        prince_rounds_Sbox_Input_s2[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n68) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U5 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n75), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n67), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n71) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U4 ( .A1(
        prince_rounds_Sbox_Input_s2[61]), .A2(prince_rounds_Sbox_Input_s2[62]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n67) );
  NOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U3 ( .A1(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n83), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n75) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U2 ( .A(
        prince_rounds_Sbox_Input_s2[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n83) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_U1 ( .A(
        prince_rounds_Sbox_Input_s2[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_N_F8_n88) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_U3 ( .A(
        roundHalf_Select_Signal), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n6) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n6), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_0_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_0_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_0_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_0_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_1_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_1_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_1_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_1_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_2_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_2_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_2_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_2_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_3_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_3_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_3_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_3_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_4_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_4_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_4_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_4_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_5_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_5_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_5_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_5_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_6_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_6_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_6_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_6_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_7_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_e_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_7_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_7_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_7_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_8_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_8_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_8_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_8_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_9_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_9_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_9_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_9_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_10_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_10_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_10_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_10_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_11_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_11_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_11_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_11_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_12_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_12_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_12_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_12_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_13_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_13_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_13_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_13_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_14_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_14_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_14_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_14_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_15_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_f_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_15_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_15_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_15_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_16_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[1]), .S(
        roundHalf_Select_Signal), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_16_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_16_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_16_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_17_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[2]), .S(
        roundHalf_Select_Signal), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_17_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_17_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_17_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_18_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_18_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_18_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_18_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_19_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[4]), .S(
        roundHalf_Select_Signal), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_19_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_19_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_19_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_20_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[5]), .S(
        roundHalf_Select_Signal), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_20_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_20_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_20_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_21_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_21_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_21_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_21_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_22_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_22_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_22_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_22_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_23_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_g_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_23_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_23_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_23_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[8]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_24_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[1]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_24_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_24_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_24_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[1]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_25_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[2]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_25_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_25_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_25_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[2]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_26_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[3]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_26_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_26_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_26_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[3]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_27_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[4]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[4]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_27_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_27_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_27_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[4]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_28_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[5]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_28_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_28_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_28_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[5]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_29_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[6]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_29_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_29_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_29_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[6]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_30_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[7]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n5), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_30_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_30_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_30_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[7]) , .QN());
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_31_SFFInst_U3 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_h_s[8]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_si[8]), .S(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_31_SFFInst_N3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_31_SFFInst_Q_reg ( 
        .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_ScanFF_GEN_SFF_31_SFFInst_N3), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[8]) , .QN());
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[60]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst1_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_n5), .ZN(
        output_s2[60]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_e_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst2_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[61]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst3_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_n5), .ZN(
        output_s2[61]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_f_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst4_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[62]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst5_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_n5), .ZN(
        output_s2[62]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_g_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst6_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_n5), .ZN(
        prince_rounds_sub_Inv_Result_s1[63]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst7_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_n5), .ZN(
        output_s2[63]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[6]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[7]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_h_reg[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Inst_L_XORInst8_n6) );
  XNOR2_X1 prince_rounds_mul_s1_U96 ( .A(prince_rounds_mul_input_s1[59]), .B(
        prince_rounds_mul_s1_n32), .ZN(prince_rounds_mul_result_s1[63]) );
  XNOR2_X1 prince_rounds_mul_s1_U95 ( .A(prince_rounds_mul_input_s1[63]), .B(
        prince_rounds_mul_s1_n32), .ZN(prince_rounds_mul_result_s1[51]) );
  XNOR2_X1 prince_rounds_mul_s1_U94 ( .A(prince_rounds_mul_input_s1[51]), .B(
        prince_rounds_mul_input_s1[55]), .ZN(prince_rounds_mul_s1_n32) );
  XNOR2_X1 prince_rounds_mul_s1_U93 ( .A(prince_rounds_mul_input_s1[62]), .B(
        prince_rounds_mul_s1_n31), .ZN(prince_rounds_mul_result_s1[62]) );
  XNOR2_X1 prince_rounds_mul_s1_U92 ( .A(prince_rounds_mul_input_s1[58]), .B(
        prince_rounds_mul_s1_n31), .ZN(prince_rounds_mul_result_s1[58]) );
  XNOR2_X1 prince_rounds_mul_s1_U91 ( .A(prince_rounds_mul_input_s1[50]), .B(
        prince_rounds_mul_input_s1[54]), .ZN(prince_rounds_mul_s1_n31) );
  XNOR2_X1 prince_rounds_mul_s1_U90 ( .A(prince_rounds_mul_input_s1[60]), .B(
        prince_rounds_mul_s1_n30), .ZN(prince_rounds_mul_result_s1[60]) );
  XNOR2_X1 prince_rounds_mul_s1_U89 ( .A(prince_rounds_mul_input_s1[48]), .B(
        prince_rounds_mul_s1_n30), .ZN(prince_rounds_mul_result_s1[48]) );
  XNOR2_X1 prince_rounds_mul_s1_U88 ( .A(prince_rounds_mul_input_s1[52]), .B(
        prince_rounds_mul_input_s1[56]), .ZN(prince_rounds_mul_s1_n30) );
  XNOR2_X1 prince_rounds_mul_s1_U87 ( .A(prince_rounds_mul_input_s1[42]), .B(
        prince_rounds_mul_s1_n29), .ZN(prince_rounds_mul_result_s1[46]) );
  XNOR2_X1 prince_rounds_mul_s1_U86 ( .A(prince_rounds_mul_input_s1[46]), .B(
        prince_rounds_mul_s1_n29), .ZN(prince_rounds_mul_result_s1[34]) );
  XNOR2_X1 prince_rounds_mul_s1_U85 ( .A(prince_rounds_mul_input_s1[34]), .B(
        prince_rounds_mul_input_s1[38]), .ZN(prince_rounds_mul_s1_n29) );
  XNOR2_X1 prince_rounds_mul_s1_U84 ( .A(prince_rounds_mul_input_s1[28]), .B(
        prince_rounds_mul_s1_n28), .ZN(prince_rounds_mul_result_s1[28]) );
  XNOR2_X1 prince_rounds_mul_s1_U83 ( .A(prince_rounds_mul_input_s1[20]), .B(
        prince_rounds_mul_s1_n28), .ZN(prince_rounds_mul_result_s1[20]) );
  XNOR2_X1 prince_rounds_mul_s1_U82 ( .A(prince_rounds_mul_input_s1[24]), .B(
        prince_rounds_mul_input_s1[16]), .ZN(prince_rounds_mul_s1_n28) );
  XNOR2_X1 prince_rounds_mul_s1_U81 ( .A(prince_rounds_mul_input_s1[31]), .B(
        prince_rounds_mul_s1_n27), .ZN(prince_rounds_mul_result_s1[27]) );
  XNOR2_X1 prince_rounds_mul_s1_U80 ( .A(prince_rounds_mul_input_s1[23]), .B(
        prince_rounds_mul_s1_n27), .ZN(prince_rounds_mul_result_s1[19]) );
  XNOR2_X1 prince_rounds_mul_s1_U79 ( .A(prince_rounds_mul_input_s1[19]), .B(
        prince_rounds_mul_input_s1[27]), .ZN(prince_rounds_mul_s1_n27) );
  XNOR2_X1 prince_rounds_mul_s1_U78 ( .A(prince_rounds_mul_input_s1[45]), .B(
        prince_rounds_mul_s1_n26), .ZN(prince_rounds_mul_result_s1[45]) );
  XNOR2_X1 prince_rounds_mul_s1_U77 ( .A(prince_rounds_mul_input_s1[41]), .B(
        prince_rounds_mul_s1_n26), .ZN(prince_rounds_mul_result_s1[41]) );
  XNOR2_X1 prince_rounds_mul_s1_U76 ( .A(prince_rounds_mul_input_s1[33]), .B(
        prince_rounds_mul_input_s1[37]), .ZN(prince_rounds_mul_s1_n26) );
  XNOR2_X1 prince_rounds_mul_s1_U75 ( .A(prince_rounds_mul_input_s1[22]), .B(
        prince_rounds_mul_s1_n25), .ZN(prince_rounds_mul_result_s1[26]) );
  XNOR2_X1 prince_rounds_mul_s1_U74 ( .A(prince_rounds_mul_input_s1[18]), .B(
        prince_rounds_mul_s1_n25), .ZN(prince_rounds_mul_result_s1[22]) );
  XNOR2_X1 prince_rounds_mul_s1_U73 ( .A(prince_rounds_mul_input_s1[30]), .B(
        prince_rounds_mul_input_s1[26]), .ZN(prince_rounds_mul_s1_n25) );
  XNOR2_X1 prince_rounds_mul_s1_U72 ( .A(prince_rounds_mul_input_s1[16]), .B(
        prince_rounds_mul_s1_n24), .ZN(prince_rounds_mul_result_s1[24]) );
  XNOR2_X1 prince_rounds_mul_s1_U71 ( .A(prince_rounds_mul_input_s1[24]), .B(
        prince_rounds_mul_s1_n24), .ZN(prince_rounds_mul_result_s1[16]) );
  XNOR2_X1 prince_rounds_mul_s1_U70 ( .A(prince_rounds_mul_input_s1[28]), .B(
        prince_rounds_mul_input_s1[20]), .ZN(prince_rounds_mul_s1_n24) );
  XNOR2_X1 prince_rounds_mul_s1_U69 ( .A(prince_rounds_mul_input_s1[55]), .B(
        prince_rounds_mul_s1_n23), .ZN(prince_rounds_mul_result_s1[59]) );
  XNOR2_X1 prince_rounds_mul_s1_U68 ( .A(prince_rounds_mul_input_s1[51]), .B(
        prince_rounds_mul_s1_n23), .ZN(prince_rounds_mul_result_s1[55]) );
  XNOR2_X1 prince_rounds_mul_s1_U67 ( .A(prince_rounds_mul_input_s1[59]), .B(
        prince_rounds_mul_input_s1[63]), .ZN(prince_rounds_mul_s1_n23) );
  XNOR2_X1 prince_rounds_mul_s1_U66 ( .A(prince_rounds_mul_input_s1[21]), .B(
        prince_rounds_mul_s1_n22), .ZN(prince_rounds_mul_result_s1[21]) );
  XNOR2_X1 prince_rounds_mul_s1_U65 ( .A(prince_rounds_mul_input_s1[17]), .B(
        prince_rounds_mul_s1_n22), .ZN(prince_rounds_mul_result_s1[17]) );
  XNOR2_X1 prince_rounds_mul_s1_U64 ( .A(prince_rounds_mul_input_s1[25]), .B(
        prince_rounds_mul_input_s1[29]), .ZN(prince_rounds_mul_s1_n22) );
  XNOR2_X1 prince_rounds_mul_s1_U63 ( .A(prince_rounds_mul_input_s1[7]), .B(
        prince_rounds_mul_s1_n21), .ZN(prince_rounds_mul_result_s1[15]) );
  XNOR2_X1 prince_rounds_mul_s1_U62 ( .A(prince_rounds_mul_input_s1[15]), .B(
        prince_rounds_mul_s1_n21), .ZN(prince_rounds_mul_result_s1[7]) );
  XNOR2_X1 prince_rounds_mul_s1_U61 ( .A(prince_rounds_mul_input_s1[3]), .B(
        prince_rounds_mul_input_s1[11]), .ZN(prince_rounds_mul_s1_n21) );
  XNOR2_X1 prince_rounds_mul_s1_U60 ( .A(prince_rounds_mul_input_s1[44]), .B(
        prince_rounds_mul_s1_n20), .ZN(prince_rounds_mul_result_s1[44]) );
  XNOR2_X1 prince_rounds_mul_s1_U59 ( .A(prince_rounds_mul_input_s1[36]), .B(
        prince_rounds_mul_s1_n20), .ZN(prince_rounds_mul_result_s1[36]) );
  XNOR2_X1 prince_rounds_mul_s1_U58 ( .A(prince_rounds_mul_input_s1[40]), .B(
        prince_rounds_mul_input_s1[32]), .ZN(prince_rounds_mul_s1_n20) );
  XNOR2_X1 prince_rounds_mul_s1_U57 ( .A(prince_rounds_mul_input_s1[11]), .B(
        prince_rounds_mul_s1_n19), .ZN(prince_rounds_mul_result_s1[11]) );
  XNOR2_X1 prince_rounds_mul_s1_U56 ( .A(prince_rounds_mul_input_s1[3]), .B(
        prince_rounds_mul_s1_n19), .ZN(prince_rounds_mul_result_s1[3]) );
  XNOR2_X1 prince_rounds_mul_s1_U55 ( .A(prince_rounds_mul_input_s1[7]), .B(
        prince_rounds_mul_input_s1[15]), .ZN(prince_rounds_mul_s1_n19) );
  XNOR2_X1 prince_rounds_mul_s1_U54 ( .A(prince_rounds_mul_input_s1[6]), .B(
        prince_rounds_mul_s1_n18), .ZN(prince_rounds_mul_result_s1[14]) );
  XNOR2_X1 prince_rounds_mul_s1_U53 ( .A(prince_rounds_mul_input_s1[10]), .B(
        prince_rounds_mul_s1_n18), .ZN(prince_rounds_mul_result_s1[2]) );
  XNOR2_X1 prince_rounds_mul_s1_U52 ( .A(prince_rounds_mul_input_s1[14]), .B(
        prince_rounds_mul_input_s1[2]), .ZN(prince_rounds_mul_s1_n18) );
  XNOR2_X1 prince_rounds_mul_s1_U51 ( .A(prince_rounds_mul_input_s1[61]), .B(
        prince_rounds_mul_s1_n17), .ZN(prince_rounds_mul_result_s1[61]) );
  XNOR2_X1 prince_rounds_mul_s1_U50 ( .A(prince_rounds_mul_input_s1[53]), .B(
        prince_rounds_mul_s1_n17), .ZN(prince_rounds_mul_result_s1[53]) );
  XNOR2_X1 prince_rounds_mul_s1_U49 ( .A(prince_rounds_mul_input_s1[57]), .B(
        prince_rounds_mul_input_s1[49]), .ZN(prince_rounds_mul_s1_n17) );
  XNOR2_X1 prince_rounds_mul_s1_U48 ( .A(prince_rounds_mul_input_s1[49]), .B(
        prince_rounds_mul_s1_n16), .ZN(prince_rounds_mul_result_s1[57]) );
  XNOR2_X1 prince_rounds_mul_s1_U47 ( .A(prince_rounds_mul_input_s1[57]), .B(
        prince_rounds_mul_s1_n16), .ZN(prince_rounds_mul_result_s1[49]) );
  XNOR2_X1 prince_rounds_mul_s1_U46 ( .A(prince_rounds_mul_input_s1[61]), .B(
        prince_rounds_mul_input_s1[53]), .ZN(prince_rounds_mul_s1_n16) );
  XNOR2_X1 prince_rounds_mul_s1_U45 ( .A(prince_rounds_mul_input_s1[2]), .B(
        prince_rounds_mul_s1_n15), .ZN(prince_rounds_mul_result_s1[10]) );
  XNOR2_X1 prince_rounds_mul_s1_U44 ( .A(prince_rounds_mul_input_s1[14]), .B(
        prince_rounds_mul_s1_n15), .ZN(prince_rounds_mul_result_s1[6]) );
  XNOR2_X1 prince_rounds_mul_s1_U43 ( .A(prince_rounds_mul_input_s1[6]), .B(
        prince_rounds_mul_input_s1[10]), .ZN(prince_rounds_mul_s1_n15) );
  XNOR2_X1 prince_rounds_mul_s1_U42 ( .A(prince_rounds_mul_input_s1[9]), .B(
        prince_rounds_mul_s1_n14), .ZN(prince_rounds_mul_result_s1[13]) );
  XNOR2_X1 prince_rounds_mul_s1_U41 ( .A(prince_rounds_mul_input_s1[5]), .B(
        prince_rounds_mul_s1_n14), .ZN(prince_rounds_mul_result_s1[9]) );
  XNOR2_X1 prince_rounds_mul_s1_U40 ( .A(prince_rounds_mul_input_s1[13]), .B(
        prince_rounds_mul_input_s1[1]), .ZN(prince_rounds_mul_s1_n14) );
  XNOR2_X1 prince_rounds_mul_s1_U39 ( .A(prince_rounds_mul_input_s1[47]), .B(
        prince_rounds_mul_s1_n13), .ZN(prince_rounds_mul_result_s1[43]) );
  XNOR2_X1 prince_rounds_mul_s1_U38 ( .A(prince_rounds_mul_input_s1[39]), .B(
        prince_rounds_mul_s1_n13), .ZN(prince_rounds_mul_result_s1[35]) );
  XNOR2_X1 prince_rounds_mul_s1_U37 ( .A(prince_rounds_mul_input_s1[35]), .B(
        prince_rounds_mul_input_s1[43]), .ZN(prince_rounds_mul_s1_n13) );
  XNOR2_X1 prince_rounds_mul_s1_U36 ( .A(prince_rounds_mul_input_s1[8]), .B(
        prince_rounds_mul_s1_n12), .ZN(prince_rounds_mul_result_s1[12]) );
  XNOR2_X1 prince_rounds_mul_s1_U35 ( .A(prince_rounds_mul_input_s1[0]), .B(
        prince_rounds_mul_s1_n12), .ZN(prince_rounds_mul_result_s1[4]) );
  XNOR2_X1 prince_rounds_mul_s1_U34 ( .A(prince_rounds_mul_input_s1[4]), .B(
        prince_rounds_mul_input_s1[12]), .ZN(prince_rounds_mul_s1_n12) );
  XNOR2_X1 prince_rounds_mul_s1_U33 ( .A(prince_rounds_mul_input_s1[56]), .B(
        prince_rounds_mul_s1_n11), .ZN(prince_rounds_mul_result_s1[56]) );
  XNOR2_X1 prince_rounds_mul_s1_U32 ( .A(prince_rounds_mul_input_s1[52]), .B(
        prince_rounds_mul_s1_n11), .ZN(prince_rounds_mul_result_s1[52]) );
  XNOR2_X1 prince_rounds_mul_s1_U31 ( .A(prince_rounds_mul_input_s1[60]), .B(
        prince_rounds_mul_input_s1[48]), .ZN(prince_rounds_mul_s1_n11) );
  XNOR2_X1 prince_rounds_mul_s1_U30 ( .A(prince_rounds_mul_input_s1[38]), .B(
        prince_rounds_mul_s1_n10), .ZN(prince_rounds_mul_result_s1[42]) );
  XNOR2_X1 prince_rounds_mul_s1_U29 ( .A(prince_rounds_mul_input_s1[34]), .B(
        prince_rounds_mul_s1_n10), .ZN(prince_rounds_mul_result_s1[38]) );
  XNOR2_X1 prince_rounds_mul_s1_U28 ( .A(prince_rounds_mul_input_s1[42]), .B(
        prince_rounds_mul_input_s1[46]), .ZN(prince_rounds_mul_s1_n10) );
  XNOR2_X1 prince_rounds_mul_s1_U27 ( .A(prince_rounds_mul_input_s1[32]), .B(
        prince_rounds_mul_s1_n9), .ZN(prince_rounds_mul_result_s1[40]) );
  XNOR2_X1 prince_rounds_mul_s1_U26 ( .A(prince_rounds_mul_input_s1[40]), .B(
        prince_rounds_mul_s1_n9), .ZN(prince_rounds_mul_result_s1[32]) );
  XNOR2_X1 prince_rounds_mul_s1_U25 ( .A(prince_rounds_mul_input_s1[44]), .B(
        prince_rounds_mul_input_s1[36]), .ZN(prince_rounds_mul_s1_n9) );
  XNOR2_X1 prince_rounds_mul_s1_U24 ( .A(prince_rounds_mul_input_s1[1]), .B(
        prince_rounds_mul_s1_n8), .ZN(prince_rounds_mul_result_s1[5]) );
  XNOR2_X1 prince_rounds_mul_s1_U23 ( .A(prince_rounds_mul_input_s1[13]), .B(
        prince_rounds_mul_s1_n8), .ZN(prince_rounds_mul_result_s1[1]) );
  XNOR2_X1 prince_rounds_mul_s1_U22 ( .A(prince_rounds_mul_input_s1[9]), .B(
        prince_rounds_mul_input_s1[5]), .ZN(prince_rounds_mul_s1_n8) );
  XNOR2_X1 prince_rounds_mul_s1_U21 ( .A(prince_rounds_mul_input_s1[12]), .B(
        prince_rounds_mul_s1_n7), .ZN(prince_rounds_mul_result_s1[8]) );
  XNOR2_X1 prince_rounds_mul_s1_U20 ( .A(prince_rounds_mul_input_s1[4]), .B(
        prince_rounds_mul_s1_n7), .ZN(prince_rounds_mul_result_s1[0]) );
  XNOR2_X1 prince_rounds_mul_s1_U19 ( .A(prince_rounds_mul_input_s1[8]), .B(
        prince_rounds_mul_input_s1[0]), .ZN(prince_rounds_mul_s1_n7) );
  XNOR2_X1 prince_rounds_mul_s1_U18 ( .A(prince_rounds_mul_input_s1[54]), .B(
        prince_rounds_mul_s1_n6), .ZN(prince_rounds_mul_result_s1[54]) );
  XNOR2_X1 prince_rounds_mul_s1_U17 ( .A(prince_rounds_mul_input_s1[50]), .B(
        prince_rounds_mul_s1_n6), .ZN(prince_rounds_mul_result_s1[50]) );
  XNOR2_X1 prince_rounds_mul_s1_U16 ( .A(prince_rounds_mul_input_s1[62]), .B(
        prince_rounds_mul_input_s1[58]), .ZN(prince_rounds_mul_s1_n6) );
  XNOR2_X1 prince_rounds_mul_s1_U15 ( .A(prince_rounds_mul_input_s1[37]), .B(
        prince_rounds_mul_s1_n5), .ZN(prince_rounds_mul_result_s1[37]) );
  XNOR2_X1 prince_rounds_mul_s1_U14 ( .A(prince_rounds_mul_input_s1[33]), .B(
        prince_rounds_mul_s1_n5), .ZN(prince_rounds_mul_result_s1[33]) );
  XNOR2_X1 prince_rounds_mul_s1_U13 ( .A(prince_rounds_mul_input_s1[45]), .B(
        prince_rounds_mul_input_s1[41]), .ZN(prince_rounds_mul_s1_n5) );
  XNOR2_X1 prince_rounds_mul_s1_U12 ( .A(prince_rounds_mul_input_s1[27]), .B(
        prince_rounds_mul_s1_n4), .ZN(prince_rounds_mul_result_s1[31]) );
  XNOR2_X1 prince_rounds_mul_s1_U11 ( .A(prince_rounds_mul_input_s1[19]), .B(
        prince_rounds_mul_s1_n4), .ZN(prince_rounds_mul_result_s1[23]) );
  XNOR2_X1 prince_rounds_mul_s1_U10 ( .A(prince_rounds_mul_input_s1[31]), .B(
        prince_rounds_mul_input_s1[23]), .ZN(prince_rounds_mul_s1_n4) );
  XNOR2_X1 prince_rounds_mul_s1_U9 ( .A(prince_rounds_mul_input_s1[43]), .B(
        prince_rounds_mul_s1_n3), .ZN(prince_rounds_mul_result_s1[47]) );
  XNOR2_X1 prince_rounds_mul_s1_U8 ( .A(prince_rounds_mul_input_s1[35]), .B(
        prince_rounds_mul_s1_n3), .ZN(prince_rounds_mul_result_s1[39]) );
  XNOR2_X1 prince_rounds_mul_s1_U7 ( .A(prince_rounds_mul_input_s1[47]), .B(
        prince_rounds_mul_input_s1[39]), .ZN(prince_rounds_mul_s1_n3) );
  XNOR2_X1 prince_rounds_mul_s1_U6 ( .A(prince_rounds_mul_input_s1[26]), .B(
        prince_rounds_mul_s1_n2), .ZN(prince_rounds_mul_result_s1[30]) );
  XNOR2_X1 prince_rounds_mul_s1_U5 ( .A(prince_rounds_mul_input_s1[30]), .B(
        prince_rounds_mul_s1_n2), .ZN(prince_rounds_mul_result_s1[18]) );
  XNOR2_X1 prince_rounds_mul_s1_U4 ( .A(prince_rounds_mul_input_s1[22]), .B(
        prince_rounds_mul_input_s1[18]), .ZN(prince_rounds_mul_s1_n2) );
  XNOR2_X1 prince_rounds_mul_s1_U3 ( .A(prince_rounds_mul_input_s1[29]), .B(
        prince_rounds_mul_s1_n1), .ZN(prince_rounds_mul_result_s1[29]) );
  XNOR2_X1 prince_rounds_mul_s1_U2 ( .A(prince_rounds_mul_input_s1[25]), .B(
        prince_rounds_mul_s1_n1), .ZN(prince_rounds_mul_result_s1[25]) );
  XNOR2_X1 prince_rounds_mul_s1_U1 ( .A(prince_rounds_mul_input_s1[21]), .B(
        prince_rounds_mul_input_s1[17]), .ZN(prince_rounds_mul_s1_n1) );
  XNOR2_X1 prince_rounds_mul_s2_U96 ( .A(prince_rounds_mul_input_s2[59]), .B(
        prince_rounds_mul_s2_n96), .ZN(prince_rounds_mul_result_s2[63]) );
  XNOR2_X1 prince_rounds_mul_s2_U95 ( .A(prince_rounds_mul_input_s2[63]), .B(
        prince_rounds_mul_s2_n96), .ZN(prince_rounds_mul_result_s2[51]) );
  XNOR2_X1 prince_rounds_mul_s2_U94 ( .A(prince_rounds_mul_input_s2[51]), .B(
        prince_rounds_mul_input_s2[55]), .ZN(prince_rounds_mul_s2_n96) );
  XNOR2_X1 prince_rounds_mul_s2_U93 ( .A(prince_rounds_mul_input_s2[62]), .B(
        prince_rounds_mul_s2_n95), .ZN(prince_rounds_mul_result_s2[62]) );
  XNOR2_X1 prince_rounds_mul_s2_U92 ( .A(prince_rounds_mul_input_s2[58]), .B(
        prince_rounds_mul_s2_n95), .ZN(prince_rounds_mul_result_s2[58]) );
  XNOR2_X1 prince_rounds_mul_s2_U91 ( .A(prince_rounds_mul_input_s2[50]), .B(
        prince_rounds_mul_input_s2[54]), .ZN(prince_rounds_mul_s2_n95) );
  XNOR2_X1 prince_rounds_mul_s2_U90 ( .A(prince_rounds_mul_input_s2[60]), .B(
        prince_rounds_mul_s2_n94), .ZN(prince_rounds_mul_result_s2[60]) );
  XNOR2_X1 prince_rounds_mul_s2_U89 ( .A(prince_rounds_mul_input_s2[48]), .B(
        prince_rounds_mul_s2_n94), .ZN(prince_rounds_mul_result_s2[48]) );
  XNOR2_X1 prince_rounds_mul_s2_U88 ( .A(prince_rounds_mul_input_s2[52]), .B(
        prince_rounds_mul_input_s2[56]), .ZN(prince_rounds_mul_s2_n94) );
  XNOR2_X1 prince_rounds_mul_s2_U87 ( .A(prince_rounds_mul_input_s2[42]), .B(
        prince_rounds_mul_s2_n93), .ZN(prince_rounds_mul_result_s2[46]) );
  XNOR2_X1 prince_rounds_mul_s2_U86 ( .A(prince_rounds_mul_input_s2[46]), .B(
        prince_rounds_mul_s2_n93), .ZN(prince_rounds_mul_result_s2[34]) );
  XNOR2_X1 prince_rounds_mul_s2_U85 ( .A(prince_rounds_mul_input_s2[34]), .B(
        prince_rounds_mul_input_s2[38]), .ZN(prince_rounds_mul_s2_n93) );
  XNOR2_X1 prince_rounds_mul_s2_U84 ( .A(prince_rounds_mul_input_s2[28]), .B(
        prince_rounds_mul_s2_n92), .ZN(prince_rounds_mul_result_s2[28]) );
  XNOR2_X1 prince_rounds_mul_s2_U83 ( .A(prince_rounds_mul_input_s2[20]), .B(
        prince_rounds_mul_s2_n92), .ZN(prince_rounds_mul_result_s2[20]) );
  XNOR2_X1 prince_rounds_mul_s2_U82 ( .A(prince_rounds_mul_input_s2[24]), .B(
        prince_rounds_mul_input_s2[16]), .ZN(prince_rounds_mul_s2_n92) );
  XNOR2_X1 prince_rounds_mul_s2_U81 ( .A(prince_rounds_mul_input_s2[31]), .B(
        prince_rounds_mul_s2_n91), .ZN(prince_rounds_mul_result_s2[27]) );
  XNOR2_X1 prince_rounds_mul_s2_U80 ( .A(prince_rounds_mul_input_s2[23]), .B(
        prince_rounds_mul_s2_n91), .ZN(prince_rounds_mul_result_s2[19]) );
  XNOR2_X1 prince_rounds_mul_s2_U79 ( .A(prince_rounds_mul_input_s2[19]), .B(
        prince_rounds_mul_input_s2[27]), .ZN(prince_rounds_mul_s2_n91) );
  XNOR2_X1 prince_rounds_mul_s2_U78 ( .A(prince_rounds_mul_input_s2[45]), .B(
        prince_rounds_mul_s2_n90), .ZN(prince_rounds_mul_result_s2[45]) );
  XNOR2_X1 prince_rounds_mul_s2_U77 ( .A(prince_rounds_mul_input_s2[41]), .B(
        prince_rounds_mul_s2_n90), .ZN(prince_rounds_mul_result_s2[41]) );
  XNOR2_X1 prince_rounds_mul_s2_U76 ( .A(prince_rounds_mul_input_s2[33]), .B(
        prince_rounds_mul_input_s2[37]), .ZN(prince_rounds_mul_s2_n90) );
  XNOR2_X1 prince_rounds_mul_s2_U75 ( .A(prince_rounds_mul_input_s2[22]), .B(
        prince_rounds_mul_s2_n89), .ZN(prince_rounds_mul_result_s2[26]) );
  XNOR2_X1 prince_rounds_mul_s2_U74 ( .A(prince_rounds_mul_input_s2[18]), .B(
        prince_rounds_mul_s2_n89), .ZN(prince_rounds_mul_result_s2[22]) );
  XNOR2_X1 prince_rounds_mul_s2_U73 ( .A(prince_rounds_mul_input_s2[30]), .B(
        prince_rounds_mul_input_s2[26]), .ZN(prince_rounds_mul_s2_n89) );
  XNOR2_X1 prince_rounds_mul_s2_U72 ( .A(prince_rounds_mul_input_s2[16]), .B(
        prince_rounds_mul_s2_n88), .ZN(prince_rounds_mul_result_s2[24]) );
  XNOR2_X1 prince_rounds_mul_s2_U71 ( .A(prince_rounds_mul_input_s2[24]), .B(
        prince_rounds_mul_s2_n88), .ZN(prince_rounds_mul_result_s2[16]) );
  XNOR2_X1 prince_rounds_mul_s2_U70 ( .A(prince_rounds_mul_input_s2[28]), .B(
        prince_rounds_mul_input_s2[20]), .ZN(prince_rounds_mul_s2_n88) );
  XNOR2_X1 prince_rounds_mul_s2_U69 ( .A(prince_rounds_mul_input_s2[55]), .B(
        prince_rounds_mul_s2_n87), .ZN(prince_rounds_mul_result_s2[59]) );
  XNOR2_X1 prince_rounds_mul_s2_U68 ( .A(prince_rounds_mul_input_s2[51]), .B(
        prince_rounds_mul_s2_n87), .ZN(prince_rounds_mul_result_s2[55]) );
  XNOR2_X1 prince_rounds_mul_s2_U67 ( .A(prince_rounds_mul_input_s2[59]), .B(
        prince_rounds_mul_input_s2[63]), .ZN(prince_rounds_mul_s2_n87) );
  XNOR2_X1 prince_rounds_mul_s2_U66 ( .A(prince_rounds_mul_input_s2[21]), .B(
        prince_rounds_mul_s2_n86), .ZN(prince_rounds_mul_result_s2[21]) );
  XNOR2_X1 prince_rounds_mul_s2_U65 ( .A(prince_rounds_mul_input_s2[17]), .B(
        prince_rounds_mul_s2_n86), .ZN(prince_rounds_mul_result_s2[17]) );
  XNOR2_X1 prince_rounds_mul_s2_U64 ( .A(prince_rounds_mul_input_s2[25]), .B(
        prince_rounds_mul_input_s2[29]), .ZN(prince_rounds_mul_s2_n86) );
  XNOR2_X1 prince_rounds_mul_s2_U63 ( .A(prince_rounds_mul_input_s2[7]), .B(
        prince_rounds_mul_s2_n85), .ZN(prince_rounds_mul_result_s2[15]) );
  XNOR2_X1 prince_rounds_mul_s2_U62 ( .A(prince_rounds_mul_input_s2[15]), .B(
        prince_rounds_mul_s2_n85), .ZN(prince_rounds_mul_result_s2[7]) );
  XNOR2_X1 prince_rounds_mul_s2_U61 ( .A(prince_rounds_mul_input_s2[3]), .B(
        prince_rounds_mul_input_s2[11]), .ZN(prince_rounds_mul_s2_n85) );
  XNOR2_X1 prince_rounds_mul_s2_U60 ( .A(prince_rounds_mul_input_s2[44]), .B(
        prince_rounds_mul_s2_n84), .ZN(prince_rounds_mul_result_s2[44]) );
  XNOR2_X1 prince_rounds_mul_s2_U59 ( .A(prince_rounds_mul_input_s2[36]), .B(
        prince_rounds_mul_s2_n84), .ZN(prince_rounds_mul_result_s2[36]) );
  XNOR2_X1 prince_rounds_mul_s2_U58 ( .A(prince_rounds_mul_input_s2[40]), .B(
        prince_rounds_mul_input_s2[32]), .ZN(prince_rounds_mul_s2_n84) );
  XNOR2_X1 prince_rounds_mul_s2_U57 ( .A(prince_rounds_mul_input_s2[11]), .B(
        prince_rounds_mul_s2_n83), .ZN(prince_rounds_mul_result_s2[11]) );
  XNOR2_X1 prince_rounds_mul_s2_U56 ( .A(prince_rounds_mul_input_s2[3]), .B(
        prince_rounds_mul_s2_n83), .ZN(prince_rounds_mul_result_s2[3]) );
  XNOR2_X1 prince_rounds_mul_s2_U55 ( .A(prince_rounds_mul_input_s2[7]), .B(
        prince_rounds_mul_input_s2[15]), .ZN(prince_rounds_mul_s2_n83) );
  XNOR2_X1 prince_rounds_mul_s2_U54 ( .A(prince_rounds_mul_input_s2[6]), .B(
        prince_rounds_mul_s2_n82), .ZN(prince_rounds_mul_result_s2[14]) );
  XNOR2_X1 prince_rounds_mul_s2_U53 ( .A(prince_rounds_mul_input_s2[10]), .B(
        prince_rounds_mul_s2_n82), .ZN(prince_rounds_mul_result_s2[2]) );
  XNOR2_X1 prince_rounds_mul_s2_U52 ( .A(prince_rounds_mul_input_s2[14]), .B(
        prince_rounds_mul_input_s2[2]), .ZN(prince_rounds_mul_s2_n82) );
  XNOR2_X1 prince_rounds_mul_s2_U51 ( .A(prince_rounds_mul_input_s2[61]), .B(
        prince_rounds_mul_s2_n81), .ZN(prince_rounds_mul_result_s2[61]) );
  XNOR2_X1 prince_rounds_mul_s2_U50 ( .A(prince_rounds_mul_input_s2[53]), .B(
        prince_rounds_mul_s2_n81), .ZN(prince_rounds_mul_result_s2[53]) );
  XNOR2_X1 prince_rounds_mul_s2_U49 ( .A(prince_rounds_mul_input_s2[57]), .B(
        prince_rounds_mul_input_s2[49]), .ZN(prince_rounds_mul_s2_n81) );
  XNOR2_X1 prince_rounds_mul_s2_U48 ( .A(prince_rounds_mul_input_s2[49]), .B(
        prince_rounds_mul_s2_n80), .ZN(prince_rounds_mul_result_s2[57]) );
  XNOR2_X1 prince_rounds_mul_s2_U47 ( .A(prince_rounds_mul_input_s2[57]), .B(
        prince_rounds_mul_s2_n80), .ZN(prince_rounds_mul_result_s2[49]) );
  XNOR2_X1 prince_rounds_mul_s2_U46 ( .A(prince_rounds_mul_input_s2[61]), .B(
        prince_rounds_mul_input_s2[53]), .ZN(prince_rounds_mul_s2_n80) );
  XNOR2_X1 prince_rounds_mul_s2_U45 ( .A(prince_rounds_mul_input_s2[2]), .B(
        prince_rounds_mul_s2_n79), .ZN(prince_rounds_mul_result_s2[10]) );
  XNOR2_X1 prince_rounds_mul_s2_U44 ( .A(prince_rounds_mul_input_s2[14]), .B(
        prince_rounds_mul_s2_n79), .ZN(prince_rounds_mul_result_s2[6]) );
  XNOR2_X1 prince_rounds_mul_s2_U43 ( .A(prince_rounds_mul_input_s2[6]), .B(
        prince_rounds_mul_input_s2[10]), .ZN(prince_rounds_mul_s2_n79) );
  XNOR2_X1 prince_rounds_mul_s2_U42 ( .A(prince_rounds_mul_input_s2[9]), .B(
        prince_rounds_mul_s2_n78), .ZN(prince_rounds_mul_result_s2[13]) );
  XNOR2_X1 prince_rounds_mul_s2_U41 ( .A(prince_rounds_mul_input_s2[5]), .B(
        prince_rounds_mul_s2_n78), .ZN(prince_rounds_mul_result_s2[9]) );
  XNOR2_X1 prince_rounds_mul_s2_U40 ( .A(prince_rounds_mul_input_s2[13]), .B(
        prince_rounds_mul_input_s2[1]), .ZN(prince_rounds_mul_s2_n78) );
  XNOR2_X1 prince_rounds_mul_s2_U39 ( .A(prince_rounds_mul_input_s2[47]), .B(
        prince_rounds_mul_s2_n77), .ZN(prince_rounds_mul_result_s2[43]) );
  XNOR2_X1 prince_rounds_mul_s2_U38 ( .A(prince_rounds_mul_input_s2[39]), .B(
        prince_rounds_mul_s2_n77), .ZN(prince_rounds_mul_result_s2[35]) );
  XNOR2_X1 prince_rounds_mul_s2_U37 ( .A(prince_rounds_mul_input_s2[35]), .B(
        prince_rounds_mul_input_s2[43]), .ZN(prince_rounds_mul_s2_n77) );
  XNOR2_X1 prince_rounds_mul_s2_U36 ( .A(prince_rounds_mul_input_s2[8]), .B(
        prince_rounds_mul_s2_n76), .ZN(prince_rounds_mul_result_s2[12]) );
  XNOR2_X1 prince_rounds_mul_s2_U35 ( .A(prince_rounds_mul_input_s2[0]), .B(
        prince_rounds_mul_s2_n76), .ZN(prince_rounds_mul_result_s2[4]) );
  XNOR2_X1 prince_rounds_mul_s2_U34 ( .A(prince_rounds_mul_input_s2[4]), .B(
        prince_rounds_mul_input_s2[12]), .ZN(prince_rounds_mul_s2_n76) );
  XNOR2_X1 prince_rounds_mul_s2_U33 ( .A(prince_rounds_mul_input_s2[56]), .B(
        prince_rounds_mul_s2_n75), .ZN(prince_rounds_mul_result_s2[56]) );
  XNOR2_X1 prince_rounds_mul_s2_U32 ( .A(prince_rounds_mul_input_s2[52]), .B(
        prince_rounds_mul_s2_n75), .ZN(prince_rounds_mul_result_s2[52]) );
  XNOR2_X1 prince_rounds_mul_s2_U31 ( .A(prince_rounds_mul_input_s2[60]), .B(
        prince_rounds_mul_input_s2[48]), .ZN(prince_rounds_mul_s2_n75) );
  XNOR2_X1 prince_rounds_mul_s2_U30 ( .A(prince_rounds_mul_input_s2[38]), .B(
        prince_rounds_mul_s2_n74), .ZN(prince_rounds_mul_result_s2[42]) );
  XNOR2_X1 prince_rounds_mul_s2_U29 ( .A(prince_rounds_mul_input_s2[34]), .B(
        prince_rounds_mul_s2_n74), .ZN(prince_rounds_mul_result_s2[38]) );
  XNOR2_X1 prince_rounds_mul_s2_U28 ( .A(prince_rounds_mul_input_s2[42]), .B(
        prince_rounds_mul_input_s2[46]), .ZN(prince_rounds_mul_s2_n74) );
  XNOR2_X1 prince_rounds_mul_s2_U27 ( .A(prince_rounds_mul_input_s2[32]), .B(
        prince_rounds_mul_s2_n73), .ZN(prince_rounds_mul_result_s2[40]) );
  XNOR2_X1 prince_rounds_mul_s2_U26 ( .A(prince_rounds_mul_input_s2[40]), .B(
        prince_rounds_mul_s2_n73), .ZN(prince_rounds_mul_result_s2[32]) );
  XNOR2_X1 prince_rounds_mul_s2_U25 ( .A(prince_rounds_mul_input_s2[44]), .B(
        prince_rounds_mul_input_s2[36]), .ZN(prince_rounds_mul_s2_n73) );
  XNOR2_X1 prince_rounds_mul_s2_U24 ( .A(prince_rounds_mul_input_s2[1]), .B(
        prince_rounds_mul_s2_n72), .ZN(prince_rounds_mul_result_s2[5]) );
  XNOR2_X1 prince_rounds_mul_s2_U23 ( .A(prince_rounds_mul_input_s2[13]), .B(
        prince_rounds_mul_s2_n72), .ZN(prince_rounds_mul_result_s2[1]) );
  XNOR2_X1 prince_rounds_mul_s2_U22 ( .A(prince_rounds_mul_input_s2[9]), .B(
        prince_rounds_mul_input_s2[5]), .ZN(prince_rounds_mul_s2_n72) );
  XNOR2_X1 prince_rounds_mul_s2_U21 ( .A(prince_rounds_mul_input_s2[12]), .B(
        prince_rounds_mul_s2_n71), .ZN(prince_rounds_mul_result_s2[8]) );
  XNOR2_X1 prince_rounds_mul_s2_U20 ( .A(prince_rounds_mul_input_s2[4]), .B(
        prince_rounds_mul_s2_n71), .ZN(prince_rounds_mul_result_s2[0]) );
  XNOR2_X1 prince_rounds_mul_s2_U19 ( .A(prince_rounds_mul_input_s2[8]), .B(
        prince_rounds_mul_input_s2[0]), .ZN(prince_rounds_mul_s2_n71) );
  XNOR2_X1 prince_rounds_mul_s2_U18 ( .A(prince_rounds_mul_input_s2[54]), .B(
        prince_rounds_mul_s2_n70), .ZN(prince_rounds_mul_result_s2[54]) );
  XNOR2_X1 prince_rounds_mul_s2_U17 ( .A(prince_rounds_mul_input_s2[50]), .B(
        prince_rounds_mul_s2_n70), .ZN(prince_rounds_mul_result_s2[50]) );
  XNOR2_X1 prince_rounds_mul_s2_U16 ( .A(prince_rounds_mul_input_s2[62]), .B(
        prince_rounds_mul_input_s2[58]), .ZN(prince_rounds_mul_s2_n70) );
  XNOR2_X1 prince_rounds_mul_s2_U15 ( .A(prince_rounds_mul_input_s2[37]), .B(
        prince_rounds_mul_s2_n69), .ZN(prince_rounds_mul_result_s2[37]) );
  XNOR2_X1 prince_rounds_mul_s2_U14 ( .A(prince_rounds_mul_input_s2[33]), .B(
        prince_rounds_mul_s2_n69), .ZN(prince_rounds_mul_result_s2[33]) );
  XNOR2_X1 prince_rounds_mul_s2_U13 ( .A(prince_rounds_mul_input_s2[45]), .B(
        prince_rounds_mul_input_s2[41]), .ZN(prince_rounds_mul_s2_n69) );
  XNOR2_X1 prince_rounds_mul_s2_U12 ( .A(prince_rounds_mul_input_s2[27]), .B(
        prince_rounds_mul_s2_n68), .ZN(prince_rounds_mul_result_s2[31]) );
  XNOR2_X1 prince_rounds_mul_s2_U11 ( .A(prince_rounds_mul_input_s2[19]), .B(
        prince_rounds_mul_s2_n68), .ZN(prince_rounds_mul_result_s2[23]) );
  XNOR2_X1 prince_rounds_mul_s2_U10 ( .A(prince_rounds_mul_input_s2[31]), .B(
        prince_rounds_mul_input_s2[23]), .ZN(prince_rounds_mul_s2_n68) );
  XNOR2_X1 prince_rounds_mul_s2_U9 ( .A(prince_rounds_mul_input_s2[43]), .B(
        prince_rounds_mul_s2_n67), .ZN(prince_rounds_mul_result_s2[47]) );
  XNOR2_X1 prince_rounds_mul_s2_U8 ( .A(prince_rounds_mul_input_s2[35]), .B(
        prince_rounds_mul_s2_n67), .ZN(prince_rounds_mul_result_s2[39]) );
  XNOR2_X1 prince_rounds_mul_s2_U7 ( .A(prince_rounds_mul_input_s2[47]), .B(
        prince_rounds_mul_input_s2[39]), .ZN(prince_rounds_mul_s2_n67) );
  XNOR2_X1 prince_rounds_mul_s2_U6 ( .A(prince_rounds_mul_input_s2[26]), .B(
        prince_rounds_mul_s2_n66), .ZN(prince_rounds_mul_result_s2[30]) );
  XNOR2_X1 prince_rounds_mul_s2_U5 ( .A(prince_rounds_mul_input_s2[30]), .B(
        prince_rounds_mul_s2_n66), .ZN(prince_rounds_mul_result_s2[18]) );
  XNOR2_X1 prince_rounds_mul_s2_U4 ( .A(prince_rounds_mul_input_s2[22]), .B(
        prince_rounds_mul_input_s2[18]), .ZN(prince_rounds_mul_s2_n66) );
  XNOR2_X1 prince_rounds_mul_s2_U3 ( .A(prince_rounds_mul_input_s2[29]), .B(
        prince_rounds_mul_s2_n65), .ZN(prince_rounds_mul_result_s2[29]) );
  XNOR2_X1 prince_rounds_mul_s2_U2 ( .A(prince_rounds_mul_input_s2[25]), .B(
        prince_rounds_mul_s2_n65), .ZN(prince_rounds_mul_result_s2[25]) );
  XNOR2_X1 prince_rounds_mul_s2_U1 ( .A(prince_rounds_mul_input_s2[21]), .B(
        prince_rounds_mul_input_s2[17]), .ZN(prince_rounds_mul_s2_n65) );
endmodule

