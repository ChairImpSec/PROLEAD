
module circuit ( clk, rst, Plaintext0, Plaintext1, Plaintext2, Key0, Key1, 
        Key2, r, Ciphertext0, Ciphertext1, Ciphertext2, done );
  input [63:0] Plaintext0;
  input [63:0] Plaintext1;
  input [63:0] Plaintext2;
  input [127:0] Key0;
  input [127:0] Key1;
  input [127:0] Key2;
  input [71:0] r;
  output [63:0] Ciphertext0;
  output [63:0] Ciphertext1;
  output [63:0] Ciphertext2;
  input clk, rst;
  output done;
  wire   RoundFunctionEN, AddKey, SelKey, LED_RoundFunction0_n562,
         LED_RoundFunction0_n561, LED_RoundFunction0_n560,
         LED_RoundFunction0_n559, LED_RoundFunction0_n558,
         LED_RoundFunction0_n557, LED_RoundFunction0_n556,
         LED_RoundFunction0_n555, LED_RoundFunction0_n554,
         LED_RoundFunction0_n553, LED_RoundFunction0_n552,
         LED_RoundFunction0_n551, LED_RoundFunction0_n550,
         LED_RoundFunction0_n549, LED_RoundFunction0_n548,
         LED_RoundFunction0_n547, LED_RoundFunction0_n546,
         LED_RoundFunction0_n545, LED_RoundFunction0_n544,
         LED_RoundFunction0_n543, LED_RoundFunction0_n542,
         LED_RoundFunction0_n541, LED_RoundFunction0_n540,
         LED_RoundFunction0_n539, LED_RoundFunction0_n538,
         LED_RoundFunction0_n537, LED_RoundFunction0_n536,
         LED_RoundFunction0_n535, LED_RoundFunction0_n534,
         LED_RoundFunction0_n533, LED_RoundFunction0_n532,
         LED_RoundFunction0_n531, LED_RoundFunction0_n530,
         LED_RoundFunction0_n529, LED_RoundFunction0_n528,
         LED_RoundFunction0_n527, LED_RoundFunction0_n526,
         LED_RoundFunction0_n525, LED_RoundFunction0_n524,
         LED_RoundFunction0_n523, LED_RoundFunction0_n522,
         LED_RoundFunction0_n521, LED_RoundFunction0_n520,
         LED_RoundFunction0_n519, LED_RoundFunction0_n518,
         LED_RoundFunction0_n517, LED_RoundFunction0_n516,
         LED_RoundFunction0_n515, LED_RoundFunction0_n514,
         LED_RoundFunction0_n513, LED_RoundFunction0_n512,
         LED_RoundFunction0_n511, LED_RoundFunction0_n510,
         LED_RoundFunction0_n509, LED_RoundFunction0_n508,
         LED_RoundFunction0_n507, LED_RoundFunction0_n506,
         LED_RoundFunction0_n505, LED_RoundFunction0_n504,
         LED_RoundFunction0_n503, LED_RoundFunction0_n502,
         LED_RoundFunction0_n501, LED_RoundFunction0_n500,
         LED_RoundFunction0_n499, LED_RoundFunction0_n498,
         LED_RoundFunction0_n497, LED_RoundFunction0_n496,
         LED_RoundFunction0_n495, LED_RoundFunction0_n494,
         LED_RoundFunction0_n493, LED_RoundFunction0_n492,
         LED_RoundFunction0_n491, LED_RoundFunction0_n490,
         LED_RoundFunction0_n489, LED_RoundFunction0_n488,
         LED_RoundFunction0_n487, LED_RoundFunction0_n486,
         LED_RoundFunction0_n485, LED_RoundFunction0_n484,
         LED_RoundFunction0_n483, LED_RoundFunction0_n482,
         LED_RoundFunction0_n481, LED_RoundFunction0_n480,
         LED_RoundFunction0_n479, LED_RoundFunction0_n478,
         LED_RoundFunction0_n477, LED_RoundFunction0_n476,
         LED_RoundFunction0_n475, LED_RoundFunction0_n474,
         LED_RoundFunction0_n473, LED_RoundFunction0_n472,
         LED_RoundFunction0_n471, LED_RoundFunction0_n470,
         LED_RoundFunction0_n469, LED_RoundFunction0_n468,
         LED_RoundFunction0_n467, LED_RoundFunction0_n466,
         LED_RoundFunction0_n465, LED_RoundFunction0_n464,
         LED_RoundFunction0_n463, LED_RoundFunction0_n462,
         LED_RoundFunction0_n461, LED_RoundFunction0_n460,
         LED_RoundFunction0_n459, LED_RoundFunction0_n458,
         LED_RoundFunction0_n457, LED_RoundFunction0_n456,
         LED_RoundFunction0_n455, LED_RoundFunction0_n454,
         LED_RoundFunction0_n453, LED_RoundFunction0_n452,
         LED_RoundFunction0_n451, LED_RoundFunction0_n450,
         LED_RoundFunction0_n449, LED_RoundFunction0_n448,
         LED_RoundFunction0_n447, LED_RoundFunction0_n446,
         LED_RoundFunction0_n445, LED_RoundFunction0_n444,
         LED_RoundFunction0_n443, LED_RoundFunction0_n442,
         LED_RoundFunction0_n441, LED_RoundFunction0_n440,
         LED_RoundFunction0_n439, LED_RoundFunction0_n438,
         LED_RoundFunction0_n437, LED_RoundFunction0_n436,
         LED_RoundFunction0_n435, LED_RoundFunction0_n434,
         LED_RoundFunction0_n433, LED_RoundFunction0_n432,
         LED_RoundFunction0_n431, LED_RoundFunction0_n430,
         LED_RoundFunction0_n429, LED_RoundFunction0_n428,
         LED_RoundFunction0_n427, LED_RoundFunction0_n426,
         LED_RoundFunction0_n425, LED_RoundFunction0_n424,
         LED_RoundFunction0_n423, LED_RoundFunction0_n422,
         LED_RoundFunction0_n421, LED_RoundFunction0_n420,
         LED_RoundFunction0_n419, LED_RoundFunction0_n418,
         LED_RoundFunction0_n417, LED_RoundFunction0_n416,
         LED_RoundFunction0_n415, LED_RoundFunction0_n414,
         LED_RoundFunction0_n413, LED_RoundFunction0_n412,
         LED_RoundFunction0_n411, LED_RoundFunction0_n410,
         LED_RoundFunction0_n409, LED_RoundFunction0_n408,
         LED_RoundFunction0_n407, LED_RoundFunction0_n406,
         LED_RoundFunction0_n405, LED_RoundFunction0_n404,
         LED_RoundFunction0_n403, LED_RoundFunction0_n402,
         LED_RoundFunction0_n401, LED_RoundFunction0_n400,
         LED_RoundFunction0_n399, LED_RoundFunction0_n398,
         LED_RoundFunction0_n397, LED_RoundFunction0_n396,
         LED_RoundFunction0_n395, LED_RoundFunction0_n394,
         LED_RoundFunction0_n393, LED_RoundFunction0_n392,
         LED_RoundFunction0_n391, LED_RoundFunction0_n390,
         LED_RoundFunction0_n389, LED_RoundFunction0_n388,
         LED_RoundFunction0_n387, LED_RoundFunction0_n386,
         LED_RoundFunction0_n385, LED_RoundFunction0_n384,
         LED_RoundFunction0_n383, LED_RoundFunction0_n382,
         LED_RoundFunction0_n381, LED_RoundFunction0_n380,
         LED_RoundFunction0_n379, LED_RoundFunction0_n378,
         LED_RoundFunction0_n377, LED_RoundFunction0_n376,
         LED_RoundFunction0_n375, LED_RoundFunction0_n374,
         LED_RoundFunction0_n373, LED_RoundFunction0_n372,
         LED_RoundFunction0_n371, LED_RoundFunction0_n370,
         LED_RoundFunction0_n369, LED_RoundFunction0_n368,
         LED_RoundFunction0_n367, LED_RoundFunction0_n366,
         LED_RoundFunction0_n365, LED_RoundFunction0_n364,
         LED_RoundFunction0_n363, LED_RoundFunction0_n362,
         LED_RoundFunction0_n361, LED_RoundFunction0_n360,
         LED_RoundFunction0_n359, LED_RoundFunction0_n358,
         LED_RoundFunction0_n357, LED_RoundFunction0_n356,
         LED_RoundFunction0_n355, LED_RoundFunction0_n354,
         LED_RoundFunction0_n353, LED_RoundFunction0_n352,
         LED_RoundFunction0_n351, LED_RoundFunction0_n350,
         LED_RoundFunction0_n349, LED_RoundFunction0_n348,
         LED_RoundFunction0_n347, LED_RoundFunction0_n346,
         LED_RoundFunction0_n345, LED_RoundFunction0_n344,
         LED_RoundFunction0_n343, LED_RoundFunction0_n342,
         LED_RoundFunction0_n341, LED_RoundFunction0_n340,
         LED_RoundFunction0_n339, LED_RoundFunction0_n338,
         LED_RoundFunction0_n337, LED_RoundFunction0_n336,
         LED_RoundFunction0_n335, LED_RoundFunction0_n334,
         LED_RoundFunction0_n333, LED_RoundFunction0_n332,
         LED_RoundFunction0_n331, LED_RoundFunction0_n330,
         LED_RoundFunction0_n329, LED_RoundFunction0_n328,
         LED_RoundFunction0_n327, LED_RoundFunction0_n326,
         LED_RoundFunction0_n325, LED_RoundFunction0_n324,
         LED_RoundFunction0_n323, LED_RoundFunction0_n322,
         LED_RoundFunction0_n321, LED_RoundFunction0_n320,
         LED_RoundFunction0_n319, LED_RoundFunction0_n318,
         LED_RoundFunction0_n317, LED_RoundFunction0_n316,
         LED_RoundFunction0_n315, LED_RoundFunction0_n314,
         LED_RoundFunction0_n313, LED_RoundFunction0_n312,
         LED_RoundFunction0_n311, LED_RoundFunction0_n310,
         LED_RoundFunction0_n309, LED_RoundFunction0_n308,
         LED_RoundFunction0_n307, LED_RoundFunction0_n306,
         LED_RoundFunction0_n305, LED_RoundFunction0_n304,
         LED_RoundFunction0_n303, LED_RoundFunction0_n302,
         LED_RoundFunction0_n301, LED_RoundFunction0_n300,
         LED_RoundFunction0_n299, LED_RoundFunction0_n298,
         LED_RoundFunction0_n297, LED_RoundFunction0_n296,
         LED_RoundFunction0_n295, LED_RoundFunction0_n294,
         LED_RoundFunction0_n293, LED_RoundFunction0_n292,
         LED_RoundFunction0_n291, LED_RoundFunction0_n290,
         LED_RoundFunction0_n289, LED_RoundFunction0_n288,
         LED_RoundFunction0_n287, LED_RoundFunction0_n286,
         LED_RoundFunction0_n285, LED_RoundFunction0_n284,
         LED_RoundFunction0_n283, LED_RoundFunction0_n282,
         LED_RoundFunction0_n281, LED_RoundFunction0_Feedback_0_,
         LED_RoundFunction0_Feedback_1_, LED_RoundFunction0_Feedback_2_,
         LED_RoundFunction0_Feedback_3_, LED_RoundFunction0_Feedback_4_,
         LED_RoundFunction0_Feedback_5_, LED_RoundFunction0_Feedback_6_,
         LED_RoundFunction0_Feedback_7_, LED_RoundFunction0_Feedback_8_,
         LED_RoundFunction0_Feedback_9_, LED_RoundFunction0_Feedback_10_,
         LED_RoundFunction0_Feedback_11_, LED_RoundFunction0_Feedback_12_,
         LED_RoundFunction0_Feedback_13_, LED_RoundFunction0_Feedback_14_,
         LED_RoundFunction0_Feedback_15_, LED_RoundFunction0_Feedback_16_,
         LED_RoundFunction0_Feedback_17_, LED_RoundFunction0_Feedback_18_,
         LED_RoundFunction0_Feedback_19_, LED_RoundFunction0_Feedback_20_,
         LED_RoundFunction0_Feedback_21_, LED_RoundFunction0_Feedback_22_,
         LED_RoundFunction0_Feedback_23_, LED_RoundFunction0_Feedback_24_,
         LED_RoundFunction0_Feedback_25_, LED_RoundFunction0_Feedback_26_,
         LED_RoundFunction0_Feedback_27_, LED_RoundFunction0_Feedback_28_,
         LED_RoundFunction0_Feedback_29_, LED_RoundFunction0_Feedback_30_,
         LED_RoundFunction0_Feedback_31_, LED_RoundFunction0_Feedback_32_,
         LED_RoundFunction0_Feedback_33_, LED_RoundFunction0_Feedback_34_,
         LED_RoundFunction0_Feedback_35_, LED_RoundFunction0_Feedback_36_,
         LED_RoundFunction0_Feedback_37_, LED_RoundFunction0_Feedback_38_,
         LED_RoundFunction0_Feedback_39_, LED_RoundFunction0_Feedback_40_,
         LED_RoundFunction0_Feedback_41_, LED_RoundFunction0_Feedback_42_,
         LED_RoundFunction0_Feedback_43_, LED_RoundFunction0_Feedback_44_,
         LED_RoundFunction0_Feedback_45_, LED_RoundFunction0_Feedback_46_,
         LED_RoundFunction0_Feedback_47_, LED_RoundFunction0_Feedback_48_,
         LED_RoundFunction0_Feedback_49_, LED_RoundFunction0_Feedback_50_,
         LED_RoundFunction0_Feedback_51_, LED_RoundFunction0_Feedback_52_,
         LED_RoundFunction0_Feedback_53_, LED_RoundFunction0_Feedback_54_,
         LED_RoundFunction0_Feedback_55_, LED_RoundFunction0_Feedback_56_,
         LED_RoundFunction0_Feedback_57_, LED_RoundFunction0_Feedback_58_,
         LED_RoundFunction0_Feedback_59_, LED_RoundFunction0_Feedback_60_,
         LED_RoundFunction0_Feedback_61_, LED_RoundFunction0_Feedback_62_,
         LED_RoundFunction0_Feedback_63_, LED_RoundFunction0_MCInst1_MC0_n160,
         LED_RoundFunction0_MCInst1_MC0_n159,
         LED_RoundFunction0_MCInst1_MC0_n158,
         LED_RoundFunction0_MCInst1_MC0_n157,
         LED_RoundFunction0_MCInst1_MC0_n156,
         LED_RoundFunction0_MCInst1_MC0_n155,
         LED_RoundFunction0_MCInst1_MC0_n154,
         LED_RoundFunction0_MCInst1_MC0_n153,
         LED_RoundFunction0_MCInst1_MC0_n152,
         LED_RoundFunction0_MCInst1_MC0_n151,
         LED_RoundFunction0_MCInst1_MC0_n150,
         LED_RoundFunction0_MCInst1_MC0_n149,
         LED_RoundFunction0_MCInst1_MC0_n148,
         LED_RoundFunction0_MCInst1_MC0_n147,
         LED_RoundFunction0_MCInst1_MC0_n146,
         LED_RoundFunction0_MCInst1_MC0_n145,
         LED_RoundFunction0_MCInst1_MC0_n144,
         LED_RoundFunction0_MCInst1_MC0_n143,
         LED_RoundFunction0_MCInst1_MC0_n142,
         LED_RoundFunction0_MCInst1_MC0_n141,
         LED_RoundFunction0_MCInst1_MC0_n140,
         LED_RoundFunction0_MCInst1_MC0_n139,
         LED_RoundFunction0_MCInst1_MC0_n138,
         LED_RoundFunction0_MCInst1_MC0_n137,
         LED_RoundFunction0_MCInst1_MC0_n136,
         LED_RoundFunction0_MCInst1_MC0_n135,
         LED_RoundFunction0_MCInst1_MC0_n134,
         LED_RoundFunction0_MCInst1_MC0_n133,
         LED_RoundFunction0_MCInst1_MC0_n132,
         LED_RoundFunction0_MCInst1_MC0_n131,
         LED_RoundFunction0_MCInst1_MC0_n130,
         LED_RoundFunction0_MCInst1_MC0_n129,
         LED_RoundFunction0_MCInst1_MC0_n128,
         LED_RoundFunction0_MCInst1_MC0_n127,
         LED_RoundFunction0_MCInst1_MC0_n126,
         LED_RoundFunction0_MCInst1_MC0_n125,
         LED_RoundFunction0_MCInst1_MC0_n124,
         LED_RoundFunction0_MCInst1_MC0_n123,
         LED_RoundFunction0_MCInst1_MC0_n122,
         LED_RoundFunction0_MCInst1_MC0_n121,
         LED_RoundFunction0_MCInst1_MC0_n120,
         LED_RoundFunction0_MCInst1_MC0_n119,
         LED_RoundFunction0_MCInst1_MC0_n118,
         LED_RoundFunction0_MCInst1_MC0_n117,
         LED_RoundFunction0_MCInst1_MC0_n116,
         LED_RoundFunction0_MCInst1_MC0_n115,
         LED_RoundFunction0_MCInst1_MC0_n114,
         LED_RoundFunction0_MCInst1_MC0_n113,
         LED_RoundFunction0_MCInst1_MC0_n112,
         LED_RoundFunction0_MCInst1_MC0_n111,
         LED_RoundFunction0_MCInst1_MC0_n110,
         LED_RoundFunction0_MCInst1_MC0_n109,
         LED_RoundFunction0_MCInst1_MC1_n160,
         LED_RoundFunction0_MCInst1_MC1_n159,
         LED_RoundFunction0_MCInst1_MC1_n158,
         LED_RoundFunction0_MCInst1_MC1_n157,
         LED_RoundFunction0_MCInst1_MC1_n156,
         LED_RoundFunction0_MCInst1_MC1_n155,
         LED_RoundFunction0_MCInst1_MC1_n154,
         LED_RoundFunction0_MCInst1_MC1_n153,
         LED_RoundFunction0_MCInst1_MC1_n152,
         LED_RoundFunction0_MCInst1_MC1_n151,
         LED_RoundFunction0_MCInst1_MC1_n150,
         LED_RoundFunction0_MCInst1_MC1_n149,
         LED_RoundFunction0_MCInst1_MC1_n148,
         LED_RoundFunction0_MCInst1_MC1_n147,
         LED_RoundFunction0_MCInst1_MC1_n146,
         LED_RoundFunction0_MCInst1_MC1_n145,
         LED_RoundFunction0_MCInst1_MC1_n144,
         LED_RoundFunction0_MCInst1_MC1_n143,
         LED_RoundFunction0_MCInst1_MC1_n142,
         LED_RoundFunction0_MCInst1_MC1_n141,
         LED_RoundFunction0_MCInst1_MC1_n140,
         LED_RoundFunction0_MCInst1_MC1_n139,
         LED_RoundFunction0_MCInst1_MC1_n138,
         LED_RoundFunction0_MCInst1_MC1_n137,
         LED_RoundFunction0_MCInst1_MC1_n136,
         LED_RoundFunction0_MCInst1_MC1_n135,
         LED_RoundFunction0_MCInst1_MC1_n134,
         LED_RoundFunction0_MCInst1_MC1_n133,
         LED_RoundFunction0_MCInst1_MC1_n132,
         LED_RoundFunction0_MCInst1_MC1_n131,
         LED_RoundFunction0_MCInst1_MC1_n130,
         LED_RoundFunction0_MCInst1_MC1_n129,
         LED_RoundFunction0_MCInst1_MC1_n128,
         LED_RoundFunction0_MCInst1_MC1_n127,
         LED_RoundFunction0_MCInst1_MC1_n126,
         LED_RoundFunction0_MCInst1_MC1_n125,
         LED_RoundFunction0_MCInst1_MC1_n124,
         LED_RoundFunction0_MCInst1_MC1_n123,
         LED_RoundFunction0_MCInst1_MC1_n122,
         LED_RoundFunction0_MCInst1_MC1_n121,
         LED_RoundFunction0_MCInst1_MC1_n120,
         LED_RoundFunction0_MCInst1_MC1_n119,
         LED_RoundFunction0_MCInst1_MC1_n118,
         LED_RoundFunction0_MCInst1_MC1_n117,
         LED_RoundFunction0_MCInst1_MC1_n116,
         LED_RoundFunction0_MCInst1_MC1_n115,
         LED_RoundFunction0_MCInst1_MC1_n114,
         LED_RoundFunction0_MCInst1_MC1_n113,
         LED_RoundFunction0_MCInst1_MC1_n112,
         LED_RoundFunction0_MCInst1_MC1_n111,
         LED_RoundFunction0_MCInst1_MC1_n110,
         LED_RoundFunction0_MCInst1_MC1_n109,
         LED_RoundFunction0_MCInst1_MC2_n160,
         LED_RoundFunction0_MCInst1_MC2_n159,
         LED_RoundFunction0_MCInst1_MC2_n158,
         LED_RoundFunction0_MCInst1_MC2_n157,
         LED_RoundFunction0_MCInst1_MC2_n156,
         LED_RoundFunction0_MCInst1_MC2_n155,
         LED_RoundFunction0_MCInst1_MC2_n154,
         LED_RoundFunction0_MCInst1_MC2_n153,
         LED_RoundFunction0_MCInst1_MC2_n152,
         LED_RoundFunction0_MCInst1_MC2_n151,
         LED_RoundFunction0_MCInst1_MC2_n150,
         LED_RoundFunction0_MCInst1_MC2_n149,
         LED_RoundFunction0_MCInst1_MC2_n148,
         LED_RoundFunction0_MCInst1_MC2_n147,
         LED_RoundFunction0_MCInst1_MC2_n146,
         LED_RoundFunction0_MCInst1_MC2_n145,
         LED_RoundFunction0_MCInst1_MC2_n144,
         LED_RoundFunction0_MCInst1_MC2_n143,
         LED_RoundFunction0_MCInst1_MC2_n142,
         LED_RoundFunction0_MCInst1_MC2_n141,
         LED_RoundFunction0_MCInst1_MC2_n140,
         LED_RoundFunction0_MCInst1_MC2_n139,
         LED_RoundFunction0_MCInst1_MC2_n138,
         LED_RoundFunction0_MCInst1_MC2_n137,
         LED_RoundFunction0_MCInst1_MC2_n136,
         LED_RoundFunction0_MCInst1_MC2_n135,
         LED_RoundFunction0_MCInst1_MC2_n134,
         LED_RoundFunction0_MCInst1_MC2_n133,
         LED_RoundFunction0_MCInst1_MC2_n132,
         LED_RoundFunction0_MCInst1_MC2_n131,
         LED_RoundFunction0_MCInst1_MC2_n130,
         LED_RoundFunction0_MCInst1_MC2_n129,
         LED_RoundFunction0_MCInst1_MC2_n128,
         LED_RoundFunction0_MCInst1_MC2_n127,
         LED_RoundFunction0_MCInst1_MC2_n126,
         LED_RoundFunction0_MCInst1_MC2_n125,
         LED_RoundFunction0_MCInst1_MC2_n124,
         LED_RoundFunction0_MCInst1_MC2_n123,
         LED_RoundFunction0_MCInst1_MC2_n122,
         LED_RoundFunction0_MCInst1_MC2_n121,
         LED_RoundFunction0_MCInst1_MC2_n120,
         LED_RoundFunction0_MCInst1_MC2_n119,
         LED_RoundFunction0_MCInst1_MC2_n118,
         LED_RoundFunction0_MCInst1_MC2_n117,
         LED_RoundFunction0_MCInst1_MC2_n116,
         LED_RoundFunction0_MCInst1_MC2_n115,
         LED_RoundFunction0_MCInst1_MC2_n114,
         LED_RoundFunction0_MCInst1_MC2_n113,
         LED_RoundFunction0_MCInst1_MC2_n112,
         LED_RoundFunction0_MCInst1_MC2_n111,
         LED_RoundFunction0_MCInst1_MC2_n110,
         LED_RoundFunction0_MCInst1_MC2_n109,
         LED_RoundFunction0_MCInst1_MC3_n160,
         LED_RoundFunction0_MCInst1_MC3_n159,
         LED_RoundFunction0_MCInst1_MC3_n158,
         LED_RoundFunction0_MCInst1_MC3_n157,
         LED_RoundFunction0_MCInst1_MC3_n156,
         LED_RoundFunction0_MCInst1_MC3_n155,
         LED_RoundFunction0_MCInst1_MC3_n154,
         LED_RoundFunction0_MCInst1_MC3_n153,
         LED_RoundFunction0_MCInst1_MC3_n152,
         LED_RoundFunction0_MCInst1_MC3_n151,
         LED_RoundFunction0_MCInst1_MC3_n150,
         LED_RoundFunction0_MCInst1_MC3_n149,
         LED_RoundFunction0_MCInst1_MC3_n148,
         LED_RoundFunction0_MCInst1_MC3_n147,
         LED_RoundFunction0_MCInst1_MC3_n146,
         LED_RoundFunction0_MCInst1_MC3_n145,
         LED_RoundFunction0_MCInst1_MC3_n144,
         LED_RoundFunction0_MCInst1_MC3_n143,
         LED_RoundFunction0_MCInst1_MC3_n142,
         LED_RoundFunction0_MCInst1_MC3_n141,
         LED_RoundFunction0_MCInst1_MC3_n140,
         LED_RoundFunction0_MCInst1_MC3_n139,
         LED_RoundFunction0_MCInst1_MC3_n138,
         LED_RoundFunction0_MCInst1_MC3_n137,
         LED_RoundFunction0_MCInst1_MC3_n136,
         LED_RoundFunction0_MCInst1_MC3_n135,
         LED_RoundFunction0_MCInst1_MC3_n134,
         LED_RoundFunction0_MCInst1_MC3_n133,
         LED_RoundFunction0_MCInst1_MC3_n132,
         LED_RoundFunction0_MCInst1_MC3_n131,
         LED_RoundFunction0_MCInst1_MC3_n130,
         LED_RoundFunction0_MCInst1_MC3_n129,
         LED_RoundFunction0_MCInst1_MC3_n128,
         LED_RoundFunction0_MCInst1_MC3_n127,
         LED_RoundFunction0_MCInst1_MC3_n126,
         LED_RoundFunction0_MCInst1_MC3_n125,
         LED_RoundFunction0_MCInst1_MC3_n124,
         LED_RoundFunction0_MCInst1_MC3_n123,
         LED_RoundFunction0_MCInst1_MC3_n122,
         LED_RoundFunction0_MCInst1_MC3_n121,
         LED_RoundFunction0_MCInst1_MC3_n120,
         LED_RoundFunction0_MCInst1_MC3_n119,
         LED_RoundFunction0_MCInst1_MC3_n118,
         LED_RoundFunction0_MCInst1_MC3_n117,
         LED_RoundFunction0_MCInst1_MC3_n116,
         LED_RoundFunction0_MCInst1_MC3_n115,
         LED_RoundFunction0_MCInst1_MC3_n114,
         LED_RoundFunction0_MCInst1_MC3_n113,
         LED_RoundFunction0_MCInst1_MC3_n112,
         LED_RoundFunction0_MCInst1_MC3_n111,
         LED_RoundFunction0_MCInst1_MC3_n110,
         LED_RoundFunction0_MCInst1_MC3_n109, LED_RoundFunction1_n836,
         LED_RoundFunction1_n835, LED_RoundFunction1_n834,
         LED_RoundFunction1_n833, LED_RoundFunction1_n832,
         LED_RoundFunction1_n831, LED_RoundFunction1_n830,
         LED_RoundFunction1_n829, LED_RoundFunction1_n828,
         LED_RoundFunction1_n827, LED_RoundFunction1_n826,
         LED_RoundFunction1_n825, LED_RoundFunction1_n824,
         LED_RoundFunction1_n823, LED_RoundFunction1_n822,
         LED_RoundFunction1_n821, LED_RoundFunction1_n820,
         LED_RoundFunction1_n819, LED_RoundFunction1_n818,
         LED_RoundFunction1_n817, LED_RoundFunction1_n816,
         LED_RoundFunction1_n815, LED_RoundFunction1_n814,
         LED_RoundFunction1_n813, LED_RoundFunction1_n812,
         LED_RoundFunction1_n811, LED_RoundFunction1_n810,
         LED_RoundFunction1_n809, LED_RoundFunction1_n808,
         LED_RoundFunction1_n807, LED_RoundFunction1_n806,
         LED_RoundFunction1_n805, LED_RoundFunction1_n804,
         LED_RoundFunction1_n803, LED_RoundFunction1_n802,
         LED_RoundFunction1_n801, LED_RoundFunction1_n800,
         LED_RoundFunction1_n799, LED_RoundFunction1_n798,
         LED_RoundFunction1_n797, LED_RoundFunction1_n796,
         LED_RoundFunction1_n795, LED_RoundFunction1_n794,
         LED_RoundFunction1_n793, LED_RoundFunction1_n792,
         LED_RoundFunction1_n791, LED_RoundFunction1_n790,
         LED_RoundFunction1_n789, LED_RoundFunction1_n788,
         LED_RoundFunction1_n787, LED_RoundFunction1_n786,
         LED_RoundFunction1_n785, LED_RoundFunction1_n784,
         LED_RoundFunction1_n783, LED_RoundFunction1_n782,
         LED_RoundFunction1_n781, LED_RoundFunction1_n780,
         LED_RoundFunction1_n779, LED_RoundFunction1_n778,
         LED_RoundFunction1_n777, LED_RoundFunction1_n776,
         LED_RoundFunction1_n775, LED_RoundFunction1_n774,
         LED_RoundFunction1_n773, LED_RoundFunction1_n772,
         LED_RoundFunction1_n771, LED_RoundFunction1_n770,
         LED_RoundFunction1_n769, LED_RoundFunction1_n768,
         LED_RoundFunction1_n767, LED_RoundFunction1_n766,
         LED_RoundFunction1_n765, LED_RoundFunction1_n764,
         LED_RoundFunction1_n763, LED_RoundFunction1_n762,
         LED_RoundFunction1_n761, LED_RoundFunction1_n760,
         LED_RoundFunction1_n759, LED_RoundFunction1_n758,
         LED_RoundFunction1_n757, LED_RoundFunction1_n756,
         LED_RoundFunction1_n755, LED_RoundFunction1_n754,
         LED_RoundFunction1_n753, LED_RoundFunction1_n752,
         LED_RoundFunction1_n751, LED_RoundFunction1_n750,
         LED_RoundFunction1_n749, LED_RoundFunction1_n748,
         LED_RoundFunction1_n747, LED_RoundFunction1_n746,
         LED_RoundFunction1_n745, LED_RoundFunction1_n744,
         LED_RoundFunction1_n743, LED_RoundFunction1_n742,
         LED_RoundFunction1_n741, LED_RoundFunction1_n740,
         LED_RoundFunction1_n739, LED_RoundFunction1_n738,
         LED_RoundFunction1_n737, LED_RoundFunction1_n736,
         LED_RoundFunction1_n735, LED_RoundFunction1_n734,
         LED_RoundFunction1_n733, LED_RoundFunction1_n732,
         LED_RoundFunction1_n731, LED_RoundFunction1_n730,
         LED_RoundFunction1_n729, LED_RoundFunction1_n728,
         LED_RoundFunction1_n727, LED_RoundFunction1_n726,
         LED_RoundFunction1_n725, LED_RoundFunction1_n724,
         LED_RoundFunction1_n723, LED_RoundFunction1_n722,
         LED_RoundFunction1_n721, LED_RoundFunction1_n720,
         LED_RoundFunction1_n719, LED_RoundFunction1_n718,
         LED_RoundFunction1_n717, LED_RoundFunction1_n716,
         LED_RoundFunction1_n715, LED_RoundFunction1_n714,
         LED_RoundFunction1_n713, LED_RoundFunction1_n712,
         LED_RoundFunction1_n711, LED_RoundFunction1_n710,
         LED_RoundFunction1_n709, LED_RoundFunction1_n708,
         LED_RoundFunction1_n707, LED_RoundFunction1_n706,
         LED_RoundFunction1_n705, LED_RoundFunction1_n704,
         LED_RoundFunction1_n703, LED_RoundFunction1_n702,
         LED_RoundFunction1_n701, LED_RoundFunction1_n700,
         LED_RoundFunction1_n699, LED_RoundFunction1_n698,
         LED_RoundFunction1_n697, LED_RoundFunction1_n696,
         LED_RoundFunction1_n695, LED_RoundFunction1_n694,
         LED_RoundFunction1_n693, LED_RoundFunction1_n692,
         LED_RoundFunction1_n691, LED_RoundFunction1_n690,
         LED_RoundFunction1_n689, LED_RoundFunction1_n688,
         LED_RoundFunction1_n687, LED_RoundFunction1_n686,
         LED_RoundFunction1_n685, LED_RoundFunction1_n684,
         LED_RoundFunction1_n683, LED_RoundFunction1_n682,
         LED_RoundFunction1_n681, LED_RoundFunction1_n680,
         LED_RoundFunction1_n679, LED_RoundFunction1_n678,
         LED_RoundFunction1_n677, LED_RoundFunction1_n676,
         LED_RoundFunction1_n675, LED_RoundFunction1_n674,
         LED_RoundFunction1_n673, LED_RoundFunction1_n672,
         LED_RoundFunction1_n671, LED_RoundFunction1_n670,
         LED_RoundFunction1_n669, LED_RoundFunction1_n668,
         LED_RoundFunction1_n667, LED_RoundFunction1_n666,
         LED_RoundFunction1_n665, LED_RoundFunction1_n664,
         LED_RoundFunction1_n663, LED_RoundFunction1_n662,
         LED_RoundFunction1_n661, LED_RoundFunction1_n660,
         LED_RoundFunction1_n659, LED_RoundFunction1_n658,
         LED_RoundFunction1_n657, LED_RoundFunction1_n656,
         LED_RoundFunction1_n655, LED_RoundFunction1_n654,
         LED_RoundFunction1_n653, LED_RoundFunction1_n652,
         LED_RoundFunction1_n651, LED_RoundFunction1_n650,
         LED_RoundFunction1_n649, LED_RoundFunction1_n648,
         LED_RoundFunction1_n647, LED_RoundFunction1_n646,
         LED_RoundFunction1_n645, LED_RoundFunction1_n644,
         LED_RoundFunction1_n643, LED_RoundFunction1_n642,
         LED_RoundFunction1_n641, LED_RoundFunction1_n640,
         LED_RoundFunction1_n639, LED_RoundFunction1_n638,
         LED_RoundFunction1_n637, LED_RoundFunction1_n636,
         LED_RoundFunction1_n635, LED_RoundFunction1_n634,
         LED_RoundFunction1_n633, LED_RoundFunction1_n632,
         LED_RoundFunction1_n631, LED_RoundFunction1_n630,
         LED_RoundFunction1_n629, LED_RoundFunction1_n628,
         LED_RoundFunction1_n627, LED_RoundFunction1_n626,
         LED_RoundFunction1_n625, LED_RoundFunction1_n624,
         LED_RoundFunction1_n623, LED_RoundFunction1_n622,
         LED_RoundFunction1_n621, LED_RoundFunction1_n620,
         LED_RoundFunction1_n619, LED_RoundFunction1_n618,
         LED_RoundFunction1_n617, LED_RoundFunction1_n616,
         LED_RoundFunction1_n615, LED_RoundFunction1_n614,
         LED_RoundFunction1_n613, LED_RoundFunction1_n612,
         LED_RoundFunction1_n611, LED_RoundFunction1_n610,
         LED_RoundFunction1_n609, LED_RoundFunction1_n608,
         LED_RoundFunction1_n607, LED_RoundFunction1_n606,
         LED_RoundFunction1_n605, LED_RoundFunction1_n604,
         LED_RoundFunction1_n603, LED_RoundFunction1_n602,
         LED_RoundFunction1_n601, LED_RoundFunction1_n600,
         LED_RoundFunction1_n599, LED_RoundFunction1_n598,
         LED_RoundFunction1_n597, LED_RoundFunction1_n596,
         LED_RoundFunction1_n595, LED_RoundFunction1_n594,
         LED_RoundFunction1_n593, LED_RoundFunction1_n592,
         LED_RoundFunction1_n591, LED_RoundFunction1_n590,
         LED_RoundFunction1_n589, LED_RoundFunction1_n588,
         LED_RoundFunction1_n587, LED_RoundFunction1_n586,
         LED_RoundFunction1_n585, LED_RoundFunction1_n584,
         LED_RoundFunction1_n583, LED_RoundFunction1_n582,
         LED_RoundFunction1_n581, LED_RoundFunction1_n580,
         LED_RoundFunction1_n579, LED_RoundFunction1_n578,
         LED_RoundFunction1_n577, LED_RoundFunction1_n576,
         LED_RoundFunction1_n575, LED_RoundFunction1_n574,
         LED_RoundFunction1_n573, LED_RoundFunction1_n572,
         LED_RoundFunction1_n571, LED_RoundFunction1_n570,
         LED_RoundFunction1_n569, LED_RoundFunction1_n568,
         LED_RoundFunction1_n567, LED_RoundFunction1_n566,
         LED_RoundFunction1_n565, LED_RoundFunction1_n564,
         LED_RoundFunction1_n563, LED_RoundFunction1_n562,
         LED_RoundFunction1_n561, LED_RoundFunction1_n560,
         LED_RoundFunction1_n559, LED_RoundFunction1_n558,
         LED_RoundFunction1_n557, LED_RoundFunction1_n556,
         LED_RoundFunction1_n555, LED_RoundFunction1_Feedback_0_,
         LED_RoundFunction1_Feedback_1_, LED_RoundFunction1_Feedback_2_,
         LED_RoundFunction1_Feedback_3_, LED_RoundFunction1_Feedback_4_,
         LED_RoundFunction1_Feedback_5_, LED_RoundFunction1_Feedback_6_,
         LED_RoundFunction1_Feedback_7_, LED_RoundFunction1_Feedback_8_,
         LED_RoundFunction1_Feedback_9_, LED_RoundFunction1_Feedback_10_,
         LED_RoundFunction1_Feedback_11_, LED_RoundFunction1_Feedback_12_,
         LED_RoundFunction1_Feedback_13_, LED_RoundFunction1_Feedback_14_,
         LED_RoundFunction1_Feedback_15_, LED_RoundFunction1_Feedback_16_,
         LED_RoundFunction1_Feedback_17_, LED_RoundFunction1_Feedback_18_,
         LED_RoundFunction1_Feedback_19_, LED_RoundFunction1_Feedback_20_,
         LED_RoundFunction1_Feedback_21_, LED_RoundFunction1_Feedback_22_,
         LED_RoundFunction1_Feedback_23_, LED_RoundFunction1_Feedback_24_,
         LED_RoundFunction1_Feedback_25_, LED_RoundFunction1_Feedback_26_,
         LED_RoundFunction1_Feedback_27_, LED_RoundFunction1_Feedback_28_,
         LED_RoundFunction1_Feedback_29_, LED_RoundFunction1_Feedback_30_,
         LED_RoundFunction1_Feedback_31_, LED_RoundFunction1_Feedback_32_,
         LED_RoundFunction1_Feedback_33_, LED_RoundFunction1_Feedback_34_,
         LED_RoundFunction1_Feedback_35_, LED_RoundFunction1_Feedback_36_,
         LED_RoundFunction1_Feedback_37_, LED_RoundFunction1_Feedback_38_,
         LED_RoundFunction1_Feedback_39_, LED_RoundFunction1_Feedback_40_,
         LED_RoundFunction1_Feedback_41_, LED_RoundFunction1_Feedback_42_,
         LED_RoundFunction1_Feedback_43_, LED_RoundFunction1_Feedback_44_,
         LED_RoundFunction1_Feedback_45_, LED_RoundFunction1_Feedback_46_,
         LED_RoundFunction1_Feedback_47_, LED_RoundFunction1_Feedback_48_,
         LED_RoundFunction1_Feedback_49_, LED_RoundFunction1_Feedback_50_,
         LED_RoundFunction1_Feedback_51_, LED_RoundFunction1_Feedback_52_,
         LED_RoundFunction1_Feedback_53_, LED_RoundFunction1_Feedback_54_,
         LED_RoundFunction1_Feedback_55_, LED_RoundFunction1_Feedback_56_,
         LED_RoundFunction1_Feedback_57_, LED_RoundFunction1_Feedback_58_,
         LED_RoundFunction1_Feedback_59_, LED_RoundFunction1_Feedback_60_,
         LED_RoundFunction1_Feedback_61_, LED_RoundFunction1_Feedback_62_,
         LED_RoundFunction1_Feedback_63_, LED_RoundFunction1_MCInst1_MC0_n160,
         LED_RoundFunction1_MCInst1_MC0_n159,
         LED_RoundFunction1_MCInst1_MC0_n158,
         LED_RoundFunction1_MCInst1_MC0_n157,
         LED_RoundFunction1_MCInst1_MC0_n156,
         LED_RoundFunction1_MCInst1_MC0_n155,
         LED_RoundFunction1_MCInst1_MC0_n154,
         LED_RoundFunction1_MCInst1_MC0_n153,
         LED_RoundFunction1_MCInst1_MC0_n152,
         LED_RoundFunction1_MCInst1_MC0_n151,
         LED_RoundFunction1_MCInst1_MC0_n150,
         LED_RoundFunction1_MCInst1_MC0_n149,
         LED_RoundFunction1_MCInst1_MC0_n148,
         LED_RoundFunction1_MCInst1_MC0_n147,
         LED_RoundFunction1_MCInst1_MC0_n146,
         LED_RoundFunction1_MCInst1_MC0_n145,
         LED_RoundFunction1_MCInst1_MC0_n144,
         LED_RoundFunction1_MCInst1_MC0_n143,
         LED_RoundFunction1_MCInst1_MC0_n142,
         LED_RoundFunction1_MCInst1_MC0_n141,
         LED_RoundFunction1_MCInst1_MC0_n140,
         LED_RoundFunction1_MCInst1_MC0_n139,
         LED_RoundFunction1_MCInst1_MC0_n138,
         LED_RoundFunction1_MCInst1_MC0_n137,
         LED_RoundFunction1_MCInst1_MC0_n136,
         LED_RoundFunction1_MCInst1_MC0_n135,
         LED_RoundFunction1_MCInst1_MC0_n134,
         LED_RoundFunction1_MCInst1_MC0_n133,
         LED_RoundFunction1_MCInst1_MC0_n132,
         LED_RoundFunction1_MCInst1_MC0_n131,
         LED_RoundFunction1_MCInst1_MC0_n130,
         LED_RoundFunction1_MCInst1_MC0_n129,
         LED_RoundFunction1_MCInst1_MC0_n128,
         LED_RoundFunction1_MCInst1_MC0_n127,
         LED_RoundFunction1_MCInst1_MC0_n126,
         LED_RoundFunction1_MCInst1_MC0_n125,
         LED_RoundFunction1_MCInst1_MC0_n124,
         LED_RoundFunction1_MCInst1_MC0_n123,
         LED_RoundFunction1_MCInst1_MC0_n122,
         LED_RoundFunction1_MCInst1_MC0_n121,
         LED_RoundFunction1_MCInst1_MC0_n120,
         LED_RoundFunction1_MCInst1_MC0_n119,
         LED_RoundFunction1_MCInst1_MC0_n118,
         LED_RoundFunction1_MCInst1_MC0_n117,
         LED_RoundFunction1_MCInst1_MC0_n116,
         LED_RoundFunction1_MCInst1_MC0_n115,
         LED_RoundFunction1_MCInst1_MC0_n114,
         LED_RoundFunction1_MCInst1_MC0_n113,
         LED_RoundFunction1_MCInst1_MC0_n112,
         LED_RoundFunction1_MCInst1_MC0_n111,
         LED_RoundFunction1_MCInst1_MC0_n110,
         LED_RoundFunction1_MCInst1_MC0_n109,
         LED_RoundFunction1_MCInst1_MC1_n160,
         LED_RoundFunction1_MCInst1_MC1_n159,
         LED_RoundFunction1_MCInst1_MC1_n158,
         LED_RoundFunction1_MCInst1_MC1_n157,
         LED_RoundFunction1_MCInst1_MC1_n156,
         LED_RoundFunction1_MCInst1_MC1_n155,
         LED_RoundFunction1_MCInst1_MC1_n154,
         LED_RoundFunction1_MCInst1_MC1_n153,
         LED_RoundFunction1_MCInst1_MC1_n152,
         LED_RoundFunction1_MCInst1_MC1_n151,
         LED_RoundFunction1_MCInst1_MC1_n150,
         LED_RoundFunction1_MCInst1_MC1_n149,
         LED_RoundFunction1_MCInst1_MC1_n148,
         LED_RoundFunction1_MCInst1_MC1_n147,
         LED_RoundFunction1_MCInst1_MC1_n146,
         LED_RoundFunction1_MCInst1_MC1_n145,
         LED_RoundFunction1_MCInst1_MC1_n144,
         LED_RoundFunction1_MCInst1_MC1_n143,
         LED_RoundFunction1_MCInst1_MC1_n142,
         LED_RoundFunction1_MCInst1_MC1_n141,
         LED_RoundFunction1_MCInst1_MC1_n140,
         LED_RoundFunction1_MCInst1_MC1_n139,
         LED_RoundFunction1_MCInst1_MC1_n138,
         LED_RoundFunction1_MCInst1_MC1_n137,
         LED_RoundFunction1_MCInst1_MC1_n136,
         LED_RoundFunction1_MCInst1_MC1_n135,
         LED_RoundFunction1_MCInst1_MC1_n134,
         LED_RoundFunction1_MCInst1_MC1_n133,
         LED_RoundFunction1_MCInst1_MC1_n132,
         LED_RoundFunction1_MCInst1_MC1_n131,
         LED_RoundFunction1_MCInst1_MC1_n130,
         LED_RoundFunction1_MCInst1_MC1_n129,
         LED_RoundFunction1_MCInst1_MC1_n128,
         LED_RoundFunction1_MCInst1_MC1_n127,
         LED_RoundFunction1_MCInst1_MC1_n126,
         LED_RoundFunction1_MCInst1_MC1_n125,
         LED_RoundFunction1_MCInst1_MC1_n124,
         LED_RoundFunction1_MCInst1_MC1_n123,
         LED_RoundFunction1_MCInst1_MC1_n122,
         LED_RoundFunction1_MCInst1_MC1_n121,
         LED_RoundFunction1_MCInst1_MC1_n120,
         LED_RoundFunction1_MCInst1_MC1_n119,
         LED_RoundFunction1_MCInst1_MC1_n118,
         LED_RoundFunction1_MCInst1_MC1_n117,
         LED_RoundFunction1_MCInst1_MC1_n116,
         LED_RoundFunction1_MCInst1_MC1_n115,
         LED_RoundFunction1_MCInst1_MC1_n114,
         LED_RoundFunction1_MCInst1_MC1_n113,
         LED_RoundFunction1_MCInst1_MC1_n112,
         LED_RoundFunction1_MCInst1_MC1_n111,
         LED_RoundFunction1_MCInst1_MC1_n110,
         LED_RoundFunction1_MCInst1_MC1_n109,
         LED_RoundFunction1_MCInst1_MC2_n160,
         LED_RoundFunction1_MCInst1_MC2_n159,
         LED_RoundFunction1_MCInst1_MC2_n158,
         LED_RoundFunction1_MCInst1_MC2_n157,
         LED_RoundFunction1_MCInst1_MC2_n156,
         LED_RoundFunction1_MCInst1_MC2_n155,
         LED_RoundFunction1_MCInst1_MC2_n154,
         LED_RoundFunction1_MCInst1_MC2_n153,
         LED_RoundFunction1_MCInst1_MC2_n152,
         LED_RoundFunction1_MCInst1_MC2_n151,
         LED_RoundFunction1_MCInst1_MC2_n150,
         LED_RoundFunction1_MCInst1_MC2_n149,
         LED_RoundFunction1_MCInst1_MC2_n148,
         LED_RoundFunction1_MCInst1_MC2_n147,
         LED_RoundFunction1_MCInst1_MC2_n146,
         LED_RoundFunction1_MCInst1_MC2_n145,
         LED_RoundFunction1_MCInst1_MC2_n144,
         LED_RoundFunction1_MCInst1_MC2_n143,
         LED_RoundFunction1_MCInst1_MC2_n142,
         LED_RoundFunction1_MCInst1_MC2_n141,
         LED_RoundFunction1_MCInst1_MC2_n140,
         LED_RoundFunction1_MCInst1_MC2_n139,
         LED_RoundFunction1_MCInst1_MC2_n138,
         LED_RoundFunction1_MCInst1_MC2_n137,
         LED_RoundFunction1_MCInst1_MC2_n136,
         LED_RoundFunction1_MCInst1_MC2_n135,
         LED_RoundFunction1_MCInst1_MC2_n134,
         LED_RoundFunction1_MCInst1_MC2_n133,
         LED_RoundFunction1_MCInst1_MC2_n132,
         LED_RoundFunction1_MCInst1_MC2_n131,
         LED_RoundFunction1_MCInst1_MC2_n130,
         LED_RoundFunction1_MCInst1_MC2_n129,
         LED_RoundFunction1_MCInst1_MC2_n128,
         LED_RoundFunction1_MCInst1_MC2_n127,
         LED_RoundFunction1_MCInst1_MC2_n126,
         LED_RoundFunction1_MCInst1_MC2_n125,
         LED_RoundFunction1_MCInst1_MC2_n124,
         LED_RoundFunction1_MCInst1_MC2_n123,
         LED_RoundFunction1_MCInst1_MC2_n122,
         LED_RoundFunction1_MCInst1_MC2_n121,
         LED_RoundFunction1_MCInst1_MC2_n120,
         LED_RoundFunction1_MCInst1_MC2_n119,
         LED_RoundFunction1_MCInst1_MC2_n118,
         LED_RoundFunction1_MCInst1_MC2_n117,
         LED_RoundFunction1_MCInst1_MC2_n116,
         LED_RoundFunction1_MCInst1_MC2_n115,
         LED_RoundFunction1_MCInst1_MC2_n114,
         LED_RoundFunction1_MCInst1_MC2_n113,
         LED_RoundFunction1_MCInst1_MC2_n112,
         LED_RoundFunction1_MCInst1_MC2_n111,
         LED_RoundFunction1_MCInst1_MC2_n110,
         LED_RoundFunction1_MCInst1_MC2_n109,
         LED_RoundFunction1_MCInst1_MC3_n160,
         LED_RoundFunction1_MCInst1_MC3_n159,
         LED_RoundFunction1_MCInst1_MC3_n158,
         LED_RoundFunction1_MCInst1_MC3_n157,
         LED_RoundFunction1_MCInst1_MC3_n156,
         LED_RoundFunction1_MCInst1_MC3_n155,
         LED_RoundFunction1_MCInst1_MC3_n154,
         LED_RoundFunction1_MCInst1_MC3_n153,
         LED_RoundFunction1_MCInst1_MC3_n152,
         LED_RoundFunction1_MCInst1_MC3_n151,
         LED_RoundFunction1_MCInst1_MC3_n150,
         LED_RoundFunction1_MCInst1_MC3_n149,
         LED_RoundFunction1_MCInst1_MC3_n148,
         LED_RoundFunction1_MCInst1_MC3_n147,
         LED_RoundFunction1_MCInst1_MC3_n146,
         LED_RoundFunction1_MCInst1_MC3_n145,
         LED_RoundFunction1_MCInst1_MC3_n144,
         LED_RoundFunction1_MCInst1_MC3_n143,
         LED_RoundFunction1_MCInst1_MC3_n142,
         LED_RoundFunction1_MCInst1_MC3_n141,
         LED_RoundFunction1_MCInst1_MC3_n140,
         LED_RoundFunction1_MCInst1_MC3_n139,
         LED_RoundFunction1_MCInst1_MC3_n138,
         LED_RoundFunction1_MCInst1_MC3_n137,
         LED_RoundFunction1_MCInst1_MC3_n136,
         LED_RoundFunction1_MCInst1_MC3_n135,
         LED_RoundFunction1_MCInst1_MC3_n134,
         LED_RoundFunction1_MCInst1_MC3_n133,
         LED_RoundFunction1_MCInst1_MC3_n132,
         LED_RoundFunction1_MCInst1_MC3_n131,
         LED_RoundFunction1_MCInst1_MC3_n130,
         LED_RoundFunction1_MCInst1_MC3_n129,
         LED_RoundFunction1_MCInst1_MC3_n128,
         LED_RoundFunction1_MCInst1_MC3_n127,
         LED_RoundFunction1_MCInst1_MC3_n126,
         LED_RoundFunction1_MCInst1_MC3_n125,
         LED_RoundFunction1_MCInst1_MC3_n124,
         LED_RoundFunction1_MCInst1_MC3_n123,
         LED_RoundFunction1_MCInst1_MC3_n122,
         LED_RoundFunction1_MCInst1_MC3_n121,
         LED_RoundFunction1_MCInst1_MC3_n120,
         LED_RoundFunction1_MCInst1_MC3_n119,
         LED_RoundFunction1_MCInst1_MC3_n118,
         LED_RoundFunction1_MCInst1_MC3_n117,
         LED_RoundFunction1_MCInst1_MC3_n116,
         LED_RoundFunction1_MCInst1_MC3_n115,
         LED_RoundFunction1_MCInst1_MC3_n114,
         LED_RoundFunction1_MCInst1_MC3_n113,
         LED_RoundFunction1_MCInst1_MC3_n112,
         LED_RoundFunction1_MCInst1_MC3_n111,
         LED_RoundFunction1_MCInst1_MC3_n110,
         LED_RoundFunction1_MCInst1_MC3_n109, LED_RoundFunction2_n836,
         LED_RoundFunction2_n835, LED_RoundFunction2_n834,
         LED_RoundFunction2_n833, LED_RoundFunction2_n832,
         LED_RoundFunction2_n831, LED_RoundFunction2_n830,
         LED_RoundFunction2_n829, LED_RoundFunction2_n828,
         LED_RoundFunction2_n827, LED_RoundFunction2_n826,
         LED_RoundFunction2_n825, LED_RoundFunction2_n824,
         LED_RoundFunction2_n823, LED_RoundFunction2_n822,
         LED_RoundFunction2_n821, LED_RoundFunction2_n820,
         LED_RoundFunction2_n819, LED_RoundFunction2_n818,
         LED_RoundFunction2_n817, LED_RoundFunction2_n816,
         LED_RoundFunction2_n815, LED_RoundFunction2_n814,
         LED_RoundFunction2_n813, LED_RoundFunction2_n812,
         LED_RoundFunction2_n811, LED_RoundFunction2_n810,
         LED_RoundFunction2_n809, LED_RoundFunction2_n808,
         LED_RoundFunction2_n807, LED_RoundFunction2_n806,
         LED_RoundFunction2_n805, LED_RoundFunction2_n804,
         LED_RoundFunction2_n803, LED_RoundFunction2_n802,
         LED_RoundFunction2_n801, LED_RoundFunction2_n800,
         LED_RoundFunction2_n799, LED_RoundFunction2_n798,
         LED_RoundFunction2_n797, LED_RoundFunction2_n796,
         LED_RoundFunction2_n795, LED_RoundFunction2_n794,
         LED_RoundFunction2_n793, LED_RoundFunction2_n792,
         LED_RoundFunction2_n791, LED_RoundFunction2_n790,
         LED_RoundFunction2_n789, LED_RoundFunction2_n788,
         LED_RoundFunction2_n787, LED_RoundFunction2_n786,
         LED_RoundFunction2_n785, LED_RoundFunction2_n784,
         LED_RoundFunction2_n783, LED_RoundFunction2_n782,
         LED_RoundFunction2_n781, LED_RoundFunction2_n780,
         LED_RoundFunction2_n779, LED_RoundFunction2_n778,
         LED_RoundFunction2_n777, LED_RoundFunction2_n776,
         LED_RoundFunction2_n775, LED_RoundFunction2_n774,
         LED_RoundFunction2_n773, LED_RoundFunction2_n772,
         LED_RoundFunction2_n771, LED_RoundFunction2_n770,
         LED_RoundFunction2_n769, LED_RoundFunction2_n768,
         LED_RoundFunction2_n767, LED_RoundFunction2_n766,
         LED_RoundFunction2_n765, LED_RoundFunction2_n764,
         LED_RoundFunction2_n763, LED_RoundFunction2_n762,
         LED_RoundFunction2_n761, LED_RoundFunction2_n760,
         LED_RoundFunction2_n759, LED_RoundFunction2_n758,
         LED_RoundFunction2_n757, LED_RoundFunction2_n756,
         LED_RoundFunction2_n755, LED_RoundFunction2_n754,
         LED_RoundFunction2_n753, LED_RoundFunction2_n752,
         LED_RoundFunction2_n751, LED_RoundFunction2_n750,
         LED_RoundFunction2_n749, LED_RoundFunction2_n748,
         LED_RoundFunction2_n747, LED_RoundFunction2_n746,
         LED_RoundFunction2_n745, LED_RoundFunction2_n744,
         LED_RoundFunction2_n743, LED_RoundFunction2_n742,
         LED_RoundFunction2_n741, LED_RoundFunction2_n740,
         LED_RoundFunction2_n739, LED_RoundFunction2_n738,
         LED_RoundFunction2_n737, LED_RoundFunction2_n736,
         LED_RoundFunction2_n735, LED_RoundFunction2_n734,
         LED_RoundFunction2_n733, LED_RoundFunction2_n732,
         LED_RoundFunction2_n731, LED_RoundFunction2_n730,
         LED_RoundFunction2_n729, LED_RoundFunction2_n728,
         LED_RoundFunction2_n727, LED_RoundFunction2_n726,
         LED_RoundFunction2_n725, LED_RoundFunction2_n724,
         LED_RoundFunction2_n723, LED_RoundFunction2_n722,
         LED_RoundFunction2_n721, LED_RoundFunction2_n720,
         LED_RoundFunction2_n719, LED_RoundFunction2_n718,
         LED_RoundFunction2_n717, LED_RoundFunction2_n716,
         LED_RoundFunction2_n715, LED_RoundFunction2_n714,
         LED_RoundFunction2_n713, LED_RoundFunction2_n712,
         LED_RoundFunction2_n711, LED_RoundFunction2_n710,
         LED_RoundFunction2_n709, LED_RoundFunction2_n708,
         LED_RoundFunction2_n707, LED_RoundFunction2_n706,
         LED_RoundFunction2_n705, LED_RoundFunction2_n704,
         LED_RoundFunction2_n703, LED_RoundFunction2_n702,
         LED_RoundFunction2_n701, LED_RoundFunction2_n700,
         LED_RoundFunction2_n699, LED_RoundFunction2_n698,
         LED_RoundFunction2_n697, LED_RoundFunction2_n696,
         LED_RoundFunction2_n695, LED_RoundFunction2_n694,
         LED_RoundFunction2_n693, LED_RoundFunction2_n692,
         LED_RoundFunction2_n691, LED_RoundFunction2_n690,
         LED_RoundFunction2_n689, LED_RoundFunction2_n688,
         LED_RoundFunction2_n687, LED_RoundFunction2_n686,
         LED_RoundFunction2_n685, LED_RoundFunction2_n684,
         LED_RoundFunction2_n683, LED_RoundFunction2_n682,
         LED_RoundFunction2_n681, LED_RoundFunction2_n680,
         LED_RoundFunction2_n679, LED_RoundFunction2_n678,
         LED_RoundFunction2_n677, LED_RoundFunction2_n676,
         LED_RoundFunction2_n675, LED_RoundFunction2_n674,
         LED_RoundFunction2_n673, LED_RoundFunction2_n672,
         LED_RoundFunction2_n671, LED_RoundFunction2_n670,
         LED_RoundFunction2_n669, LED_RoundFunction2_n668,
         LED_RoundFunction2_n667, LED_RoundFunction2_n666,
         LED_RoundFunction2_n665, LED_RoundFunction2_n664,
         LED_RoundFunction2_n663, LED_RoundFunction2_n662,
         LED_RoundFunction2_n661, LED_RoundFunction2_n660,
         LED_RoundFunction2_n659, LED_RoundFunction2_n658,
         LED_RoundFunction2_n657, LED_RoundFunction2_n656,
         LED_RoundFunction2_n655, LED_RoundFunction2_n654,
         LED_RoundFunction2_n653, LED_RoundFunction2_n652,
         LED_RoundFunction2_n651, LED_RoundFunction2_n650,
         LED_RoundFunction2_n649, LED_RoundFunction2_n648,
         LED_RoundFunction2_n647, LED_RoundFunction2_n646,
         LED_RoundFunction2_n645, LED_RoundFunction2_n644,
         LED_RoundFunction2_n643, LED_RoundFunction2_n642,
         LED_RoundFunction2_n641, LED_RoundFunction2_n640,
         LED_RoundFunction2_n639, LED_RoundFunction2_n638,
         LED_RoundFunction2_n637, LED_RoundFunction2_n636,
         LED_RoundFunction2_n635, LED_RoundFunction2_n634,
         LED_RoundFunction2_n633, LED_RoundFunction2_n632,
         LED_RoundFunction2_n631, LED_RoundFunction2_n630,
         LED_RoundFunction2_n629, LED_RoundFunction2_n628,
         LED_RoundFunction2_n627, LED_RoundFunction2_n626,
         LED_RoundFunction2_n625, LED_RoundFunction2_n624,
         LED_RoundFunction2_n623, LED_RoundFunction2_n622,
         LED_RoundFunction2_n621, LED_RoundFunction2_n620,
         LED_RoundFunction2_n619, LED_RoundFunction2_n618,
         LED_RoundFunction2_n617, LED_RoundFunction2_n616,
         LED_RoundFunction2_n615, LED_RoundFunction2_n614,
         LED_RoundFunction2_n613, LED_RoundFunction2_n612,
         LED_RoundFunction2_n611, LED_RoundFunction2_n610,
         LED_RoundFunction2_n609, LED_RoundFunction2_n608,
         LED_RoundFunction2_n607, LED_RoundFunction2_n606,
         LED_RoundFunction2_n605, LED_RoundFunction2_n604,
         LED_RoundFunction2_n603, LED_RoundFunction2_n602,
         LED_RoundFunction2_n601, LED_RoundFunction2_n600,
         LED_RoundFunction2_n599, LED_RoundFunction2_n598,
         LED_RoundFunction2_n597, LED_RoundFunction2_n596,
         LED_RoundFunction2_n595, LED_RoundFunction2_n594,
         LED_RoundFunction2_n593, LED_RoundFunction2_n592,
         LED_RoundFunction2_n591, LED_RoundFunction2_n590,
         LED_RoundFunction2_n589, LED_RoundFunction2_n588,
         LED_RoundFunction2_n587, LED_RoundFunction2_n586,
         LED_RoundFunction2_n585, LED_RoundFunction2_n584,
         LED_RoundFunction2_n583, LED_RoundFunction2_n582,
         LED_RoundFunction2_n581, LED_RoundFunction2_n580,
         LED_RoundFunction2_n579, LED_RoundFunction2_n578,
         LED_RoundFunction2_n577, LED_RoundFunction2_n576,
         LED_RoundFunction2_n575, LED_RoundFunction2_n574,
         LED_RoundFunction2_n573, LED_RoundFunction2_n572,
         LED_RoundFunction2_n571, LED_RoundFunction2_n570,
         LED_RoundFunction2_n569, LED_RoundFunction2_n568,
         LED_RoundFunction2_n567, LED_RoundFunction2_n566,
         LED_RoundFunction2_n565, LED_RoundFunction2_n564,
         LED_RoundFunction2_n563, LED_RoundFunction2_n562,
         LED_RoundFunction2_n561, LED_RoundFunction2_n560,
         LED_RoundFunction2_n559, LED_RoundFunction2_n558,
         LED_RoundFunction2_n557, LED_RoundFunction2_n556,
         LED_RoundFunction2_n555, LED_RoundFunction2_Feedback_0_,
         LED_RoundFunction2_Feedback_1_, LED_RoundFunction2_Feedback_2_,
         LED_RoundFunction2_Feedback_3_, LED_RoundFunction2_Feedback_4_,
         LED_RoundFunction2_Feedback_5_, LED_RoundFunction2_Feedback_6_,
         LED_RoundFunction2_Feedback_7_, LED_RoundFunction2_Feedback_8_,
         LED_RoundFunction2_Feedback_9_, LED_RoundFunction2_Feedback_10_,
         LED_RoundFunction2_Feedback_11_, LED_RoundFunction2_Feedback_12_,
         LED_RoundFunction2_Feedback_13_, LED_RoundFunction2_Feedback_14_,
         LED_RoundFunction2_Feedback_15_, LED_RoundFunction2_Feedback_16_,
         LED_RoundFunction2_Feedback_17_, LED_RoundFunction2_Feedback_18_,
         LED_RoundFunction2_Feedback_19_, LED_RoundFunction2_Feedback_20_,
         LED_RoundFunction2_Feedback_21_, LED_RoundFunction2_Feedback_22_,
         LED_RoundFunction2_Feedback_23_, LED_RoundFunction2_Feedback_24_,
         LED_RoundFunction2_Feedback_25_, LED_RoundFunction2_Feedback_26_,
         LED_RoundFunction2_Feedback_27_, LED_RoundFunction2_Feedback_28_,
         LED_RoundFunction2_Feedback_29_, LED_RoundFunction2_Feedback_30_,
         LED_RoundFunction2_Feedback_31_, LED_RoundFunction2_Feedback_32_,
         LED_RoundFunction2_Feedback_33_, LED_RoundFunction2_Feedback_34_,
         LED_RoundFunction2_Feedback_35_, LED_RoundFunction2_Feedback_36_,
         LED_RoundFunction2_Feedback_37_, LED_RoundFunction2_Feedback_38_,
         LED_RoundFunction2_Feedback_39_, LED_RoundFunction2_Feedback_40_,
         LED_RoundFunction2_Feedback_41_, LED_RoundFunction2_Feedback_42_,
         LED_RoundFunction2_Feedback_43_, LED_RoundFunction2_Feedback_44_,
         LED_RoundFunction2_Feedback_45_, LED_RoundFunction2_Feedback_46_,
         LED_RoundFunction2_Feedback_47_, LED_RoundFunction2_Feedback_48_,
         LED_RoundFunction2_Feedback_49_, LED_RoundFunction2_Feedback_50_,
         LED_RoundFunction2_Feedback_51_, LED_RoundFunction2_Feedback_52_,
         LED_RoundFunction2_Feedback_53_, LED_RoundFunction2_Feedback_54_,
         LED_RoundFunction2_Feedback_55_, LED_RoundFunction2_Feedback_56_,
         LED_RoundFunction2_Feedback_57_, LED_RoundFunction2_Feedback_58_,
         LED_RoundFunction2_Feedback_59_, LED_RoundFunction2_Feedback_60_,
         LED_RoundFunction2_Feedback_61_, LED_RoundFunction2_Feedback_62_,
         LED_RoundFunction2_Feedback_63_, LED_RoundFunction2_MCInst1_MC0_n160,
         LED_RoundFunction2_MCInst1_MC0_n159,
         LED_RoundFunction2_MCInst1_MC0_n158,
         LED_RoundFunction2_MCInst1_MC0_n157,
         LED_RoundFunction2_MCInst1_MC0_n156,
         LED_RoundFunction2_MCInst1_MC0_n155,
         LED_RoundFunction2_MCInst1_MC0_n154,
         LED_RoundFunction2_MCInst1_MC0_n153,
         LED_RoundFunction2_MCInst1_MC0_n152,
         LED_RoundFunction2_MCInst1_MC0_n151,
         LED_RoundFunction2_MCInst1_MC0_n150,
         LED_RoundFunction2_MCInst1_MC0_n149,
         LED_RoundFunction2_MCInst1_MC0_n148,
         LED_RoundFunction2_MCInst1_MC0_n147,
         LED_RoundFunction2_MCInst1_MC0_n146,
         LED_RoundFunction2_MCInst1_MC0_n145,
         LED_RoundFunction2_MCInst1_MC0_n144,
         LED_RoundFunction2_MCInst1_MC0_n143,
         LED_RoundFunction2_MCInst1_MC0_n142,
         LED_RoundFunction2_MCInst1_MC0_n141,
         LED_RoundFunction2_MCInst1_MC0_n140,
         LED_RoundFunction2_MCInst1_MC0_n139,
         LED_RoundFunction2_MCInst1_MC0_n138,
         LED_RoundFunction2_MCInst1_MC0_n137,
         LED_RoundFunction2_MCInst1_MC0_n136,
         LED_RoundFunction2_MCInst1_MC0_n135,
         LED_RoundFunction2_MCInst1_MC0_n134,
         LED_RoundFunction2_MCInst1_MC0_n133,
         LED_RoundFunction2_MCInst1_MC0_n132,
         LED_RoundFunction2_MCInst1_MC0_n131,
         LED_RoundFunction2_MCInst1_MC0_n130,
         LED_RoundFunction2_MCInst1_MC0_n129,
         LED_RoundFunction2_MCInst1_MC0_n128,
         LED_RoundFunction2_MCInst1_MC0_n127,
         LED_RoundFunction2_MCInst1_MC0_n126,
         LED_RoundFunction2_MCInst1_MC0_n125,
         LED_RoundFunction2_MCInst1_MC0_n124,
         LED_RoundFunction2_MCInst1_MC0_n123,
         LED_RoundFunction2_MCInst1_MC0_n122,
         LED_RoundFunction2_MCInst1_MC0_n121,
         LED_RoundFunction2_MCInst1_MC0_n120,
         LED_RoundFunction2_MCInst1_MC0_n119,
         LED_RoundFunction2_MCInst1_MC0_n118,
         LED_RoundFunction2_MCInst1_MC0_n117,
         LED_RoundFunction2_MCInst1_MC0_n116,
         LED_RoundFunction2_MCInst1_MC0_n115,
         LED_RoundFunction2_MCInst1_MC0_n114,
         LED_RoundFunction2_MCInst1_MC0_n113,
         LED_RoundFunction2_MCInst1_MC0_n112,
         LED_RoundFunction2_MCInst1_MC0_n111,
         LED_RoundFunction2_MCInst1_MC0_n110,
         LED_RoundFunction2_MCInst1_MC0_n109,
         LED_RoundFunction2_MCInst1_MC1_n160,
         LED_RoundFunction2_MCInst1_MC1_n159,
         LED_RoundFunction2_MCInst1_MC1_n158,
         LED_RoundFunction2_MCInst1_MC1_n157,
         LED_RoundFunction2_MCInst1_MC1_n156,
         LED_RoundFunction2_MCInst1_MC1_n155,
         LED_RoundFunction2_MCInst1_MC1_n154,
         LED_RoundFunction2_MCInst1_MC1_n153,
         LED_RoundFunction2_MCInst1_MC1_n152,
         LED_RoundFunction2_MCInst1_MC1_n151,
         LED_RoundFunction2_MCInst1_MC1_n150,
         LED_RoundFunction2_MCInst1_MC1_n149,
         LED_RoundFunction2_MCInst1_MC1_n148,
         LED_RoundFunction2_MCInst1_MC1_n147,
         LED_RoundFunction2_MCInst1_MC1_n146,
         LED_RoundFunction2_MCInst1_MC1_n145,
         LED_RoundFunction2_MCInst1_MC1_n144,
         LED_RoundFunction2_MCInst1_MC1_n143,
         LED_RoundFunction2_MCInst1_MC1_n142,
         LED_RoundFunction2_MCInst1_MC1_n141,
         LED_RoundFunction2_MCInst1_MC1_n140,
         LED_RoundFunction2_MCInst1_MC1_n139,
         LED_RoundFunction2_MCInst1_MC1_n138,
         LED_RoundFunction2_MCInst1_MC1_n137,
         LED_RoundFunction2_MCInst1_MC1_n136,
         LED_RoundFunction2_MCInst1_MC1_n135,
         LED_RoundFunction2_MCInst1_MC1_n134,
         LED_RoundFunction2_MCInst1_MC1_n133,
         LED_RoundFunction2_MCInst1_MC1_n132,
         LED_RoundFunction2_MCInst1_MC1_n131,
         LED_RoundFunction2_MCInst1_MC1_n130,
         LED_RoundFunction2_MCInst1_MC1_n129,
         LED_RoundFunction2_MCInst1_MC1_n128,
         LED_RoundFunction2_MCInst1_MC1_n127,
         LED_RoundFunction2_MCInst1_MC1_n126,
         LED_RoundFunction2_MCInst1_MC1_n125,
         LED_RoundFunction2_MCInst1_MC1_n124,
         LED_RoundFunction2_MCInst1_MC1_n123,
         LED_RoundFunction2_MCInst1_MC1_n122,
         LED_RoundFunction2_MCInst1_MC1_n121,
         LED_RoundFunction2_MCInst1_MC1_n120,
         LED_RoundFunction2_MCInst1_MC1_n119,
         LED_RoundFunction2_MCInst1_MC1_n118,
         LED_RoundFunction2_MCInst1_MC1_n117,
         LED_RoundFunction2_MCInst1_MC1_n116,
         LED_RoundFunction2_MCInst1_MC1_n115,
         LED_RoundFunction2_MCInst1_MC1_n114,
         LED_RoundFunction2_MCInst1_MC1_n113,
         LED_RoundFunction2_MCInst1_MC1_n112,
         LED_RoundFunction2_MCInst1_MC1_n111,
         LED_RoundFunction2_MCInst1_MC1_n110,
         LED_RoundFunction2_MCInst1_MC1_n109,
         LED_RoundFunction2_MCInst1_MC2_n160,
         LED_RoundFunction2_MCInst1_MC2_n159,
         LED_RoundFunction2_MCInst1_MC2_n158,
         LED_RoundFunction2_MCInst1_MC2_n157,
         LED_RoundFunction2_MCInst1_MC2_n156,
         LED_RoundFunction2_MCInst1_MC2_n155,
         LED_RoundFunction2_MCInst1_MC2_n154,
         LED_RoundFunction2_MCInst1_MC2_n153,
         LED_RoundFunction2_MCInst1_MC2_n152,
         LED_RoundFunction2_MCInst1_MC2_n151,
         LED_RoundFunction2_MCInst1_MC2_n150,
         LED_RoundFunction2_MCInst1_MC2_n149,
         LED_RoundFunction2_MCInst1_MC2_n148,
         LED_RoundFunction2_MCInst1_MC2_n147,
         LED_RoundFunction2_MCInst1_MC2_n146,
         LED_RoundFunction2_MCInst1_MC2_n145,
         LED_RoundFunction2_MCInst1_MC2_n144,
         LED_RoundFunction2_MCInst1_MC2_n143,
         LED_RoundFunction2_MCInst1_MC2_n142,
         LED_RoundFunction2_MCInst1_MC2_n141,
         LED_RoundFunction2_MCInst1_MC2_n140,
         LED_RoundFunction2_MCInst1_MC2_n139,
         LED_RoundFunction2_MCInst1_MC2_n138,
         LED_RoundFunction2_MCInst1_MC2_n137,
         LED_RoundFunction2_MCInst1_MC2_n136,
         LED_RoundFunction2_MCInst1_MC2_n135,
         LED_RoundFunction2_MCInst1_MC2_n134,
         LED_RoundFunction2_MCInst1_MC2_n133,
         LED_RoundFunction2_MCInst1_MC2_n132,
         LED_RoundFunction2_MCInst1_MC2_n131,
         LED_RoundFunction2_MCInst1_MC2_n130,
         LED_RoundFunction2_MCInst1_MC2_n129,
         LED_RoundFunction2_MCInst1_MC2_n128,
         LED_RoundFunction2_MCInst1_MC2_n127,
         LED_RoundFunction2_MCInst1_MC2_n126,
         LED_RoundFunction2_MCInst1_MC2_n125,
         LED_RoundFunction2_MCInst1_MC2_n124,
         LED_RoundFunction2_MCInst1_MC2_n123,
         LED_RoundFunction2_MCInst1_MC2_n122,
         LED_RoundFunction2_MCInst1_MC2_n121,
         LED_RoundFunction2_MCInst1_MC2_n120,
         LED_RoundFunction2_MCInst1_MC2_n119,
         LED_RoundFunction2_MCInst1_MC2_n118,
         LED_RoundFunction2_MCInst1_MC2_n117,
         LED_RoundFunction2_MCInst1_MC2_n116,
         LED_RoundFunction2_MCInst1_MC2_n115,
         LED_RoundFunction2_MCInst1_MC2_n114,
         LED_RoundFunction2_MCInst1_MC2_n113,
         LED_RoundFunction2_MCInst1_MC2_n112,
         LED_RoundFunction2_MCInst1_MC2_n111,
         LED_RoundFunction2_MCInst1_MC2_n110,
         LED_RoundFunction2_MCInst1_MC2_n109,
         LED_RoundFunction2_MCInst1_MC3_n160,
         LED_RoundFunction2_MCInst1_MC3_n159,
         LED_RoundFunction2_MCInst1_MC3_n158,
         LED_RoundFunction2_MCInst1_MC3_n157,
         LED_RoundFunction2_MCInst1_MC3_n156,
         LED_RoundFunction2_MCInst1_MC3_n155,
         LED_RoundFunction2_MCInst1_MC3_n154,
         LED_RoundFunction2_MCInst1_MC3_n153,
         LED_RoundFunction2_MCInst1_MC3_n152,
         LED_RoundFunction2_MCInst1_MC3_n151,
         LED_RoundFunction2_MCInst1_MC3_n150,
         LED_RoundFunction2_MCInst1_MC3_n149,
         LED_RoundFunction2_MCInst1_MC3_n148,
         LED_RoundFunction2_MCInst1_MC3_n147,
         LED_RoundFunction2_MCInst1_MC3_n146,
         LED_RoundFunction2_MCInst1_MC3_n145,
         LED_RoundFunction2_MCInst1_MC3_n144,
         LED_RoundFunction2_MCInst1_MC3_n143,
         LED_RoundFunction2_MCInst1_MC3_n142,
         LED_RoundFunction2_MCInst1_MC3_n141,
         LED_RoundFunction2_MCInst1_MC3_n140,
         LED_RoundFunction2_MCInst1_MC3_n139,
         LED_RoundFunction2_MCInst1_MC3_n138,
         LED_RoundFunction2_MCInst1_MC3_n137,
         LED_RoundFunction2_MCInst1_MC3_n136,
         LED_RoundFunction2_MCInst1_MC3_n135,
         LED_RoundFunction2_MCInst1_MC3_n134,
         LED_RoundFunction2_MCInst1_MC3_n133,
         LED_RoundFunction2_MCInst1_MC3_n132,
         LED_RoundFunction2_MCInst1_MC3_n131,
         LED_RoundFunction2_MCInst1_MC3_n130,
         LED_RoundFunction2_MCInst1_MC3_n129,
         LED_RoundFunction2_MCInst1_MC3_n128,
         LED_RoundFunction2_MCInst1_MC3_n127,
         LED_RoundFunction2_MCInst1_MC3_n126,
         LED_RoundFunction2_MCInst1_MC3_n125,
         LED_RoundFunction2_MCInst1_MC3_n124,
         LED_RoundFunction2_MCInst1_MC3_n123,
         LED_RoundFunction2_MCInst1_MC3_n122,
         LED_RoundFunction2_MCInst1_MC3_n121,
         LED_RoundFunction2_MCInst1_MC3_n120,
         LED_RoundFunction2_MCInst1_MC3_n119,
         LED_RoundFunction2_MCInst1_MC3_n118,
         LED_RoundFunction2_MCInst1_MC3_n117,
         LED_RoundFunction2_MCInst1_MC3_n116,
         LED_RoundFunction2_MCInst1_MC3_n115,
         LED_RoundFunction2_MCInst1_MC3_n114,
         LED_RoundFunction2_MCInst1_MC3_n113,
         LED_RoundFunction2_MCInst1_MC3_n112,
         LED_RoundFunction2_MCInst1_MC3_n111,
         LED_RoundFunction2_MCInst1_MC3_n110,
         LED_RoundFunction2_MCInst1_MC3_n109,
         Inst_SubCell_Multi_Inst_TwoSbox_0_n1,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n36,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n35,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n34,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n33,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n32,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n31,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n30,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n29,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n28,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n27,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n26,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n25,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_n1,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_n1,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_n1,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_n1,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_n1,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_n1,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n79,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n78,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n77,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n76,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n62,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n61,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n60,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n59,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n50,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n49,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n48,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n47,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n46,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n45,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n44,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n43,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n42,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n41,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n40,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n39,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N2,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_0__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_3__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_6__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_9__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_12__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_15__CF_Inst_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n20,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n19,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n18,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n17,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n16,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n15,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n14,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n13,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_n2,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_N1,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_N0,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n12,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n11,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n10,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_n6,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_n5,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n9,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n8,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n7,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression3_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression1_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression2_n3,
         Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression3_n3,
         LED128_Controller_Inst_n48, LED128_Controller_Inst_n38,
         LED128_Controller_Inst_n37, LED128_Controller_Inst_n36,
         LED128_Controller_Inst_n35, LED128_Controller_Inst_n34,
         LED128_Controller_Inst_n33, LED128_Controller_Inst_n32,
         LED128_Controller_Inst_n31, LED128_Controller_Inst_n30,
         LED128_Controller_Inst_n29, LED128_Controller_Inst_n28,
         LED128_Controller_Inst_n27, LED128_Controller_Inst_n26,
         LED128_Controller_Inst_n25, LED128_Controller_Inst_n24,
         LED128_Controller_Inst_n23, LED128_Controller_Inst_n22,
         LED128_Controller_Inst_n21, LED128_Controller_Inst_n20,
         LED128_Controller_Inst_n18, LED128_Controller_Inst_n17,
         LED128_Controller_Inst_n16, LED128_Controller_Inst_n14,
         LED128_Controller_Inst_n13, LED128_Controller_Inst_n11,
         LED128_Controller_Inst_n10, LED128_Controller_Inst_n8,
         LED128_Controller_Inst_n47, LED128_Controller_Inst_n40,
         LED128_Controller_Inst_n39, LED128_Controller_Inst_n19,
         LED128_Controller_Inst_n2, LED128_Controller_Inst_n1,
         LED128_Controller_Inst_n46, LED128_Controller_Inst_n45,
         LED128_Controller_Inst_n44, LED128_Controller_Inst_n43,
         LED128_Controller_Inst_n42, LED128_Controller_Inst_n41,
         LED128_Controller_Inst_n15, LED128_Controller_Inst_n12,
         LED128_Controller_Inst_n9, LED128_Controller_Inst_n7,
         LED128_Controller_Inst_n6, LED128_Controller_Inst_n3;
  wire   [5:0] FSM;
  wire   [63:0] SubCellOutput0;
  wire   [62:2] SubCellInput0;
  wire   [63:0] SubCellOutput1;
  wire   [62:2] SubCellInput1;
  wire   [63:0] SubCellOutput2;
  wire   [62:2] SubCellInput2;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_0_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_0_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_1_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_1_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_2_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_2_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_3_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_3_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_4_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_4_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_5_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_5_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_6_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_6_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_7_rs1;
  wire   [7:0] Inst_SubCell_Multi_Inst_TwoSbox_7_rs2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2;
  wire   [3:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg;
  wire   [26:0] Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out;

  AOI22_X1 LED_RoundFunction0_U412 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n562), .B1(LED_RoundFunction0_n561), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U411 ( .A1(rst), .A2(Plaintext0[0]), .B1(
        LED_RoundFunction0_Feedback_0_), .B2(LED_RoundFunction0_n290), .ZN(
        LED_RoundFunction0_n561) );
  INV_X1 LED_RoundFunction0_U410 ( .A(Ciphertext0[0]), .ZN(
        LED_RoundFunction0_n562) );
  AOI22_X1 LED_RoundFunction0_U409 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n560), .B1(LED_RoundFunction0_n559), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U408 ( .A1(rst), .A2(Plaintext0[1]), .B1(
        LED_RoundFunction0_Feedback_1_), .B2(LED_RoundFunction0_n294), .ZN(
        LED_RoundFunction0_n559) );
  INV_X1 LED_RoundFunction0_U407 ( .A(Ciphertext0[1]), .ZN(
        LED_RoundFunction0_n560) );
  AOI22_X1 LED_RoundFunction0_U406 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n558), .B1(LED_RoundFunction0_n557), .B2(
        LED_RoundFunction0_n287), .ZN(SubCellInput0[2]) );
  AOI22_X1 LED_RoundFunction0_U405 ( .A1(rst), .A2(Plaintext0[2]), .B1(
        LED_RoundFunction0_Feedback_2_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n557) );
  INV_X1 LED_RoundFunction0_U404 ( .A(Ciphertext0[2]), .ZN(
        LED_RoundFunction0_n558) );
  AOI22_X1 LED_RoundFunction0_U403 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n556), .B1(LED_RoundFunction0_n555), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U402 ( .A1(rst), .A2(Plaintext0[3]), .B1(
        LED_RoundFunction0_Feedback_3_), .B2(LED_RoundFunction0_n294), .ZN(
        LED_RoundFunction0_n555) );
  INV_X1 LED_RoundFunction0_U401 ( .A(Ciphertext0[3]), .ZN(
        LED_RoundFunction0_n556) );
  AOI22_X1 LED_RoundFunction0_U400 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n554), .B1(LED_RoundFunction0_n553), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U399 ( .A1(rst), .A2(Plaintext0[4]), .B1(
        LED_RoundFunction0_Feedback_4_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n553) );
  INV_X1 LED_RoundFunction0_U398 ( .A(Ciphertext0[4]), .ZN(
        LED_RoundFunction0_n554) );
  AOI22_X1 LED_RoundFunction0_U397 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n552), .B1(LED_RoundFunction0_n551), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U396 ( .A1(rst), .A2(Plaintext0[5]), .B1(
        LED_RoundFunction0_Feedback_5_), .B2(LED_RoundFunction0_n294), .ZN(
        LED_RoundFunction0_n551) );
  INV_X1 LED_RoundFunction0_U395 ( .A(Ciphertext0[5]), .ZN(
        LED_RoundFunction0_n552) );
  AOI22_X1 LED_RoundFunction0_U394 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n550), .B1(LED_RoundFunction0_n549), .B2(
        LED_RoundFunction0_n286), .ZN(SubCellInput0[6]) );
  AOI22_X1 LED_RoundFunction0_U393 ( .A1(rst), .A2(Plaintext0[6]), .B1(
        LED_RoundFunction0_Feedback_6_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n549) );
  INV_X1 LED_RoundFunction0_U392 ( .A(Ciphertext0[6]), .ZN(
        LED_RoundFunction0_n550) );
  AOI22_X1 LED_RoundFunction0_U391 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n548), .B1(LED_RoundFunction0_n547), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U390 ( .A1(rst), .A2(Plaintext0[7]), .B1(
        LED_RoundFunction0_Feedback_7_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n547) );
  INV_X1 LED_RoundFunction0_U389 ( .A(Ciphertext0[7]), .ZN(
        LED_RoundFunction0_n548) );
  AOI22_X1 LED_RoundFunction0_U388 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n546), .B1(LED_RoundFunction0_n545), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U387 ( .A1(rst), .A2(Plaintext0[11]), .B1(
        LED_RoundFunction0_Feedback_11_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n545) );
  INV_X1 LED_RoundFunction0_U386 ( .A(Ciphertext0[11]), .ZN(
        LED_RoundFunction0_n546) );
  AOI22_X1 LED_RoundFunction0_U385 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n544), .B1(LED_RoundFunction0_n543), .B2(
        LED_RoundFunction0_n287), .ZN(SubCellInput0[14]) );
  AOI22_X1 LED_RoundFunction0_U384 ( .A1(rst), .A2(Plaintext0[14]), .B1(
        LED_RoundFunction0_Feedback_14_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n543) );
  INV_X1 LED_RoundFunction0_U383 ( .A(Ciphertext0[14]), .ZN(
        LED_RoundFunction0_n544) );
  AOI22_X1 LED_RoundFunction0_U382 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n542), .B1(LED_RoundFunction0_n541), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U381 ( .A1(rst), .A2(Plaintext0[15]), .B1(
        LED_RoundFunction0_Feedback_15_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n541) );
  INV_X1 LED_RoundFunction0_U380 ( .A(Ciphertext0[15]), .ZN(
        LED_RoundFunction0_n542) );
  AOI22_X1 LED_RoundFunction0_U379 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n540), .B1(LED_RoundFunction0_n539), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U378 ( .A1(rst), .A2(Plaintext0[16]), .B1(
        LED_RoundFunction0_Feedback_16_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n539) );
  INV_X1 LED_RoundFunction0_U377 ( .A(Ciphertext0[16]), .ZN(
        LED_RoundFunction0_n540) );
  AOI22_X1 LED_RoundFunction0_U376 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n538), .B1(LED_RoundFunction0_n537), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U375 ( .A1(rst), .A2(Plaintext0[17]), .B1(
        LED_RoundFunction0_Feedback_17_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n537) );
  INV_X1 LED_RoundFunction0_U374 ( .A(Ciphertext0[17]), .ZN(
        LED_RoundFunction0_n538) );
  AOI22_X1 LED_RoundFunction0_U373 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n536), .B1(LED_RoundFunction0_n535), .B2(
        LED_RoundFunction0_n286), .ZN(SubCellInput0[18]) );
  AOI22_X1 LED_RoundFunction0_U372 ( .A1(rst), .A2(Plaintext0[18]), .B1(
        LED_RoundFunction0_Feedback_18_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n535) );
  INV_X1 LED_RoundFunction0_U371 ( .A(Ciphertext0[18]), .ZN(
        LED_RoundFunction0_n536) );
  AOI22_X1 LED_RoundFunction0_U370 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n534), .B1(LED_RoundFunction0_n533), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U369 ( .A1(rst), .A2(Plaintext0[19]), .B1(
        LED_RoundFunction0_Feedback_19_), .B2(LED_RoundFunction0_n294), .ZN(
        LED_RoundFunction0_n533) );
  INV_X1 LED_RoundFunction0_U368 ( .A(Ciphertext0[19]), .ZN(
        LED_RoundFunction0_n534) );
  AOI22_X1 LED_RoundFunction0_U367 ( .A1(LED_RoundFunction0_n283), .A2(
        LED_RoundFunction0_n532), .B1(LED_RoundFunction0_n531), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U366 ( .A1(rst), .A2(Plaintext0[20]), .B1(
        LED_RoundFunction0_Feedback_20_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n531) );
  INV_X1 LED_RoundFunction0_U365 ( .A(Ciphertext0[20]), .ZN(
        LED_RoundFunction0_n532) );
  AOI22_X1 LED_RoundFunction0_U364 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n530), .B1(LED_RoundFunction0_n529), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U363 ( .A1(rst), .A2(Plaintext0[21]), .B1(
        LED_RoundFunction0_Feedback_21_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n529) );
  INV_X1 LED_RoundFunction0_U362 ( .A(Ciphertext0[21]), .ZN(
        LED_RoundFunction0_n530) );
  AOI22_X1 LED_RoundFunction0_U361 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n528), .B1(LED_RoundFunction0_n527), .B2(
        LED_RoundFunction0_n287), .ZN(SubCellInput0[22]) );
  AOI22_X1 LED_RoundFunction0_U360 ( .A1(rst), .A2(Plaintext0[22]), .B1(
        LED_RoundFunction0_Feedback_22_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n527) );
  INV_X1 LED_RoundFunction0_U359 ( .A(Ciphertext0[22]), .ZN(
        LED_RoundFunction0_n528) );
  AOI22_X1 LED_RoundFunction0_U358 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n526), .B1(LED_RoundFunction0_n525), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U357 ( .A1(rst), .A2(Plaintext0[23]), .B1(
        LED_RoundFunction0_Feedback_23_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n525) );
  INV_X1 LED_RoundFunction0_U356 ( .A(Ciphertext0[23]), .ZN(
        LED_RoundFunction0_n526) );
  AOI22_X1 LED_RoundFunction0_U355 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n524), .B1(LED_RoundFunction0_n523), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U354 ( .A1(rst), .A2(Plaintext0[27]), .B1(
        LED_RoundFunction0_Feedback_27_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n523) );
  INV_X1 LED_RoundFunction0_U353 ( .A(Ciphertext0[27]), .ZN(
        LED_RoundFunction0_n524) );
  AOI22_X1 LED_RoundFunction0_U352 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n522), .B1(LED_RoundFunction0_n521), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U351 ( .A1(rst), .A2(Plaintext0[28]), .B1(
        LED_RoundFunction0_Feedback_28_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n521) );
  INV_X1 LED_RoundFunction0_U350 ( .A(Ciphertext0[28]), .ZN(
        LED_RoundFunction0_n522) );
  AOI22_X1 LED_RoundFunction0_U349 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n520), .B1(LED_RoundFunction0_n519), .B2(
        LED_RoundFunction0_n286), .ZN(SubCellInput0[30]) );
  AOI22_X1 LED_RoundFunction0_U348 ( .A1(rst), .A2(Plaintext0[30]), .B1(
        LED_RoundFunction0_Feedback_30_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n519) );
  INV_X1 LED_RoundFunction0_U347 ( .A(Ciphertext0[30]), .ZN(
        LED_RoundFunction0_n520) );
  AOI22_X1 LED_RoundFunction0_U346 ( .A1(LED_RoundFunction0_n282), .A2(
        LED_RoundFunction0_n518), .B1(LED_RoundFunction0_n517), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U345 ( .A1(rst), .A2(Plaintext0[31]), .B1(
        LED_RoundFunction0_Feedback_31_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n517) );
  INV_X1 LED_RoundFunction0_U344 ( .A(Ciphertext0[31]), .ZN(
        LED_RoundFunction0_n518) );
  AOI22_X1 LED_RoundFunction0_U343 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n516), .B1(LED_RoundFunction0_n515), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U342 ( .A1(rst), .A2(Plaintext0[32]), .B1(
        LED_RoundFunction0_Feedback_32_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n515) );
  INV_X1 LED_RoundFunction0_U341 ( .A(Ciphertext0[32]), .ZN(
        LED_RoundFunction0_n516) );
  AOI22_X1 LED_RoundFunction0_U340 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n514), .B1(LED_RoundFunction0_n513), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U339 ( .A1(rst), .A2(Plaintext0[33]), .B1(
        LED_RoundFunction0_Feedback_33_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n513) );
  INV_X1 LED_RoundFunction0_U338 ( .A(Ciphertext0[33]), .ZN(
        LED_RoundFunction0_n514) );
  AOI22_X1 LED_RoundFunction0_U337 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n512), .B1(LED_RoundFunction0_n511), .B2(
        LED_RoundFunction0_n287), .ZN(SubCellInput0[34]) );
  AOI22_X1 LED_RoundFunction0_U336 ( .A1(rst), .A2(Plaintext0[34]), .B1(
        LED_RoundFunction0_Feedback_34_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n511) );
  INV_X1 LED_RoundFunction0_U335 ( .A(Ciphertext0[34]), .ZN(
        LED_RoundFunction0_n512) );
  AOI22_X1 LED_RoundFunction0_U334 ( .A1(LED_RoundFunction0_n283), .A2(
        LED_RoundFunction0_n510), .B1(LED_RoundFunction0_n509), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U333 ( .A1(rst), .A2(Plaintext0[35]), .B1(
        LED_RoundFunction0_Feedback_35_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n509) );
  INV_X1 LED_RoundFunction0_U332 ( .A(Ciphertext0[35]), .ZN(
        LED_RoundFunction0_n510) );
  AOI22_X1 LED_RoundFunction0_U331 ( .A1(LED_RoundFunction0_n282), .A2(
        LED_RoundFunction0_n508), .B1(LED_RoundFunction0_n507), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U330 ( .A1(rst), .A2(Plaintext0[36]), .B1(
        LED_RoundFunction0_Feedback_36_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n507) );
  INV_X1 LED_RoundFunction0_U329 ( .A(Ciphertext0[36]), .ZN(
        LED_RoundFunction0_n508) );
  AOI22_X1 LED_RoundFunction0_U328 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n506), .B1(LED_RoundFunction0_n505), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U327 ( .A1(rst), .A2(Plaintext0[37]), .B1(
        LED_RoundFunction0_Feedback_37_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n505) );
  INV_X1 LED_RoundFunction0_U326 ( .A(Ciphertext0[37]), .ZN(
        LED_RoundFunction0_n506) );
  AOI22_X1 LED_RoundFunction0_U325 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n504), .B1(LED_RoundFunction0_n503), .B2(
        LED_RoundFunction0_n287), .ZN(SubCellInput0[38]) );
  AOI22_X1 LED_RoundFunction0_U324 ( .A1(rst), .A2(Plaintext0[38]), .B1(
        LED_RoundFunction0_Feedback_38_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n503) );
  INV_X1 LED_RoundFunction0_U323 ( .A(Ciphertext0[38]), .ZN(
        LED_RoundFunction0_n504) );
  AOI22_X1 LED_RoundFunction0_U322 ( .A1(LED_RoundFunction0_n282), .A2(
        LED_RoundFunction0_n502), .B1(LED_RoundFunction0_n501), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U321 ( .A1(rst), .A2(Plaintext0[39]), .B1(
        LED_RoundFunction0_Feedback_39_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n501) );
  INV_X1 LED_RoundFunction0_U320 ( .A(Ciphertext0[39]), .ZN(
        LED_RoundFunction0_n502) );
  AOI22_X1 LED_RoundFunction0_U319 ( .A1(LED_RoundFunction0_n283), .A2(
        LED_RoundFunction0_n500), .B1(LED_RoundFunction0_n499), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U318 ( .A1(rst), .A2(Plaintext0[43]), .B1(
        LED_RoundFunction0_Feedback_43_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n499) );
  INV_X1 LED_RoundFunction0_U317 ( .A(Ciphertext0[43]), .ZN(
        LED_RoundFunction0_n500) );
  AOI22_X1 LED_RoundFunction0_U316 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n498), .B1(LED_RoundFunction0_n497), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U315 ( .A1(rst), .A2(Plaintext0[45]), .B1(
        LED_RoundFunction0_Feedback_45_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n497) );
  INV_X1 LED_RoundFunction0_U314 ( .A(Ciphertext0[45]), .ZN(
        LED_RoundFunction0_n498) );
  AOI22_X1 LED_RoundFunction0_U313 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n496), .B1(LED_RoundFunction0_n495), .B2(
        LED_RoundFunction0_n287), .ZN(SubCellInput0[46]) );
  AOI22_X1 LED_RoundFunction0_U312 ( .A1(rst), .A2(Plaintext0[46]), .B1(
        LED_RoundFunction0_Feedback_46_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n495) );
  INV_X1 LED_RoundFunction0_U311 ( .A(Ciphertext0[46]), .ZN(
        LED_RoundFunction0_n496) );
  AOI22_X1 LED_RoundFunction0_U310 ( .A1(LED_RoundFunction0_n283), .A2(
        LED_RoundFunction0_n494), .B1(LED_RoundFunction0_n493), .B2(
        LED_RoundFunction0_n287), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U309 ( .A1(rst), .A2(Plaintext0[48]), .B1(
        LED_RoundFunction0_Feedback_48_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n493) );
  INV_X1 LED_RoundFunction0_U308 ( .A(Ciphertext0[48]), .ZN(
        LED_RoundFunction0_n494) );
  AOI22_X1 LED_RoundFunction0_U307 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n492), .B1(LED_RoundFunction0_n491), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U306 ( .A1(rst), .A2(Plaintext0[49]), .B1(
        LED_RoundFunction0_Feedback_49_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n491) );
  INV_X1 LED_RoundFunction0_U305 ( .A(Ciphertext0[49]), .ZN(
        LED_RoundFunction0_n492) );
  AOI22_X1 LED_RoundFunction0_U304 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n490), .B1(LED_RoundFunction0_n489), .B2(
        LED_RoundFunction0_n286), .ZN(SubCellInput0[50]) );
  AOI22_X1 LED_RoundFunction0_U303 ( .A1(rst), .A2(Plaintext0[50]), .B1(
        LED_RoundFunction0_Feedback_50_), .B2(LED_RoundFunction0_n288), .ZN(
        LED_RoundFunction0_n489) );
  INV_X1 LED_RoundFunction0_U302 ( .A(Ciphertext0[50]), .ZN(
        LED_RoundFunction0_n490) );
  AOI22_X1 LED_RoundFunction0_U301 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n488), .B1(LED_RoundFunction0_n487), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U300 ( .A1(rst), .A2(Plaintext0[51]), .B1(
        LED_RoundFunction0_Feedback_51_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n487) );
  INV_X1 LED_RoundFunction0_U299 ( .A(Ciphertext0[51]), .ZN(
        LED_RoundFunction0_n488) );
  AOI22_X1 LED_RoundFunction0_U298 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n486), .B1(LED_RoundFunction0_n485), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U297 ( .A1(rst), .A2(Plaintext0[52]), .B1(
        LED_RoundFunction0_Feedback_52_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n485) );
  INV_X1 LED_RoundFunction0_U296 ( .A(Ciphertext0[52]), .ZN(
        LED_RoundFunction0_n486) );
  AOI22_X1 LED_RoundFunction0_U295 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n484), .B1(LED_RoundFunction0_n483), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U294 ( .A1(rst), .A2(Plaintext0[53]), .B1(
        LED_RoundFunction0_Feedback_53_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n483) );
  INV_X1 LED_RoundFunction0_U293 ( .A(Ciphertext0[53]), .ZN(
        LED_RoundFunction0_n484) );
  AOI22_X1 LED_RoundFunction0_U292 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n482), .B1(LED_RoundFunction0_n481), .B2(
        LED_RoundFunction0_n286), .ZN(SubCellInput0[54]) );
  AOI22_X1 LED_RoundFunction0_U291 ( .A1(rst), .A2(Plaintext0[54]), .B1(
        LED_RoundFunction0_Feedback_54_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n481) );
  INV_X1 LED_RoundFunction0_U290 ( .A(Ciphertext0[54]), .ZN(
        LED_RoundFunction0_n482) );
  AOI22_X1 LED_RoundFunction0_U289 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n480), .B1(LED_RoundFunction0_n479), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U288 ( .A1(rst), .A2(Plaintext0[55]), .B1(
        LED_RoundFunction0_Feedback_55_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n479) );
  INV_X1 LED_RoundFunction0_U287 ( .A(Ciphertext0[55]), .ZN(
        LED_RoundFunction0_n480) );
  AOI22_X1 LED_RoundFunction0_U286 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n478), .B1(LED_RoundFunction0_n477), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[1]) );
  AOI22_X1 LED_RoundFunction0_U285 ( .A1(rst), .A2(Plaintext0[59]), .B1(
        LED_RoundFunction0_Feedback_59_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n477) );
  INV_X1 LED_RoundFunction0_U284 ( .A(Ciphertext0[59]), .ZN(
        LED_RoundFunction0_n478) );
  AOI22_X1 LED_RoundFunction0_U283 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n476), .B1(LED_RoundFunction0_n475), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[0]) );
  AOI22_X1 LED_RoundFunction0_U282 ( .A1(rst), .A2(Plaintext0[60]), .B1(
        LED_RoundFunction0_Feedback_60_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n475) );
  INV_X1 LED_RoundFunction0_U281 ( .A(Ciphertext0[60]), .ZN(
        LED_RoundFunction0_n476) );
  AOI22_X1 LED_RoundFunction0_U280 ( .A1(LED_RoundFunction0_n284), .A2(
        LED_RoundFunction0_n474), .B1(LED_RoundFunction0_n473), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[2]) );
  AOI22_X1 LED_RoundFunction0_U279 ( .A1(rst), .A2(Plaintext0[61]), .B1(
        LED_RoundFunction0_Feedback_61_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n473) );
  INV_X1 LED_RoundFunction0_U278 ( .A(Ciphertext0[61]), .ZN(
        LED_RoundFunction0_n474) );
  AOI22_X1 LED_RoundFunction0_U277 ( .A1(LED_RoundFunction0_n281), .A2(
        LED_RoundFunction0_n472), .B1(LED_RoundFunction0_n471), .B2(
        LED_RoundFunction0_n286), .ZN(SubCellInput0[62]) );
  AOI22_X1 LED_RoundFunction0_U276 ( .A1(rst), .A2(Plaintext0[62]), .B1(
        LED_RoundFunction0_Feedback_62_), .B2(LED_RoundFunction0_n289), .ZN(
        LED_RoundFunction0_n471) );
  INV_X1 LED_RoundFunction0_U275 ( .A(Ciphertext0[62]), .ZN(
        LED_RoundFunction0_n472) );
  XOR2_X1 LED_RoundFunction0_U274 ( .A(FSM[1]), .B(LED_RoundFunction0_n470), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[2]) );
  AOI21_X1 LED_RoundFunction0_U273 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n469), .A(LED_RoundFunction0_n468), .ZN(
        LED_RoundFunction0_n470) );
  AOI221_X1 LED_RoundFunction0_U272 ( .B1(Plaintext0[9]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_9_), .C2(LED_RoundFunction0_n294), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n468) );
  INV_X1 LED_RoundFunction0_U271 ( .A(Ciphertext0[9]), .ZN(
        LED_RoundFunction0_n469) );
  XOR2_X1 LED_RoundFunction0_U270 ( .A(FSM[0]), .B(LED_RoundFunction0_n467), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[0]) );
  AOI21_X1 LED_RoundFunction0_U269 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n466), .A(LED_RoundFunction0_n465), .ZN(
        LED_RoundFunction0_n467) );
  AOI221_X1 LED_RoundFunction0_U268 ( .B1(Plaintext0[8]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_8_), .C2(LED_RoundFunction0_n292), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n465) );
  INV_X1 LED_RoundFunction0_U267 ( .A(Ciphertext0[8]), .ZN(
        LED_RoundFunction0_n466) );
  AOI22_X1 LED_RoundFunction0_U266 ( .A1(LED_RoundFunction0_n281), .A2(
        Ciphertext0[63]), .B1(LED_RoundFunction0_n464), .B2(
        LED_RoundFunction0_n286), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[1]) );
  INV_X1 LED_RoundFunction0_U265 ( .A(LED_RoundFunction0_n463), .ZN(
        LED_RoundFunction0_n464) );
  OAI22_X1 LED_RoundFunction0_U264 ( .A1(LED_RoundFunction0_n291), .A2(
        Plaintext0[63]), .B1(LED_RoundFunction0_Feedback_63_), .B2(rst), .ZN(
        LED_RoundFunction0_n463) );
  XOR2_X1 LED_RoundFunction0_U263 ( .A(FSM[5]), .B(LED_RoundFunction0_n462), 
        .Z(SubCellInput0[58]) );
  AOI21_X1 LED_RoundFunction0_U262 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n461), .A(LED_RoundFunction0_n460), .ZN(
        LED_RoundFunction0_n462) );
  AOI221_X1 LED_RoundFunction0_U261 ( .B1(Plaintext0[58]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_58_), .C2(LED_RoundFunction0_n291), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n460) );
  INV_X1 LED_RoundFunction0_U260 ( .A(Ciphertext0[58]), .ZN(
        LED_RoundFunction0_n461) );
  XOR2_X1 LED_RoundFunction0_U259 ( .A(FSM[4]), .B(LED_RoundFunction0_n459), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[2]) );
  AOI21_X1 LED_RoundFunction0_U258 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n458), .A(LED_RoundFunction0_n457), .ZN(
        LED_RoundFunction0_n459) );
  AOI221_X1 LED_RoundFunction0_U257 ( .B1(Plaintext0[57]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_57_), .C2(LED_RoundFunction0_n292), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n457) );
  INV_X1 LED_RoundFunction0_U256 ( .A(Ciphertext0[57]), .ZN(
        LED_RoundFunction0_n458) );
  XOR2_X1 LED_RoundFunction0_U255 ( .A(FSM[3]), .B(LED_RoundFunction0_n456), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[0]) );
  AOI21_X1 LED_RoundFunction0_U254 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n455), .A(LED_RoundFunction0_n454), .ZN(
        LED_RoundFunction0_n456) );
  AOI221_X1 LED_RoundFunction0_U253 ( .B1(Plaintext0[56]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_56_), .C2(LED_RoundFunction0_n294), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n454) );
  INV_X1 LED_RoundFunction0_U252 ( .A(Ciphertext0[56]), .ZN(
        LED_RoundFunction0_n455) );
  AOI22_X1 LED_RoundFunction0_U251 ( .A1(LED_RoundFunction0_n282), .A2(
        Ciphertext0[47]), .B1(LED_RoundFunction0_n453), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[1]) );
  INV_X1 LED_RoundFunction0_U250 ( .A(LED_RoundFunction0_n452), .ZN(
        LED_RoundFunction0_n453) );
  OAI22_X1 LED_RoundFunction0_U249 ( .A1(LED_RoundFunction0_n294), .A2(
        Plaintext0[47]), .B1(LED_RoundFunction0_Feedback_47_), .B2(rst), .ZN(
        LED_RoundFunction0_n452) );
  AOI22_X1 LED_RoundFunction0_U248 ( .A1(LED_RoundFunction0_n282), .A2(
        Ciphertext0[44]), .B1(LED_RoundFunction0_n451), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[0]) );
  INV_X1 LED_RoundFunction0_U247 ( .A(LED_RoundFunction0_n450), .ZN(
        LED_RoundFunction0_n451) );
  OAI22_X1 LED_RoundFunction0_U246 ( .A1(LED_RoundFunction0_n294), .A2(
        Plaintext0[44]), .B1(LED_RoundFunction0_Feedback_44_), .B2(rst), .ZN(
        LED_RoundFunction0_n450) );
  XOR2_X1 LED_RoundFunction0_U245 ( .A(FSM[2]), .B(LED_RoundFunction0_n449), 
        .Z(SubCellInput0[42]) );
  AOI21_X1 LED_RoundFunction0_U244 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n448), .A(LED_RoundFunction0_n447), .ZN(
        LED_RoundFunction0_n449) );
  AOI221_X1 LED_RoundFunction0_U243 ( .B1(Plaintext0[42]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_42_), .C2(LED_RoundFunction0_n294), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n447) );
  INV_X1 LED_RoundFunction0_U242 ( .A(Ciphertext0[42]), .ZN(
        LED_RoundFunction0_n448) );
  XOR2_X1 LED_RoundFunction0_U241 ( .A(FSM[1]), .B(LED_RoundFunction0_n446), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[2]) );
  AOI21_X1 LED_RoundFunction0_U240 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n445), .A(LED_RoundFunction0_n444), .ZN(
        LED_RoundFunction0_n446) );
  AOI221_X1 LED_RoundFunction0_U239 ( .B1(Plaintext0[41]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_41_), .C2(LED_RoundFunction0_n291), .A(
        LED_RoundFunction0_n283), .ZN(LED_RoundFunction0_n444) );
  INV_X1 LED_RoundFunction0_U238 ( .A(Ciphertext0[41]), .ZN(
        LED_RoundFunction0_n445) );
  XOR2_X1 LED_RoundFunction0_U237 ( .A(FSM[0]), .B(LED_RoundFunction0_n443), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[0]) );
  AOI21_X1 LED_RoundFunction0_U236 ( .B1(LED_RoundFunction0_n283), .B2(
        LED_RoundFunction0_n442), .A(LED_RoundFunction0_n441), .ZN(
        LED_RoundFunction0_n443) );
  AOI221_X1 LED_RoundFunction0_U235 ( .B1(Plaintext0[40]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_40_), .C2(LED_RoundFunction0_n294), .A(
        LED_RoundFunction0_n283), .ZN(LED_RoundFunction0_n441) );
  INV_X1 LED_RoundFunction0_U234 ( .A(Ciphertext0[40]), .ZN(
        LED_RoundFunction0_n442) );
  AOI22_X1 LED_RoundFunction0_U233 ( .A1(LED_RoundFunction0_n282), .A2(
        Ciphertext0[29]), .B1(LED_RoundFunction0_n440), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[2]) );
  INV_X1 LED_RoundFunction0_U232 ( .A(LED_RoundFunction0_n439), .ZN(
        LED_RoundFunction0_n440) );
  OAI22_X1 LED_RoundFunction0_U231 ( .A1(LED_RoundFunction0_n291), .A2(
        Plaintext0[29]), .B1(LED_RoundFunction0_Feedback_29_), .B2(rst), .ZN(
        LED_RoundFunction0_n439) );
  XOR2_X1 LED_RoundFunction0_U230 ( .A(FSM[5]), .B(LED_RoundFunction0_n438), 
        .Z(SubCellInput0[26]) );
  AOI21_X1 LED_RoundFunction0_U229 ( .B1(LED_RoundFunction0_n284), .B2(
        LED_RoundFunction0_n437), .A(LED_RoundFunction0_n436), .ZN(
        LED_RoundFunction0_n438) );
  AOI221_X1 LED_RoundFunction0_U228 ( .B1(Plaintext0[26]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_26_), .C2(LED_RoundFunction0_n294), .A(
        LED_RoundFunction0_n283), .ZN(LED_RoundFunction0_n436) );
  INV_X1 LED_RoundFunction0_U227 ( .A(Ciphertext0[26]), .ZN(
        LED_RoundFunction0_n437) );
  XOR2_X1 LED_RoundFunction0_U226 ( .A(FSM[4]), .B(LED_RoundFunction0_n435), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[2]) );
  AOI21_X1 LED_RoundFunction0_U225 ( .B1(LED_RoundFunction0_n284), .B2(
        LED_RoundFunction0_n434), .A(LED_RoundFunction0_n433), .ZN(
        LED_RoundFunction0_n435) );
  AOI221_X1 LED_RoundFunction0_U224 ( .B1(Plaintext0[25]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_25_), .C2(LED_RoundFunction0_n294), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n433) );
  INV_X1 LED_RoundFunction0_U223 ( .A(Ciphertext0[25]), .ZN(
        LED_RoundFunction0_n434) );
  XOR2_X1 LED_RoundFunction0_U222 ( .A(FSM[3]), .B(LED_RoundFunction0_n432), 
        .Z(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[0]) );
  AOI21_X1 LED_RoundFunction0_U221 ( .B1(LED_RoundFunction0_n284), .B2(
        LED_RoundFunction0_n431), .A(LED_RoundFunction0_n430), .ZN(
        LED_RoundFunction0_n432) );
  AOI221_X1 LED_RoundFunction0_U220 ( .B1(Plaintext0[24]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_24_), .C2(LED_RoundFunction0_n292), .A(
        LED_RoundFunction0_n283), .ZN(LED_RoundFunction0_n430) );
  INV_X1 LED_RoundFunction0_U219 ( .A(Ciphertext0[24]), .ZN(
        LED_RoundFunction0_n431) );
  AOI22_X1 LED_RoundFunction0_U218 ( .A1(LED_RoundFunction0_n282), .A2(
        Ciphertext0[13]), .B1(LED_RoundFunction0_n429), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[2]) );
  INV_X1 LED_RoundFunction0_U217 ( .A(LED_RoundFunction0_n428), .ZN(
        LED_RoundFunction0_n429) );
  OAI22_X1 LED_RoundFunction0_U216 ( .A1(LED_RoundFunction0_n294), .A2(
        Plaintext0[13]), .B1(LED_RoundFunction0_Feedback_13_), .B2(rst), .ZN(
        LED_RoundFunction0_n428) );
  AOI22_X1 LED_RoundFunction0_U215 ( .A1(LED_RoundFunction0_n282), .A2(
        Ciphertext0[12]), .B1(LED_RoundFunction0_n427), .B2(
        LED_RoundFunction0_n285), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[0]) );
  INV_X1 LED_RoundFunction0_U214 ( .A(LED_RoundFunction0_n426), .ZN(
        LED_RoundFunction0_n427) );
  OAI22_X1 LED_RoundFunction0_U213 ( .A1(LED_RoundFunction0_n291), .A2(
        Plaintext0[12]), .B1(LED_RoundFunction0_Feedback_12_), .B2(rst), .ZN(
        LED_RoundFunction0_n426) );
  XOR2_X1 LED_RoundFunction0_U212 ( .A(FSM[2]), .B(LED_RoundFunction0_n425), 
        .Z(SubCellInput0[10]) );
  AOI21_X1 LED_RoundFunction0_U211 ( .B1(LED_RoundFunction0_n284), .B2(
        LED_RoundFunction0_n424), .A(LED_RoundFunction0_n423), .ZN(
        LED_RoundFunction0_n425) );
  AOI221_X1 LED_RoundFunction0_U210 ( .B1(Plaintext0[10]), .B2(rst), .C1(
        LED_RoundFunction0_Feedback_10_), .C2(LED_RoundFunction0_n291), .A(
        LED_RoundFunction0_n282), .ZN(LED_RoundFunction0_n423) );
  INV_X1 LED_RoundFunction0_U209 ( .A(Ciphertext0[10]), .ZN(
        LED_RoundFunction0_n424) );
  AOI22_X1 LED_RoundFunction0_U208 ( .A1(rst), .A2(LED_RoundFunction0_n422), 
        .B1(LED_RoundFunction0_n421), .B2(LED_RoundFunction0_n289), .ZN(
        Ciphertext0[9]) );
  XNOR2_X1 LED_RoundFunction0_U207 ( .A(LED_RoundFunction0_Feedback_9_), .B(
        Key0[73]), .ZN(LED_RoundFunction0_n421) );
  XNOR2_X1 LED_RoundFunction0_U206 ( .A(Plaintext0[9]), .B(Key0[9]), .ZN(
        LED_RoundFunction0_n422) );
  AOI22_X1 LED_RoundFunction0_U205 ( .A1(rst), .A2(LED_RoundFunction0_n420), 
        .B1(LED_RoundFunction0_n419), .B2(LED_RoundFunction0_n289), .ZN(
        Ciphertext0[8]) );
  XNOR2_X1 LED_RoundFunction0_U204 ( .A(LED_RoundFunction0_Feedback_8_), .B(
        Key0[72]), .ZN(LED_RoundFunction0_n419) );
  XNOR2_X1 LED_RoundFunction0_U203 ( .A(Plaintext0[8]), .B(Key0[8]), .ZN(
        LED_RoundFunction0_n420) );
  AOI22_X1 LED_RoundFunction0_U202 ( .A1(rst), .A2(LED_RoundFunction0_n418), 
        .B1(LED_RoundFunction0_n417), .B2(LED_RoundFunction0_n289), .ZN(
        Ciphertext0[7]) );
  XNOR2_X1 LED_RoundFunction0_U201 ( .A(LED_RoundFunction0_Feedback_7_), .B(
        Key0[71]), .ZN(LED_RoundFunction0_n417) );
  XNOR2_X1 LED_RoundFunction0_U200 ( .A(Plaintext0[7]), .B(Key0[7]), .ZN(
        LED_RoundFunction0_n418) );
  AOI22_X1 LED_RoundFunction0_U199 ( .A1(rst), .A2(LED_RoundFunction0_n416), 
        .B1(LED_RoundFunction0_n415), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[6]) );
  XNOR2_X1 LED_RoundFunction0_U198 ( .A(LED_RoundFunction0_Feedback_6_), .B(
        Key0[70]), .ZN(LED_RoundFunction0_n415) );
  XNOR2_X1 LED_RoundFunction0_U197 ( .A(Plaintext0[6]), .B(Key0[6]), .ZN(
        LED_RoundFunction0_n416) );
  AOI22_X1 LED_RoundFunction0_U196 ( .A1(rst), .A2(LED_RoundFunction0_n414), 
        .B1(LED_RoundFunction0_n413), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[63]) );
  XNOR2_X1 LED_RoundFunction0_U195 ( .A(LED_RoundFunction0_Feedback_63_), .B(
        Key0[127]), .ZN(LED_RoundFunction0_n413) );
  XNOR2_X1 LED_RoundFunction0_U194 ( .A(Plaintext0[63]), .B(Key0[63]), .ZN(
        LED_RoundFunction0_n414) );
  AOI22_X1 LED_RoundFunction0_U193 ( .A1(rst), .A2(LED_RoundFunction0_n412), 
        .B1(LED_RoundFunction0_n411), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[5]) );
  XNOR2_X1 LED_RoundFunction0_U192 ( .A(LED_RoundFunction0_Feedback_5_), .B(
        Key0[69]), .ZN(LED_RoundFunction0_n411) );
  XNOR2_X1 LED_RoundFunction0_U191 ( .A(Plaintext0[5]), .B(Key0[5]), .ZN(
        LED_RoundFunction0_n412) );
  AOI22_X1 LED_RoundFunction0_U190 ( .A1(rst), .A2(LED_RoundFunction0_n410), 
        .B1(LED_RoundFunction0_n409), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[58]) );
  XNOR2_X1 LED_RoundFunction0_U189 ( .A(LED_RoundFunction0_Feedback_58_), .B(
        Key0[122]), .ZN(LED_RoundFunction0_n409) );
  XNOR2_X1 LED_RoundFunction0_U188 ( .A(Plaintext0[58]), .B(Key0[58]), .ZN(
        LED_RoundFunction0_n410) );
  AOI22_X1 LED_RoundFunction0_U187 ( .A1(rst), .A2(LED_RoundFunction0_n408), 
        .B1(LED_RoundFunction0_n407), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[57]) );
  XNOR2_X1 LED_RoundFunction0_U186 ( .A(LED_RoundFunction0_Feedback_57_), .B(
        Key0[121]), .ZN(LED_RoundFunction0_n407) );
  XNOR2_X1 LED_RoundFunction0_U185 ( .A(Plaintext0[57]), .B(Key0[57]), .ZN(
        LED_RoundFunction0_n408) );
  AOI22_X1 LED_RoundFunction0_U184 ( .A1(rst), .A2(LED_RoundFunction0_n406), 
        .B1(LED_RoundFunction0_n405), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[56]) );
  XNOR2_X1 LED_RoundFunction0_U183 ( .A(LED_RoundFunction0_Feedback_56_), .B(
        Key0[120]), .ZN(LED_RoundFunction0_n405) );
  XNOR2_X1 LED_RoundFunction0_U182 ( .A(Plaintext0[56]), .B(Key0[56]), .ZN(
        LED_RoundFunction0_n406) );
  AOI22_X1 LED_RoundFunction0_U181 ( .A1(rst), .A2(LED_RoundFunction0_n404), 
        .B1(LED_RoundFunction0_n403), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[55]) );
  XNOR2_X1 LED_RoundFunction0_U180 ( .A(LED_RoundFunction0_Feedback_55_), .B(
        Key0[119]), .ZN(LED_RoundFunction0_n403) );
  XNOR2_X1 LED_RoundFunction0_U179 ( .A(Plaintext0[55]), .B(Key0[55]), .ZN(
        LED_RoundFunction0_n404) );
  AOI22_X1 LED_RoundFunction0_U178 ( .A1(rst), .A2(LED_RoundFunction0_n402), 
        .B1(LED_RoundFunction0_n401), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[54]) );
  XNOR2_X1 LED_RoundFunction0_U177 ( .A(LED_RoundFunction0_Feedback_54_), .B(
        Key0[118]), .ZN(LED_RoundFunction0_n401) );
  XNOR2_X1 LED_RoundFunction0_U176 ( .A(Plaintext0[54]), .B(Key0[54]), .ZN(
        LED_RoundFunction0_n402) );
  AOI22_X1 LED_RoundFunction0_U175 ( .A1(rst), .A2(LED_RoundFunction0_n400), 
        .B1(LED_RoundFunction0_n399), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[53]) );
  XNOR2_X1 LED_RoundFunction0_U174 ( .A(LED_RoundFunction0_Feedback_53_), .B(
        Key0[117]), .ZN(LED_RoundFunction0_n399) );
  XNOR2_X1 LED_RoundFunction0_U173 ( .A(Plaintext0[53]), .B(Key0[53]), .ZN(
        LED_RoundFunction0_n400) );
  AOI22_X1 LED_RoundFunction0_U172 ( .A1(rst), .A2(LED_RoundFunction0_n398), 
        .B1(LED_RoundFunction0_n397), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[52]) );
  XNOR2_X1 LED_RoundFunction0_U171 ( .A(LED_RoundFunction0_Feedback_52_), .B(
        Key0[116]), .ZN(LED_RoundFunction0_n397) );
  XNOR2_X1 LED_RoundFunction0_U170 ( .A(Plaintext0[52]), .B(Key0[52]), .ZN(
        LED_RoundFunction0_n398) );
  AOI22_X1 LED_RoundFunction0_U169 ( .A1(rst), .A2(LED_RoundFunction0_n396), 
        .B1(LED_RoundFunction0_n395), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[51]) );
  XNOR2_X1 LED_RoundFunction0_U168 ( .A(LED_RoundFunction0_Feedback_51_), .B(
        Key0[115]), .ZN(LED_RoundFunction0_n395) );
  XNOR2_X1 LED_RoundFunction0_U167 ( .A(Plaintext0[51]), .B(Key0[51]), .ZN(
        LED_RoundFunction0_n396) );
  AOI22_X1 LED_RoundFunction0_U166 ( .A1(rst), .A2(LED_RoundFunction0_n394), 
        .B1(LED_RoundFunction0_n393), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[50]) );
  XNOR2_X1 LED_RoundFunction0_U165 ( .A(LED_RoundFunction0_Feedback_50_), .B(
        Key0[114]), .ZN(LED_RoundFunction0_n393) );
  XNOR2_X1 LED_RoundFunction0_U164 ( .A(Plaintext0[50]), .B(Key0[50]), .ZN(
        LED_RoundFunction0_n394) );
  AOI22_X1 LED_RoundFunction0_U163 ( .A1(rst), .A2(LED_RoundFunction0_n392), 
        .B1(LED_RoundFunction0_n391), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[4]) );
  XNOR2_X1 LED_RoundFunction0_U162 ( .A(LED_RoundFunction0_Feedback_4_), .B(
        Key0[68]), .ZN(LED_RoundFunction0_n391) );
  XNOR2_X1 LED_RoundFunction0_U161 ( .A(Plaintext0[4]), .B(Key0[4]), .ZN(
        LED_RoundFunction0_n392) );
  AOI22_X1 LED_RoundFunction0_U160 ( .A1(rst), .A2(LED_RoundFunction0_n390), 
        .B1(LED_RoundFunction0_n389), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[49]) );
  XNOR2_X1 LED_RoundFunction0_U159 ( .A(LED_RoundFunction0_Feedback_49_), .B(
        Key0[113]), .ZN(LED_RoundFunction0_n389) );
  XNOR2_X1 LED_RoundFunction0_U158 ( .A(Plaintext0[49]), .B(Key0[49]), .ZN(
        LED_RoundFunction0_n390) );
  AOI22_X1 LED_RoundFunction0_U157 ( .A1(rst), .A2(LED_RoundFunction0_n388), 
        .B1(LED_RoundFunction0_n387), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[48]) );
  XNOR2_X1 LED_RoundFunction0_U156 ( .A(LED_RoundFunction0_Feedback_48_), .B(
        Key0[112]), .ZN(LED_RoundFunction0_n387) );
  XNOR2_X1 LED_RoundFunction0_U155 ( .A(Plaintext0[48]), .B(Key0[48]), .ZN(
        LED_RoundFunction0_n388) );
  AOI22_X1 LED_RoundFunction0_U154 ( .A1(rst), .A2(LED_RoundFunction0_n386), 
        .B1(LED_RoundFunction0_n385), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[47]) );
  XNOR2_X1 LED_RoundFunction0_U153 ( .A(LED_RoundFunction0_Feedback_47_), .B(
        Key0[111]), .ZN(LED_RoundFunction0_n385) );
  XNOR2_X1 LED_RoundFunction0_U152 ( .A(Plaintext0[47]), .B(Key0[47]), .ZN(
        LED_RoundFunction0_n386) );
  AOI22_X1 LED_RoundFunction0_U151 ( .A1(rst), .A2(LED_RoundFunction0_n384), 
        .B1(LED_RoundFunction0_n383), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[44]) );
  XNOR2_X1 LED_RoundFunction0_U150 ( .A(LED_RoundFunction0_Feedback_44_), .B(
        Key0[108]), .ZN(LED_RoundFunction0_n383) );
  XNOR2_X1 LED_RoundFunction0_U149 ( .A(Plaintext0[44]), .B(Key0[44]), .ZN(
        LED_RoundFunction0_n384) );
  AOI22_X1 LED_RoundFunction0_U148 ( .A1(rst), .A2(LED_RoundFunction0_n382), 
        .B1(LED_RoundFunction0_n381), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[42]) );
  XNOR2_X1 LED_RoundFunction0_U147 ( .A(LED_RoundFunction0_Feedback_42_), .B(
        Key0[106]), .ZN(LED_RoundFunction0_n381) );
  XNOR2_X1 LED_RoundFunction0_U146 ( .A(Plaintext0[42]), .B(Key0[42]), .ZN(
        LED_RoundFunction0_n382) );
  AOI22_X1 LED_RoundFunction0_U145 ( .A1(rst), .A2(LED_RoundFunction0_n380), 
        .B1(LED_RoundFunction0_n379), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[41]) );
  XNOR2_X1 LED_RoundFunction0_U144 ( .A(LED_RoundFunction0_Feedback_41_), .B(
        Key0[105]), .ZN(LED_RoundFunction0_n379) );
  XNOR2_X1 LED_RoundFunction0_U143 ( .A(Plaintext0[41]), .B(Key0[41]), .ZN(
        LED_RoundFunction0_n380) );
  AOI22_X1 LED_RoundFunction0_U142 ( .A1(rst), .A2(LED_RoundFunction0_n378), 
        .B1(LED_RoundFunction0_n377), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[40]) );
  XNOR2_X1 LED_RoundFunction0_U141 ( .A(LED_RoundFunction0_Feedback_40_), .B(
        Key0[104]), .ZN(LED_RoundFunction0_n377) );
  XNOR2_X1 LED_RoundFunction0_U140 ( .A(Plaintext0[40]), .B(Key0[40]), .ZN(
        LED_RoundFunction0_n378) );
  AOI22_X1 LED_RoundFunction0_U139 ( .A1(rst), .A2(LED_RoundFunction0_n376), 
        .B1(LED_RoundFunction0_n375), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[3]) );
  XNOR2_X1 LED_RoundFunction0_U138 ( .A(LED_RoundFunction0_Feedback_3_), .B(
        Key0[67]), .ZN(LED_RoundFunction0_n375) );
  XNOR2_X1 LED_RoundFunction0_U137 ( .A(Plaintext0[3]), .B(Key0[3]), .ZN(
        LED_RoundFunction0_n376) );
  AOI22_X1 LED_RoundFunction0_U136 ( .A1(rst), .A2(LED_RoundFunction0_n374), 
        .B1(LED_RoundFunction0_n373), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[39]) );
  XNOR2_X1 LED_RoundFunction0_U135 ( .A(LED_RoundFunction0_Feedback_39_), .B(
        Key0[103]), .ZN(LED_RoundFunction0_n373) );
  XNOR2_X1 LED_RoundFunction0_U134 ( .A(Plaintext0[39]), .B(Key0[39]), .ZN(
        LED_RoundFunction0_n374) );
  AOI22_X1 LED_RoundFunction0_U133 ( .A1(rst), .A2(LED_RoundFunction0_n372), 
        .B1(LED_RoundFunction0_n371), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[38]) );
  XNOR2_X1 LED_RoundFunction0_U132 ( .A(LED_RoundFunction0_Feedback_38_), .B(
        Key0[102]), .ZN(LED_RoundFunction0_n371) );
  XNOR2_X1 LED_RoundFunction0_U131 ( .A(Plaintext0[38]), .B(Key0[38]), .ZN(
        LED_RoundFunction0_n372) );
  AOI22_X1 LED_RoundFunction0_U130 ( .A1(rst), .A2(LED_RoundFunction0_n370), 
        .B1(LED_RoundFunction0_n369), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[37]) );
  XNOR2_X1 LED_RoundFunction0_U129 ( .A(LED_RoundFunction0_Feedback_37_), .B(
        Key0[101]), .ZN(LED_RoundFunction0_n369) );
  XNOR2_X1 LED_RoundFunction0_U128 ( .A(Plaintext0[37]), .B(Key0[37]), .ZN(
        LED_RoundFunction0_n370) );
  AOI22_X1 LED_RoundFunction0_U127 ( .A1(rst), .A2(LED_RoundFunction0_n368), 
        .B1(LED_RoundFunction0_n367), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[36]) );
  XNOR2_X1 LED_RoundFunction0_U126 ( .A(LED_RoundFunction0_Feedback_36_), .B(
        Key0[100]), .ZN(LED_RoundFunction0_n367) );
  XNOR2_X1 LED_RoundFunction0_U125 ( .A(Plaintext0[36]), .B(Key0[36]), .ZN(
        LED_RoundFunction0_n368) );
  AOI22_X1 LED_RoundFunction0_U124 ( .A1(rst), .A2(LED_RoundFunction0_n366), 
        .B1(LED_RoundFunction0_n365), .B2(LED_RoundFunction0_n294), .ZN(
        Ciphertext0[35]) );
  XNOR2_X1 LED_RoundFunction0_U123 ( .A(LED_RoundFunction0_Feedback_35_), .B(
        Key0[99]), .ZN(LED_RoundFunction0_n365) );
  XNOR2_X1 LED_RoundFunction0_U122 ( .A(Plaintext0[35]), .B(Key0[35]), .ZN(
        LED_RoundFunction0_n366) );
  AOI22_X1 LED_RoundFunction0_U121 ( .A1(rst), .A2(LED_RoundFunction0_n364), 
        .B1(LED_RoundFunction0_n363), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[34]) );
  XNOR2_X1 LED_RoundFunction0_U120 ( .A(LED_RoundFunction0_Feedback_34_), .B(
        Key0[98]), .ZN(LED_RoundFunction0_n363) );
  XNOR2_X1 LED_RoundFunction0_U119 ( .A(Plaintext0[34]), .B(Key0[34]), .ZN(
        LED_RoundFunction0_n364) );
  AOI22_X1 LED_RoundFunction0_U118 ( .A1(rst), .A2(LED_RoundFunction0_n362), 
        .B1(LED_RoundFunction0_n361), .B2(LED_RoundFunction0_n294), .ZN(
        Ciphertext0[33]) );
  XNOR2_X1 LED_RoundFunction0_U117 ( .A(LED_RoundFunction0_Feedback_33_), .B(
        Key0[97]), .ZN(LED_RoundFunction0_n361) );
  XNOR2_X1 LED_RoundFunction0_U116 ( .A(Plaintext0[33]), .B(Key0[33]), .ZN(
        LED_RoundFunction0_n362) );
  AOI22_X1 LED_RoundFunction0_U115 ( .A1(rst), .A2(LED_RoundFunction0_n360), 
        .B1(LED_RoundFunction0_n359), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[32]) );
  XNOR2_X1 LED_RoundFunction0_U114 ( .A(LED_RoundFunction0_Feedback_32_), .B(
        Key0[96]), .ZN(LED_RoundFunction0_n359) );
  XNOR2_X1 LED_RoundFunction0_U113 ( .A(Plaintext0[32]), .B(Key0[32]), .ZN(
        LED_RoundFunction0_n360) );
  AOI22_X1 LED_RoundFunction0_U112 ( .A1(rst), .A2(LED_RoundFunction0_n358), 
        .B1(LED_RoundFunction0_n357), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[2]) );
  XNOR2_X1 LED_RoundFunction0_U111 ( .A(LED_RoundFunction0_Feedback_2_), .B(
        Key0[66]), .ZN(LED_RoundFunction0_n357) );
  XNOR2_X1 LED_RoundFunction0_U110 ( .A(Plaintext0[2]), .B(Key0[2]), .ZN(
        LED_RoundFunction0_n358) );
  AOI22_X1 LED_RoundFunction0_U109 ( .A1(rst), .A2(LED_RoundFunction0_n356), 
        .B1(LED_RoundFunction0_n355), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[29]) );
  XNOR2_X1 LED_RoundFunction0_U108 ( .A(LED_RoundFunction0_Feedback_29_), .B(
        Key0[93]), .ZN(LED_RoundFunction0_n355) );
  XNOR2_X1 LED_RoundFunction0_U107 ( .A(Plaintext0[29]), .B(Key0[29]), .ZN(
        LED_RoundFunction0_n356) );
  AOI22_X1 LED_RoundFunction0_U106 ( .A1(rst), .A2(LED_RoundFunction0_n354), 
        .B1(LED_RoundFunction0_n353), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[26]) );
  XNOR2_X1 LED_RoundFunction0_U105 ( .A(LED_RoundFunction0_Feedback_26_), .B(
        Key0[90]), .ZN(LED_RoundFunction0_n353) );
  XNOR2_X1 LED_RoundFunction0_U104 ( .A(Plaintext0[26]), .B(Key0[26]), .ZN(
        LED_RoundFunction0_n354) );
  AOI22_X1 LED_RoundFunction0_U103 ( .A1(rst), .A2(LED_RoundFunction0_n352), 
        .B1(LED_RoundFunction0_n351), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[25]) );
  XNOR2_X1 LED_RoundFunction0_U102 ( .A(LED_RoundFunction0_Feedback_25_), .B(
        Key0[89]), .ZN(LED_RoundFunction0_n351) );
  XNOR2_X1 LED_RoundFunction0_U101 ( .A(Plaintext0[25]), .B(Key0[25]), .ZN(
        LED_RoundFunction0_n352) );
  AOI22_X1 LED_RoundFunction0_U100 ( .A1(rst), .A2(LED_RoundFunction0_n350), 
        .B1(LED_RoundFunction0_n349), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[24]) );
  XNOR2_X1 LED_RoundFunction0_U99 ( .A(LED_RoundFunction0_Feedback_24_), .B(
        Key0[88]), .ZN(LED_RoundFunction0_n349) );
  XNOR2_X1 LED_RoundFunction0_U98 ( .A(Plaintext0[24]), .B(Key0[24]), .ZN(
        LED_RoundFunction0_n350) );
  AOI22_X1 LED_RoundFunction0_U97 ( .A1(rst), .A2(LED_RoundFunction0_n348), 
        .B1(LED_RoundFunction0_n347), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[23]) );
  XNOR2_X1 LED_RoundFunction0_U96 ( .A(LED_RoundFunction0_Feedback_23_), .B(
        Key0[87]), .ZN(LED_RoundFunction0_n347) );
  XNOR2_X1 LED_RoundFunction0_U95 ( .A(Plaintext0[23]), .B(Key0[23]), .ZN(
        LED_RoundFunction0_n348) );
  AOI22_X1 LED_RoundFunction0_U94 ( .A1(rst), .A2(LED_RoundFunction0_n346), 
        .B1(LED_RoundFunction0_n345), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[22]) );
  XNOR2_X1 LED_RoundFunction0_U93 ( .A(LED_RoundFunction0_Feedback_22_), .B(
        Key0[86]), .ZN(LED_RoundFunction0_n345) );
  XNOR2_X1 LED_RoundFunction0_U92 ( .A(Plaintext0[22]), .B(Key0[22]), .ZN(
        LED_RoundFunction0_n346) );
  AOI22_X1 LED_RoundFunction0_U91 ( .A1(rst), .A2(LED_RoundFunction0_n344), 
        .B1(LED_RoundFunction0_n343), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[21]) );
  XNOR2_X1 LED_RoundFunction0_U90 ( .A(LED_RoundFunction0_Feedback_21_), .B(
        Key0[85]), .ZN(LED_RoundFunction0_n343) );
  XNOR2_X1 LED_RoundFunction0_U89 ( .A(Plaintext0[21]), .B(Key0[21]), .ZN(
        LED_RoundFunction0_n344) );
  AOI22_X1 LED_RoundFunction0_U88 ( .A1(rst), .A2(LED_RoundFunction0_n342), 
        .B1(LED_RoundFunction0_n341), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[20]) );
  XNOR2_X1 LED_RoundFunction0_U87 ( .A(LED_RoundFunction0_Feedback_20_), .B(
        Key0[84]), .ZN(LED_RoundFunction0_n341) );
  XNOR2_X1 LED_RoundFunction0_U86 ( .A(Plaintext0[20]), .B(Key0[20]), .ZN(
        LED_RoundFunction0_n342) );
  AOI22_X1 LED_RoundFunction0_U85 ( .A1(rst), .A2(LED_RoundFunction0_n340), 
        .B1(LED_RoundFunction0_n339), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[1]) );
  XNOR2_X1 LED_RoundFunction0_U84 ( .A(LED_RoundFunction0_Feedback_1_), .B(
        Key0[65]), .ZN(LED_RoundFunction0_n339) );
  XNOR2_X1 LED_RoundFunction0_U83 ( .A(Plaintext0[1]), .B(Key0[1]), .ZN(
        LED_RoundFunction0_n340) );
  AOI22_X1 LED_RoundFunction0_U82 ( .A1(rst), .A2(LED_RoundFunction0_n338), 
        .B1(LED_RoundFunction0_n337), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[19]) );
  XNOR2_X1 LED_RoundFunction0_U81 ( .A(LED_RoundFunction0_Feedback_19_), .B(
        Key0[83]), .ZN(LED_RoundFunction0_n337) );
  XNOR2_X1 LED_RoundFunction0_U80 ( .A(Plaintext0[19]), .B(Key0[19]), .ZN(
        LED_RoundFunction0_n338) );
  AOI22_X1 LED_RoundFunction0_U79 ( .A1(rst), .A2(LED_RoundFunction0_n336), 
        .B1(LED_RoundFunction0_n335), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[18]) );
  XNOR2_X1 LED_RoundFunction0_U78 ( .A(LED_RoundFunction0_Feedback_18_), .B(
        Key0[82]), .ZN(LED_RoundFunction0_n335) );
  XNOR2_X1 LED_RoundFunction0_U77 ( .A(Plaintext0[18]), .B(Key0[18]), .ZN(
        LED_RoundFunction0_n336) );
  AOI22_X1 LED_RoundFunction0_U76 ( .A1(rst), .A2(LED_RoundFunction0_n334), 
        .B1(LED_RoundFunction0_n333), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[17]) );
  XNOR2_X1 LED_RoundFunction0_U75 ( .A(LED_RoundFunction0_Feedback_17_), .B(
        Key0[81]), .ZN(LED_RoundFunction0_n333) );
  XNOR2_X1 LED_RoundFunction0_U74 ( .A(Plaintext0[17]), .B(Key0[17]), .ZN(
        LED_RoundFunction0_n334) );
  AOI22_X1 LED_RoundFunction0_U73 ( .A1(rst), .A2(LED_RoundFunction0_n332), 
        .B1(LED_RoundFunction0_n331), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[16]) );
  XNOR2_X1 LED_RoundFunction0_U72 ( .A(LED_RoundFunction0_Feedback_16_), .B(
        Key0[80]), .ZN(LED_RoundFunction0_n331) );
  XNOR2_X1 LED_RoundFunction0_U71 ( .A(Plaintext0[16]), .B(Key0[16]), .ZN(
        LED_RoundFunction0_n332) );
  AOI22_X1 LED_RoundFunction0_U70 ( .A1(rst), .A2(LED_RoundFunction0_n330), 
        .B1(LED_RoundFunction0_n329), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[13]) );
  XNOR2_X1 LED_RoundFunction0_U69 ( .A(LED_RoundFunction0_Feedback_13_), .B(
        Key0[77]), .ZN(LED_RoundFunction0_n329) );
  XNOR2_X1 LED_RoundFunction0_U68 ( .A(Plaintext0[13]), .B(Key0[13]), .ZN(
        LED_RoundFunction0_n330) );
  AOI22_X1 LED_RoundFunction0_U67 ( .A1(rst), .A2(LED_RoundFunction0_n328), 
        .B1(LED_RoundFunction0_n327), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[12]) );
  XNOR2_X1 LED_RoundFunction0_U66 ( .A(LED_RoundFunction0_Feedback_12_), .B(
        Key0[76]), .ZN(LED_RoundFunction0_n327) );
  XNOR2_X1 LED_RoundFunction0_U65 ( .A(Plaintext0[12]), .B(Key0[12]), .ZN(
        LED_RoundFunction0_n328) );
  AOI22_X1 LED_RoundFunction0_U64 ( .A1(rst), .A2(LED_RoundFunction0_n326), 
        .B1(LED_RoundFunction0_n325), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[10]) );
  XNOR2_X1 LED_RoundFunction0_U63 ( .A(LED_RoundFunction0_Feedback_10_), .B(
        Key0[74]), .ZN(LED_RoundFunction0_n325) );
  XNOR2_X1 LED_RoundFunction0_U62 ( .A(Plaintext0[10]), .B(Key0[10]), .ZN(
        LED_RoundFunction0_n326) );
  AOI22_X1 LED_RoundFunction0_U61 ( .A1(rst), .A2(LED_RoundFunction0_n324), 
        .B1(LED_RoundFunction0_n323), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[0]) );
  XNOR2_X1 LED_RoundFunction0_U60 ( .A(LED_RoundFunction0_Feedback_0_), .B(
        Key0[64]), .ZN(LED_RoundFunction0_n323) );
  XNOR2_X1 LED_RoundFunction0_U59 ( .A(Plaintext0[0]), .B(Key0[0]), .ZN(
        LED_RoundFunction0_n324) );
  AOI22_X1 LED_RoundFunction0_U58 ( .A1(rst), .A2(LED_RoundFunction0_n322), 
        .B1(LED_RoundFunction0_n321), .B2(LED_RoundFunction0_n294), .ZN(
        Ciphertext0[46]) );
  XNOR2_X1 LED_RoundFunction0_U57 ( .A(LED_RoundFunction0_Feedback_46_), .B(
        Key0[110]), .ZN(LED_RoundFunction0_n321) );
  XNOR2_X1 LED_RoundFunction0_U56 ( .A(Plaintext0[46]), .B(Key0[46]), .ZN(
        LED_RoundFunction0_n322) );
  AOI22_X1 LED_RoundFunction0_U55 ( .A1(rst), .A2(LED_RoundFunction0_n320), 
        .B1(LED_RoundFunction0_n319), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[45]) );
  XNOR2_X1 LED_RoundFunction0_U54 ( .A(LED_RoundFunction0_Feedback_45_), .B(
        Key0[109]), .ZN(LED_RoundFunction0_n319) );
  XNOR2_X1 LED_RoundFunction0_U53 ( .A(Plaintext0[45]), .B(Key0[45]), .ZN(
        LED_RoundFunction0_n320) );
  AOI22_X1 LED_RoundFunction0_U52 ( .A1(rst), .A2(LED_RoundFunction0_n318), 
        .B1(LED_RoundFunction0_n317), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[43]) );
  XNOR2_X1 LED_RoundFunction0_U51 ( .A(LED_RoundFunction0_Feedback_43_), .B(
        Key0[107]), .ZN(LED_RoundFunction0_n317) );
  XNOR2_X1 LED_RoundFunction0_U50 ( .A(Plaintext0[43]), .B(Key0[43]), .ZN(
        LED_RoundFunction0_n318) );
  AOI22_X1 LED_RoundFunction0_U49 ( .A1(rst), .A2(LED_RoundFunction0_n316), 
        .B1(LED_RoundFunction0_n315), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[31]) );
  XNOR2_X1 LED_RoundFunction0_U48 ( .A(LED_RoundFunction0_Feedback_31_), .B(
        Key0[95]), .ZN(LED_RoundFunction0_n315) );
  XNOR2_X1 LED_RoundFunction0_U47 ( .A(Plaintext0[31]), .B(Key0[31]), .ZN(
        LED_RoundFunction0_n316) );
  AOI22_X1 LED_RoundFunction0_U46 ( .A1(rst), .A2(LED_RoundFunction0_n314), 
        .B1(LED_RoundFunction0_n313), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[30]) );
  XNOR2_X1 LED_RoundFunction0_U45 ( .A(LED_RoundFunction0_Feedback_30_), .B(
        Key0[94]), .ZN(LED_RoundFunction0_n313) );
  XNOR2_X1 LED_RoundFunction0_U44 ( .A(Plaintext0[30]), .B(Key0[30]), .ZN(
        LED_RoundFunction0_n314) );
  AOI22_X1 LED_RoundFunction0_U43 ( .A1(rst), .A2(LED_RoundFunction0_n312), 
        .B1(LED_RoundFunction0_n311), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[28]) );
  XNOR2_X1 LED_RoundFunction0_U42 ( .A(LED_RoundFunction0_Feedback_28_), .B(
        Key0[92]), .ZN(LED_RoundFunction0_n311) );
  XNOR2_X1 LED_RoundFunction0_U41 ( .A(Plaintext0[28]), .B(Key0[28]), .ZN(
        LED_RoundFunction0_n312) );
  AOI22_X1 LED_RoundFunction0_U40 ( .A1(rst), .A2(LED_RoundFunction0_n310), 
        .B1(LED_RoundFunction0_n309), .B2(LED_RoundFunction0_n290), .ZN(
        Ciphertext0[27]) );
  XNOR2_X1 LED_RoundFunction0_U39 ( .A(LED_RoundFunction0_Feedback_27_), .B(
        Key0[91]), .ZN(LED_RoundFunction0_n309) );
  XNOR2_X1 LED_RoundFunction0_U38 ( .A(Plaintext0[27]), .B(Key0[27]), .ZN(
        LED_RoundFunction0_n310) );
  AOI22_X1 LED_RoundFunction0_U37 ( .A1(rst), .A2(LED_RoundFunction0_n308), 
        .B1(LED_RoundFunction0_n307), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[15]) );
  XNOR2_X1 LED_RoundFunction0_U36 ( .A(LED_RoundFunction0_Feedback_15_), .B(
        Key0[79]), .ZN(LED_RoundFunction0_n307) );
  XNOR2_X1 LED_RoundFunction0_U35 ( .A(Plaintext0[15]), .B(Key0[15]), .ZN(
        LED_RoundFunction0_n308) );
  AOI22_X1 LED_RoundFunction0_U34 ( .A1(rst), .A2(LED_RoundFunction0_n306), 
        .B1(LED_RoundFunction0_n305), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[14]) );
  XNOR2_X1 LED_RoundFunction0_U33 ( .A(LED_RoundFunction0_Feedback_14_), .B(
        Key0[78]), .ZN(LED_RoundFunction0_n305) );
  XNOR2_X1 LED_RoundFunction0_U32 ( .A(Plaintext0[14]), .B(Key0[14]), .ZN(
        LED_RoundFunction0_n306) );
  AOI22_X1 LED_RoundFunction0_U31 ( .A1(rst), .A2(LED_RoundFunction0_n304), 
        .B1(LED_RoundFunction0_n303), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[11]) );
  XNOR2_X1 LED_RoundFunction0_U30 ( .A(LED_RoundFunction0_Feedback_11_), .B(
        Key0[75]), .ZN(LED_RoundFunction0_n303) );
  XNOR2_X1 LED_RoundFunction0_U29 ( .A(Plaintext0[11]), .B(Key0[11]), .ZN(
        LED_RoundFunction0_n304) );
  AOI22_X1 LED_RoundFunction0_U28 ( .A1(rst), .A2(LED_RoundFunction0_n302), 
        .B1(LED_RoundFunction0_n301), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[62]) );
  XNOR2_X1 LED_RoundFunction0_U27 ( .A(LED_RoundFunction0_Feedback_62_), .B(
        Key0[126]), .ZN(LED_RoundFunction0_n301) );
  XNOR2_X1 LED_RoundFunction0_U26 ( .A(Plaintext0[62]), .B(Key0[62]), .ZN(
        LED_RoundFunction0_n302) );
  AOI22_X1 LED_RoundFunction0_U25 ( .A1(rst), .A2(LED_RoundFunction0_n300), 
        .B1(LED_RoundFunction0_n299), .B2(LED_RoundFunction0_n291), .ZN(
        Ciphertext0[61]) );
  XNOR2_X1 LED_RoundFunction0_U24 ( .A(LED_RoundFunction0_Feedback_61_), .B(
        Key0[125]), .ZN(LED_RoundFunction0_n299) );
  XNOR2_X1 LED_RoundFunction0_U23 ( .A(Plaintext0[61]), .B(Key0[61]), .ZN(
        LED_RoundFunction0_n300) );
  AOI22_X1 LED_RoundFunction0_U22 ( .A1(rst), .A2(LED_RoundFunction0_n298), 
        .B1(LED_RoundFunction0_n297), .B2(LED_RoundFunction0_n292), .ZN(
        Ciphertext0[60]) );
  XNOR2_X1 LED_RoundFunction0_U21 ( .A(LED_RoundFunction0_Feedback_60_), .B(
        Key0[124]), .ZN(LED_RoundFunction0_n297) );
  XNOR2_X1 LED_RoundFunction0_U20 ( .A(Plaintext0[60]), .B(Key0[60]), .ZN(
        LED_RoundFunction0_n298) );
  AOI22_X1 LED_RoundFunction0_U19 ( .A1(rst), .A2(LED_RoundFunction0_n296), 
        .B1(LED_RoundFunction0_n295), .B2(LED_RoundFunction0_n293), .ZN(
        Ciphertext0[59]) );
  XNOR2_X1 LED_RoundFunction0_U18 ( .A(LED_RoundFunction0_Feedback_59_), .B(
        Key0[123]), .ZN(LED_RoundFunction0_n295) );
  XNOR2_X1 LED_RoundFunction0_U17 ( .A(Plaintext0[59]), .B(Key0[59]), .ZN(
        LED_RoundFunction0_n296) );
  INV_X1 LED_RoundFunction0_U16 ( .A(LED_RoundFunction0_n285), .ZN(
        LED_RoundFunction0_n284) );
  INV_X1 LED_RoundFunction0_U15 ( .A(rst), .ZN(LED_RoundFunction0_n294) );
  BUF_X1 LED_RoundFunction0_U14 ( .A(LED_RoundFunction0_n294), .Z(
        LED_RoundFunction0_n292) );
  INV_X1 LED_RoundFunction0_U13 ( .A(LED_RoundFunction0_n285), .ZN(
        LED_RoundFunction0_n282) );
  BUF_X1 LED_RoundFunction0_U12 ( .A(LED_RoundFunction0_n294), .Z(
        LED_RoundFunction0_n291) );
  INV_X1 LED_RoundFunction0_U11 ( .A(LED_RoundFunction0_n285), .ZN(
        LED_RoundFunction0_n283) );
  BUF_X1 LED_RoundFunction0_U10 ( .A(LED_RoundFunction0_n294), .Z(
        LED_RoundFunction0_n290) );
  BUF_X1 LED_RoundFunction0_U9 ( .A(LED_RoundFunction0_n294), .Z(
        LED_RoundFunction0_n289) );
  INV_X1 LED_RoundFunction0_U8 ( .A(LED_RoundFunction0_n285), .ZN(
        LED_RoundFunction0_n281) );
  BUF_X1 LED_RoundFunction0_U7 ( .A(LED_RoundFunction0_n294), .Z(
        LED_RoundFunction0_n293) );
  BUF_X1 LED_RoundFunction0_U6 ( .A(LED_RoundFunction0_n287), .Z(
        LED_RoundFunction0_n286) );
  BUF_X1 LED_RoundFunction0_U5 ( .A(LED_RoundFunction0_n294), .Z(
        LED_RoundFunction0_n288) );
  INV_X1 LED_RoundFunction0_U4 ( .A(AddKey), .ZN(LED_RoundFunction0_n287) );
  BUF_X1 LED_RoundFunction0_U3 ( .A(LED_RoundFunction0_n287), .Z(
        LED_RoundFunction0_n285) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U68 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n160), .B(
        LED_RoundFunction0_MCInst1_MC0_n159), .ZN(
        LED_RoundFunction0_Feedback_15_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U67 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n158), .B(SubCellOutput0[62]), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n160) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U66 ( .A(SubCellOutput0[3]), .B(
        LED_RoundFunction0_MCInst1_MC0_n157), .Z(
        LED_RoundFunction0_Feedback_14_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U65 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n156), .B(
        LED_RoundFunction0_MCInst1_MC0_n155), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n157) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U64 ( .A(SubCellOutput0[21]), .B(
        SubCellOutput0[1]), .ZN(LED_RoundFunction0_MCInst1_MC0_n155) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U63 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n154), .B(SubCellOutput0[41]), .Z(
        LED_RoundFunction0_MCInst1_MC0_n156) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U62 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n153), .B(
        LED_RoundFunction0_MCInst1_MC0_n152), .ZN(
        LED_RoundFunction0_Feedback_13_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U61 ( .A(SubCellOutput0[2]), .B(
        SubCellOutput0[40]), .ZN(LED_RoundFunction0_MCInst1_MC0_n152) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U60 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n151), .B(
        LED_RoundFunction0_MCInst1_MC0_n150), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n153) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U59 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n149), .B(
        LED_RoundFunction0_MCInst1_MC0_n148), .ZN(
        LED_RoundFunction0_Feedback_12_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U58 ( .A(SubCellOutput0[23]), .B(
        LED_RoundFunction0_MCInst1_MC0_n147), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n148) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U57 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n146), .B(
        LED_RoundFunction0_MCInst1_MC0_n150), .Z(
        LED_RoundFunction0_MCInst1_MC0_n149) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U56 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n145), .B(
        LED_RoundFunction0_MCInst1_MC0_n159), .Z(
        LED_RoundFunction0_MCInst1_MC0_n150) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC0_U55 ( .A1(SubCellOutput0[21]), .A2(
        SubCellOutput0[22]), .B1(LED_RoundFunction0_MCInst1_MC0_n144), .B2(
        LED_RoundFunction0_MCInst1_MC0_n143), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n146) );
  INV_X1 LED_RoundFunction0_MCInst1_MC0_U54 ( .A(SubCellOutput0[21]), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n143) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U53 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n142), .B(
        LED_RoundFunction0_MCInst1_MC0_n141), .ZN(
        LED_RoundFunction0_Feedback_31_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U52 ( .A(SubCellOutput0[43]), .B(
        LED_RoundFunction0_MCInst1_MC0_n140), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n141) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U51 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n139), .B(SubCellOutput0[60]), .Z(
        LED_RoundFunction0_MCInst1_MC0_n142) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC0_U50 ( .A1(SubCellOutput0[42]), .A2(
        SubCellOutput0[22]), .B1(LED_RoundFunction0_MCInst1_MC0_n144), .B2(
        LED_RoundFunction0_MCInst1_MC0_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n139) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U49 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n137), .B(
        LED_RoundFunction0_MCInst1_MC0_n136), .ZN(
        LED_RoundFunction0_Feedback_30_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U48 ( .A(SubCellOutput0[40]), .B(
        LED_RoundFunction0_MCInst1_MC0_n135), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n136) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U47 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n134), .B(
        LED_RoundFunction0_MCInst1_MC0_n133), .Z(
        LED_RoundFunction0_MCInst1_MC0_n137) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC0_U46 ( .A1(SubCellOutput0[22]), .A2(
        SubCellOutput0[61]), .B1(LED_RoundFunction0_MCInst1_MC0_n132), .B2(
        LED_RoundFunction0_MCInst1_MC0_n144), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n134) );
  INV_X1 LED_RoundFunction0_MCInst1_MC0_U45 ( .A(SubCellOutput0[22]), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n144) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U44 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n131), .B(
        LED_RoundFunction0_MCInst1_MC0_n151), .ZN(
        LED_RoundFunction0_Feedback_29_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U43 ( .A(SubCellOutput0[63]), .B(
        SubCellOutput0[60]), .ZN(LED_RoundFunction0_MCInst1_MC0_n151) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U42 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n130), .B(
        LED_RoundFunction0_MCInst1_MC0_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n131) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U41 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n128), .B(
        LED_RoundFunction0_MCInst1_MC0_n127), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n130) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U40 ( .A(SubCellOutput0[21]), .B(
        LED_RoundFunction0_MCInst1_MC0_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n127) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U39 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n125), .B(SubCellOutput0[20]), .Z(
        LED_RoundFunction0_MCInst1_MC0_n128) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U38 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n124), .B(
        LED_RoundFunction0_MCInst1_MC0_n123), .ZN(
        LED_RoundFunction0_Feedback_28_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U37 ( .A(SubCellOutput0[0]), .B(
        LED_RoundFunction0_MCInst1_MC0_n122), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n124) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U36 ( .A(SubCellOutput0[2]), .B(
        LED_RoundFunction0_MCInst1_MC0_n122), .ZN(
        LED_RoundFunction0_Feedback_47_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U35 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n135), .B(
        LED_RoundFunction0_MCInst1_MC0_n121), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n122) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U34 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n120), .B(
        LED_RoundFunction0_MCInst1_MC0_n125), .Z(
        LED_RoundFunction0_MCInst1_MC0_n135) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U33 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n119), .B(
        LED_RoundFunction0_MCInst1_MC0_n118), .ZN(
        LED_RoundFunction0_Feedback_46_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U32 ( .A(SubCellOutput0[22]), .B(
        LED_RoundFunction0_MCInst1_MC0_n145), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n118) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U31 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n140), .B(
        LED_RoundFunction0_MCInst1_MC0_n147), .Z(
        LED_RoundFunction0_MCInst1_MC0_n119) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U30 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n126), .B(
        LED_RoundFunction0_MCInst1_MC0_n117), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n140) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U29 ( .A(SubCellOutput0[0]), .B(
        LED_RoundFunction0_MCInst1_MC0_n116), .ZN(
        LED_RoundFunction0_Feedback_45_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U28 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n115), .B(
        LED_RoundFunction0_MCInst1_MC0_n114), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n116) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U27 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n158), .B(SubCellOutput0[61]), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n115) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U26 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n120), .B(
        LED_RoundFunction0_MCInst1_MC0_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n158) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U25 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n113), .B(
        LED_RoundFunction0_MCInst1_MC0_n112), .ZN(
        LED_RoundFunction0_Feedback_44_) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC0_U24 ( .A1(SubCellOutput0[42]), .A2(
        LED_RoundFunction0_MCInst1_MC0_n111), .B1(
        LED_RoundFunction0_MCInst1_MC0_n129), .B2(
        LED_RoundFunction0_MCInst1_MC0_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n112) );
  INV_X1 LED_RoundFunction0_MCInst1_MC0_U23 ( .A(SubCellOutput0[42]), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n138) );
  INV_X1 LED_RoundFunction0_MCInst1_MC0_U22 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n111), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n129) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U21 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n145), .B(
        LED_RoundFunction0_MCInst1_MC0_n154), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n113) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC0_U20 ( .A1(SubCellOutput0[61]), .A2(
        SubCellOutput0[20]), .B1(LED_RoundFunction0_MCInst1_MC0_n110), .B2(
        LED_RoundFunction0_MCInst1_MC0_n132), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n154) );
  INV_X1 LED_RoundFunction0_MCInst1_MC0_U19 ( .A(SubCellOutput0[61]), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n132) );
  INV_X1 LED_RoundFunction0_MCInst1_MC0_U18 ( .A(SubCellOutput0[20]), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n110) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U17 ( .A(SubCellOutput0[3]), .B(
        SubCellOutput0[43]), .Z(LED_RoundFunction0_MCInst1_MC0_n145) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U16 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n111), .B(
        LED_RoundFunction0_MCInst1_MC0_n123), .ZN(
        LED_RoundFunction0_Feedback_63_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U15 ( .A(SubCellOutput0[61]), .B(
        SubCellOutput0[43]), .ZN(LED_RoundFunction0_MCInst1_MC0_n123) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U14 ( .A(SubCellOutput0[22]), .B(
        SubCellOutput0[2]), .Z(LED_RoundFunction0_MCInst1_MC0_n111) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U13 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n120), .B(
        LED_RoundFunction0_MCInst1_MC0_n121), .Z(
        LED_RoundFunction0_Feedback_62_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U12 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n147), .B(SubCellOutput0[60]), .Z(
        LED_RoundFunction0_MCInst1_MC0_n121) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U11 ( .A(SubCellOutput0[1]), .B(
        SubCellOutput0[63]), .Z(LED_RoundFunction0_MCInst1_MC0_n147) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U10 ( .A(SubCellOutput0[42]), .B(
        SubCellOutput0[21]), .Z(LED_RoundFunction0_MCInst1_MC0_n120) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U9 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n117), .B(
        LED_RoundFunction0_MCInst1_MC0_n109), .ZN(
        LED_RoundFunction0_Feedback_61_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U8 ( .A(SubCellOutput0[62]), .B(
        LED_RoundFunction0_MCInst1_MC0_n133), .Z(
        LED_RoundFunction0_MCInst1_MC0_n109) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U7 ( .A(SubCellOutput0[3]), .B(
        SubCellOutput0[63]), .Z(LED_RoundFunction0_MCInst1_MC0_n133) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U6 ( .A(
        LED_RoundFunction0_MCInst1_MC0_n159), .B(
        LED_RoundFunction0_MCInst1_MC0_n125), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n117) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U5 ( .A(SubCellOutput0[23]), .B(
        SubCellOutput0[41]), .Z(LED_RoundFunction0_MCInst1_MC0_n125) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U4 ( .A(SubCellOutput0[0]), .B(
        SubCellOutput0[20]), .Z(LED_RoundFunction0_MCInst1_MC0_n159) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U3 ( .A(SubCellOutput0[3]), .B(
        LED_RoundFunction0_MCInst1_MC0_n114), .ZN(
        LED_RoundFunction0_Feedback_60_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC0_U2 ( .A(SubCellOutput0[23]), .B(
        LED_RoundFunction0_MCInst1_MC0_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC0_n114) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC0_U1 ( .A(SubCellOutput0[62]), .B(
        SubCellOutput0[40]), .Z(LED_RoundFunction0_MCInst1_MC0_n126) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U68 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n160), .B(
        LED_RoundFunction0_MCInst1_MC1_n159), .ZN(
        LED_RoundFunction0_Feedback_11_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U67 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n158), .B(SubCellOutput0[58]), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n160) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U66 ( .A(SubCellOutput0[15]), .B(
        LED_RoundFunction0_MCInst1_MC1_n157), .Z(
        LED_RoundFunction0_Feedback_10_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U65 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n156), .B(
        LED_RoundFunction0_MCInst1_MC1_n155), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n157) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U64 ( .A(SubCellOutput0[17]), .B(
        SubCellOutput0[13]), .ZN(LED_RoundFunction0_MCInst1_MC1_n155) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U63 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n154), .B(SubCellOutput0[37]), .Z(
        LED_RoundFunction0_MCInst1_MC1_n156) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U62 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n153), .B(
        LED_RoundFunction0_MCInst1_MC1_n152), .ZN(
        LED_RoundFunction0_Feedback_9_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U61 ( .A(SubCellOutput0[14]), .B(
        SubCellOutput0[36]), .ZN(LED_RoundFunction0_MCInst1_MC1_n152) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U60 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n151), .B(
        LED_RoundFunction0_MCInst1_MC1_n150), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n153) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U59 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n149), .B(
        LED_RoundFunction0_MCInst1_MC1_n148), .ZN(
        LED_RoundFunction0_Feedback_8_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U58 ( .A(SubCellOutput0[19]), .B(
        LED_RoundFunction0_MCInst1_MC1_n147), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n148) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U57 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n146), .B(
        LED_RoundFunction0_MCInst1_MC1_n150), .Z(
        LED_RoundFunction0_MCInst1_MC1_n149) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U56 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n145), .B(
        LED_RoundFunction0_MCInst1_MC1_n159), .Z(
        LED_RoundFunction0_MCInst1_MC1_n150) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC1_U55 ( .A1(SubCellOutput0[17]), .A2(
        SubCellOutput0[18]), .B1(LED_RoundFunction0_MCInst1_MC1_n144), .B2(
        LED_RoundFunction0_MCInst1_MC1_n143), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n146) );
  INV_X1 LED_RoundFunction0_MCInst1_MC1_U54 ( .A(SubCellOutput0[17]), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n143) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U53 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n142), .B(
        LED_RoundFunction0_MCInst1_MC1_n141), .ZN(
        LED_RoundFunction0_Feedback_27_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U52 ( .A(SubCellOutput0[39]), .B(
        LED_RoundFunction0_MCInst1_MC1_n140), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n141) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U51 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n139), .B(SubCellOutput0[56]), .Z(
        LED_RoundFunction0_MCInst1_MC1_n142) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC1_U50 ( .A1(SubCellOutput0[38]), .A2(
        SubCellOutput0[18]), .B1(LED_RoundFunction0_MCInst1_MC1_n144), .B2(
        LED_RoundFunction0_MCInst1_MC1_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n139) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U49 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n137), .B(
        LED_RoundFunction0_MCInst1_MC1_n136), .ZN(
        LED_RoundFunction0_Feedback_26_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U48 ( .A(SubCellOutput0[36]), .B(
        LED_RoundFunction0_MCInst1_MC1_n135), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n136) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U47 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n134), .B(
        LED_RoundFunction0_MCInst1_MC1_n133), .Z(
        LED_RoundFunction0_MCInst1_MC1_n137) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC1_U46 ( .A1(SubCellOutput0[18]), .A2(
        SubCellOutput0[57]), .B1(LED_RoundFunction0_MCInst1_MC1_n132), .B2(
        LED_RoundFunction0_MCInst1_MC1_n144), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n134) );
  INV_X1 LED_RoundFunction0_MCInst1_MC1_U45 ( .A(SubCellOutput0[18]), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n144) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U44 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n131), .B(
        LED_RoundFunction0_MCInst1_MC1_n151), .ZN(
        LED_RoundFunction0_Feedback_25_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U43 ( .A(SubCellOutput0[59]), .B(
        SubCellOutput0[56]), .ZN(LED_RoundFunction0_MCInst1_MC1_n151) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U42 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n130), .B(
        LED_RoundFunction0_MCInst1_MC1_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n131) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U41 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n128), .B(
        LED_RoundFunction0_MCInst1_MC1_n127), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n130) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U40 ( .A(SubCellOutput0[17]), .B(
        LED_RoundFunction0_MCInst1_MC1_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n127) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U39 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n125), .B(SubCellOutput0[16]), .Z(
        LED_RoundFunction0_MCInst1_MC1_n128) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U38 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n124), .B(
        LED_RoundFunction0_MCInst1_MC1_n123), .ZN(
        LED_RoundFunction0_Feedback_24_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U37 ( .A(SubCellOutput0[12]), .B(
        LED_RoundFunction0_MCInst1_MC1_n122), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n124) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U36 ( .A(SubCellOutput0[14]), .B(
        LED_RoundFunction0_MCInst1_MC1_n122), .ZN(
        LED_RoundFunction0_Feedback_43_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U35 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n135), .B(
        LED_RoundFunction0_MCInst1_MC1_n121), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n122) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U34 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n120), .B(
        LED_RoundFunction0_MCInst1_MC1_n125), .Z(
        LED_RoundFunction0_MCInst1_MC1_n135) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U33 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n119), .B(
        LED_RoundFunction0_MCInst1_MC1_n118), .ZN(
        LED_RoundFunction0_Feedback_42_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U32 ( .A(SubCellOutput0[18]), .B(
        LED_RoundFunction0_MCInst1_MC1_n145), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n118) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U31 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n140), .B(
        LED_RoundFunction0_MCInst1_MC1_n147), .Z(
        LED_RoundFunction0_MCInst1_MC1_n119) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U30 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n126), .B(
        LED_RoundFunction0_MCInst1_MC1_n117), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n140) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U29 ( .A(SubCellOutput0[12]), .B(
        LED_RoundFunction0_MCInst1_MC1_n116), .ZN(
        LED_RoundFunction0_Feedback_41_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U28 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n115), .B(
        LED_RoundFunction0_MCInst1_MC1_n114), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n116) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U27 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n158), .B(SubCellOutput0[57]), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n115) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U26 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n120), .B(
        LED_RoundFunction0_MCInst1_MC1_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n158) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U25 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n113), .B(
        LED_RoundFunction0_MCInst1_MC1_n112), .ZN(
        LED_RoundFunction0_Feedback_40_) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC1_U24 ( .A1(SubCellOutput0[38]), .A2(
        LED_RoundFunction0_MCInst1_MC1_n111), .B1(
        LED_RoundFunction0_MCInst1_MC1_n129), .B2(
        LED_RoundFunction0_MCInst1_MC1_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n112) );
  INV_X1 LED_RoundFunction0_MCInst1_MC1_U23 ( .A(SubCellOutput0[38]), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n138) );
  INV_X1 LED_RoundFunction0_MCInst1_MC1_U22 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n111), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n129) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U21 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n145), .B(
        LED_RoundFunction0_MCInst1_MC1_n154), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n113) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC1_U20 ( .A1(SubCellOutput0[57]), .A2(
        SubCellOutput0[16]), .B1(LED_RoundFunction0_MCInst1_MC1_n110), .B2(
        LED_RoundFunction0_MCInst1_MC1_n132), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n154) );
  INV_X1 LED_RoundFunction0_MCInst1_MC1_U19 ( .A(SubCellOutput0[57]), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n132) );
  INV_X1 LED_RoundFunction0_MCInst1_MC1_U18 ( .A(SubCellOutput0[16]), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n110) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U17 ( .A(SubCellOutput0[15]), .B(
        SubCellOutput0[39]), .Z(LED_RoundFunction0_MCInst1_MC1_n145) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U16 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n111), .B(
        LED_RoundFunction0_MCInst1_MC1_n123), .ZN(
        LED_RoundFunction0_Feedback_59_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U15 ( .A(SubCellOutput0[57]), .B(
        SubCellOutput0[39]), .ZN(LED_RoundFunction0_MCInst1_MC1_n123) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U14 ( .A(SubCellOutput0[18]), .B(
        SubCellOutput0[14]), .Z(LED_RoundFunction0_MCInst1_MC1_n111) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U13 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n120), .B(
        LED_RoundFunction0_MCInst1_MC1_n121), .Z(
        LED_RoundFunction0_Feedback_58_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U12 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n147), .B(SubCellOutput0[56]), .Z(
        LED_RoundFunction0_MCInst1_MC1_n121) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U11 ( .A(SubCellOutput0[13]), .B(
        SubCellOutput0[59]), .Z(LED_RoundFunction0_MCInst1_MC1_n147) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U10 ( .A(SubCellOutput0[38]), .B(
        SubCellOutput0[17]), .Z(LED_RoundFunction0_MCInst1_MC1_n120) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U9 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n117), .B(
        LED_RoundFunction0_MCInst1_MC1_n109), .ZN(
        LED_RoundFunction0_Feedback_57_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U8 ( .A(SubCellOutput0[58]), .B(
        LED_RoundFunction0_MCInst1_MC1_n133), .Z(
        LED_RoundFunction0_MCInst1_MC1_n109) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U7 ( .A(SubCellOutput0[15]), .B(
        SubCellOutput0[59]), .Z(LED_RoundFunction0_MCInst1_MC1_n133) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U6 ( .A(
        LED_RoundFunction0_MCInst1_MC1_n159), .B(
        LED_RoundFunction0_MCInst1_MC1_n125), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n117) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U5 ( .A(SubCellOutput0[19]), .B(
        SubCellOutput0[37]), .Z(LED_RoundFunction0_MCInst1_MC1_n125) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U4 ( .A(SubCellOutput0[12]), .B(
        SubCellOutput0[16]), .Z(LED_RoundFunction0_MCInst1_MC1_n159) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U3 ( .A(SubCellOutput0[15]), .B(
        LED_RoundFunction0_MCInst1_MC1_n114), .ZN(
        LED_RoundFunction0_Feedback_56_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC1_U2 ( .A(SubCellOutput0[19]), .B(
        LED_RoundFunction0_MCInst1_MC1_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC1_n114) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC1_U1 ( .A(SubCellOutput0[58]), .B(
        SubCellOutput0[36]), .Z(LED_RoundFunction0_MCInst1_MC1_n126) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U68 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n160), .B(
        LED_RoundFunction0_MCInst1_MC2_n159), .ZN(
        LED_RoundFunction0_Feedback_7_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U67 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n158), .B(SubCellOutput0[54]), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n160) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U66 ( .A(SubCellOutput0[11]), .B(
        LED_RoundFunction0_MCInst1_MC2_n157), .Z(
        LED_RoundFunction0_Feedback_6_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U65 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n156), .B(
        LED_RoundFunction0_MCInst1_MC2_n155), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n157) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U64 ( .A(SubCellOutput0[29]), .B(
        SubCellOutput0[9]), .ZN(LED_RoundFunction0_MCInst1_MC2_n155) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U63 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n154), .B(SubCellOutput0[33]), .Z(
        LED_RoundFunction0_MCInst1_MC2_n156) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U62 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n153), .B(
        LED_RoundFunction0_MCInst1_MC2_n152), .ZN(
        LED_RoundFunction0_Feedback_5_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U61 ( .A(SubCellOutput0[10]), .B(
        SubCellOutput0[32]), .ZN(LED_RoundFunction0_MCInst1_MC2_n152) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U60 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n151), .B(
        LED_RoundFunction0_MCInst1_MC2_n150), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n153) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U59 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n149), .B(
        LED_RoundFunction0_MCInst1_MC2_n148), .ZN(
        LED_RoundFunction0_Feedback_4_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U58 ( .A(SubCellOutput0[31]), .B(
        LED_RoundFunction0_MCInst1_MC2_n147), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n148) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U57 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n146), .B(
        LED_RoundFunction0_MCInst1_MC2_n150), .Z(
        LED_RoundFunction0_MCInst1_MC2_n149) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U56 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n145), .B(
        LED_RoundFunction0_MCInst1_MC2_n159), .Z(
        LED_RoundFunction0_MCInst1_MC2_n150) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC2_U55 ( .A1(SubCellOutput0[29]), .A2(
        SubCellOutput0[30]), .B1(LED_RoundFunction0_MCInst1_MC2_n144), .B2(
        LED_RoundFunction0_MCInst1_MC2_n143), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n146) );
  INV_X1 LED_RoundFunction0_MCInst1_MC2_U54 ( .A(SubCellOutput0[29]), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n143) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U53 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n142), .B(
        LED_RoundFunction0_MCInst1_MC2_n141), .ZN(
        LED_RoundFunction0_Feedback_23_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U52 ( .A(SubCellOutput0[35]), .B(
        LED_RoundFunction0_MCInst1_MC2_n140), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n141) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U51 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n139), .B(SubCellOutput0[52]), .Z(
        LED_RoundFunction0_MCInst1_MC2_n142) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC2_U50 ( .A1(SubCellOutput0[34]), .A2(
        SubCellOutput0[30]), .B1(LED_RoundFunction0_MCInst1_MC2_n144), .B2(
        LED_RoundFunction0_MCInst1_MC2_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n139) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U49 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n137), .B(
        LED_RoundFunction0_MCInst1_MC2_n136), .ZN(
        LED_RoundFunction0_Feedback_22_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U48 ( .A(SubCellOutput0[32]), .B(
        LED_RoundFunction0_MCInst1_MC2_n135), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n136) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U47 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n134), .B(
        LED_RoundFunction0_MCInst1_MC2_n133), .Z(
        LED_RoundFunction0_MCInst1_MC2_n137) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC2_U46 ( .A1(SubCellOutput0[30]), .A2(
        SubCellOutput0[53]), .B1(LED_RoundFunction0_MCInst1_MC2_n132), .B2(
        LED_RoundFunction0_MCInst1_MC2_n144), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n134) );
  INV_X1 LED_RoundFunction0_MCInst1_MC2_U45 ( .A(SubCellOutput0[30]), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n144) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U44 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n131), .B(
        LED_RoundFunction0_MCInst1_MC2_n151), .ZN(
        LED_RoundFunction0_Feedback_21_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U43 ( .A(SubCellOutput0[55]), .B(
        SubCellOutput0[52]), .ZN(LED_RoundFunction0_MCInst1_MC2_n151) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U42 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n130), .B(
        LED_RoundFunction0_MCInst1_MC2_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n131) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U41 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n128), .B(
        LED_RoundFunction0_MCInst1_MC2_n127), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n130) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U40 ( .A(SubCellOutput0[29]), .B(
        LED_RoundFunction0_MCInst1_MC2_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n127) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U39 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n125), .B(SubCellOutput0[28]), .Z(
        LED_RoundFunction0_MCInst1_MC2_n128) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U38 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n124), .B(
        LED_RoundFunction0_MCInst1_MC2_n123), .ZN(
        LED_RoundFunction0_Feedback_20_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U37 ( .A(SubCellOutput0[8]), .B(
        LED_RoundFunction0_MCInst1_MC2_n122), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n124) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U36 ( .A(SubCellOutput0[10]), .B(
        LED_RoundFunction0_MCInst1_MC2_n122), .ZN(
        LED_RoundFunction0_Feedback_39_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U35 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n135), .B(
        LED_RoundFunction0_MCInst1_MC2_n121), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n122) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U34 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n120), .B(
        LED_RoundFunction0_MCInst1_MC2_n125), .Z(
        LED_RoundFunction0_MCInst1_MC2_n135) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U33 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n119), .B(
        LED_RoundFunction0_MCInst1_MC2_n118), .ZN(
        LED_RoundFunction0_Feedback_38_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U32 ( .A(SubCellOutput0[30]), .B(
        LED_RoundFunction0_MCInst1_MC2_n145), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n118) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U31 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n140), .B(
        LED_RoundFunction0_MCInst1_MC2_n147), .Z(
        LED_RoundFunction0_MCInst1_MC2_n119) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U30 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n126), .B(
        LED_RoundFunction0_MCInst1_MC2_n117), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n140) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U29 ( .A(SubCellOutput0[8]), .B(
        LED_RoundFunction0_MCInst1_MC2_n116), .ZN(
        LED_RoundFunction0_Feedback_37_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U28 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n115), .B(
        LED_RoundFunction0_MCInst1_MC2_n114), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n116) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U27 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n158), .B(SubCellOutput0[53]), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n115) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U26 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n120), .B(
        LED_RoundFunction0_MCInst1_MC2_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n158) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U25 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n113), .B(
        LED_RoundFunction0_MCInst1_MC2_n112), .ZN(
        LED_RoundFunction0_Feedback_36_) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC2_U24 ( .A1(SubCellOutput0[34]), .A2(
        LED_RoundFunction0_MCInst1_MC2_n111), .B1(
        LED_RoundFunction0_MCInst1_MC2_n129), .B2(
        LED_RoundFunction0_MCInst1_MC2_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n112) );
  INV_X1 LED_RoundFunction0_MCInst1_MC2_U23 ( .A(SubCellOutput0[34]), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n138) );
  INV_X1 LED_RoundFunction0_MCInst1_MC2_U22 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n111), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n129) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U21 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n145), .B(
        LED_RoundFunction0_MCInst1_MC2_n154), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n113) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC2_U20 ( .A1(SubCellOutput0[53]), .A2(
        SubCellOutput0[28]), .B1(LED_RoundFunction0_MCInst1_MC2_n110), .B2(
        LED_RoundFunction0_MCInst1_MC2_n132), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n154) );
  INV_X1 LED_RoundFunction0_MCInst1_MC2_U19 ( .A(SubCellOutput0[53]), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n132) );
  INV_X1 LED_RoundFunction0_MCInst1_MC2_U18 ( .A(SubCellOutput0[28]), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n110) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U17 ( .A(SubCellOutput0[11]), .B(
        SubCellOutput0[35]), .Z(LED_RoundFunction0_MCInst1_MC2_n145) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U16 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n111), .B(
        LED_RoundFunction0_MCInst1_MC2_n123), .ZN(
        LED_RoundFunction0_Feedback_55_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U15 ( .A(SubCellOutput0[53]), .B(
        SubCellOutput0[35]), .ZN(LED_RoundFunction0_MCInst1_MC2_n123) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U14 ( .A(SubCellOutput0[30]), .B(
        SubCellOutput0[10]), .Z(LED_RoundFunction0_MCInst1_MC2_n111) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U13 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n120), .B(
        LED_RoundFunction0_MCInst1_MC2_n121), .Z(
        LED_RoundFunction0_Feedback_54_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U12 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n147), .B(SubCellOutput0[52]), .Z(
        LED_RoundFunction0_MCInst1_MC2_n121) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U11 ( .A(SubCellOutput0[9]), .B(
        SubCellOutput0[55]), .Z(LED_RoundFunction0_MCInst1_MC2_n147) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U10 ( .A(SubCellOutput0[34]), .B(
        SubCellOutput0[29]), .Z(LED_RoundFunction0_MCInst1_MC2_n120) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U9 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n117), .B(
        LED_RoundFunction0_MCInst1_MC2_n109), .ZN(
        LED_RoundFunction0_Feedback_53_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U8 ( .A(SubCellOutput0[54]), .B(
        LED_RoundFunction0_MCInst1_MC2_n133), .Z(
        LED_RoundFunction0_MCInst1_MC2_n109) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U7 ( .A(SubCellOutput0[11]), .B(
        SubCellOutput0[55]), .Z(LED_RoundFunction0_MCInst1_MC2_n133) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U6 ( .A(
        LED_RoundFunction0_MCInst1_MC2_n159), .B(
        LED_RoundFunction0_MCInst1_MC2_n125), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n117) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U5 ( .A(SubCellOutput0[31]), .B(
        SubCellOutput0[33]), .Z(LED_RoundFunction0_MCInst1_MC2_n125) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U4 ( .A(SubCellOutput0[8]), .B(
        SubCellOutput0[28]), .Z(LED_RoundFunction0_MCInst1_MC2_n159) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U3 ( .A(SubCellOutput0[11]), .B(
        LED_RoundFunction0_MCInst1_MC2_n114), .ZN(
        LED_RoundFunction0_Feedback_52_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC2_U2 ( .A(SubCellOutput0[31]), .B(
        LED_RoundFunction0_MCInst1_MC2_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC2_n114) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC2_U1 ( .A(SubCellOutput0[54]), .B(
        SubCellOutput0[32]), .Z(LED_RoundFunction0_MCInst1_MC2_n126) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U68 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n160), .B(
        LED_RoundFunction0_MCInst1_MC3_n159), .ZN(
        LED_RoundFunction0_Feedback_3_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U67 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n158), .B(SubCellOutput0[50]), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n160) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U66 ( .A(SubCellOutput0[7]), .B(
        LED_RoundFunction0_MCInst1_MC3_n157), .Z(
        LED_RoundFunction0_Feedback_2_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U65 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n156), .B(
        LED_RoundFunction0_MCInst1_MC3_n155), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n157) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U64 ( .A(SubCellOutput0[25]), .B(
        SubCellOutput0[5]), .ZN(LED_RoundFunction0_MCInst1_MC3_n155) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U63 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n154), .B(SubCellOutput0[45]), .Z(
        LED_RoundFunction0_MCInst1_MC3_n156) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U62 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n153), .B(
        LED_RoundFunction0_MCInst1_MC3_n152), .ZN(
        LED_RoundFunction0_Feedback_1_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U61 ( .A(SubCellOutput0[6]), .B(
        SubCellOutput0[44]), .ZN(LED_RoundFunction0_MCInst1_MC3_n152) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U60 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n151), .B(
        LED_RoundFunction0_MCInst1_MC3_n150), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n153) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U59 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n149), .B(
        LED_RoundFunction0_MCInst1_MC3_n148), .ZN(
        LED_RoundFunction0_Feedback_0_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U58 ( .A(SubCellOutput0[27]), .B(
        LED_RoundFunction0_MCInst1_MC3_n147), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n148) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U57 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n146), .B(
        LED_RoundFunction0_MCInst1_MC3_n150), .Z(
        LED_RoundFunction0_MCInst1_MC3_n149) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U56 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n145), .B(
        LED_RoundFunction0_MCInst1_MC3_n159), .Z(
        LED_RoundFunction0_MCInst1_MC3_n150) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC3_U55 ( .A1(SubCellOutput0[25]), .A2(
        SubCellOutput0[26]), .B1(LED_RoundFunction0_MCInst1_MC3_n144), .B2(
        LED_RoundFunction0_MCInst1_MC3_n143), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n146) );
  INV_X1 LED_RoundFunction0_MCInst1_MC3_U54 ( .A(SubCellOutput0[25]), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n143) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U53 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n142), .B(
        LED_RoundFunction0_MCInst1_MC3_n141), .ZN(
        LED_RoundFunction0_Feedback_19_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U52 ( .A(SubCellOutput0[47]), .B(
        LED_RoundFunction0_MCInst1_MC3_n140), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n141) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U51 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n139), .B(SubCellOutput0[48]), .Z(
        LED_RoundFunction0_MCInst1_MC3_n142) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC3_U50 ( .A1(SubCellOutput0[46]), .A2(
        SubCellOutput0[26]), .B1(LED_RoundFunction0_MCInst1_MC3_n144), .B2(
        LED_RoundFunction0_MCInst1_MC3_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n139) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U49 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n137), .B(
        LED_RoundFunction0_MCInst1_MC3_n136), .ZN(
        LED_RoundFunction0_Feedback_18_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U48 ( .A(SubCellOutput0[44]), .B(
        LED_RoundFunction0_MCInst1_MC3_n135), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n136) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U47 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n134), .B(
        LED_RoundFunction0_MCInst1_MC3_n133), .Z(
        LED_RoundFunction0_MCInst1_MC3_n137) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC3_U46 ( .A1(SubCellOutput0[26]), .A2(
        SubCellOutput0[49]), .B1(LED_RoundFunction0_MCInst1_MC3_n132), .B2(
        LED_RoundFunction0_MCInst1_MC3_n144), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n134) );
  INV_X1 LED_RoundFunction0_MCInst1_MC3_U45 ( .A(SubCellOutput0[26]), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n144) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U44 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n131), .B(
        LED_RoundFunction0_MCInst1_MC3_n151), .ZN(
        LED_RoundFunction0_Feedback_17_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U43 ( .A(SubCellOutput0[51]), .B(
        SubCellOutput0[48]), .ZN(LED_RoundFunction0_MCInst1_MC3_n151) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U42 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n130), .B(
        LED_RoundFunction0_MCInst1_MC3_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n131) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U41 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n128), .B(
        LED_RoundFunction0_MCInst1_MC3_n127), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n130) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U40 ( .A(SubCellOutput0[25]), .B(
        LED_RoundFunction0_MCInst1_MC3_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n127) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U39 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n125), .B(SubCellOutput0[24]), .Z(
        LED_RoundFunction0_MCInst1_MC3_n128) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U38 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n124), .B(
        LED_RoundFunction0_MCInst1_MC3_n123), .ZN(
        LED_RoundFunction0_Feedback_16_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U37 ( .A(SubCellOutput0[4]), .B(
        LED_RoundFunction0_MCInst1_MC3_n122), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n124) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U36 ( .A(SubCellOutput0[6]), .B(
        LED_RoundFunction0_MCInst1_MC3_n122), .ZN(
        LED_RoundFunction0_Feedback_35_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U35 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n135), .B(
        LED_RoundFunction0_MCInst1_MC3_n121), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n122) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U34 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n120), .B(
        LED_RoundFunction0_MCInst1_MC3_n125), .Z(
        LED_RoundFunction0_MCInst1_MC3_n135) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U33 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n119), .B(
        LED_RoundFunction0_MCInst1_MC3_n118), .ZN(
        LED_RoundFunction0_Feedback_34_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U32 ( .A(SubCellOutput0[26]), .B(
        LED_RoundFunction0_MCInst1_MC3_n145), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n118) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U31 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n140), .B(
        LED_RoundFunction0_MCInst1_MC3_n147), .Z(
        LED_RoundFunction0_MCInst1_MC3_n119) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U30 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n126), .B(
        LED_RoundFunction0_MCInst1_MC3_n117), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n140) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U29 ( .A(SubCellOutput0[4]), .B(
        LED_RoundFunction0_MCInst1_MC3_n116), .ZN(
        LED_RoundFunction0_Feedback_33_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U28 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n115), .B(
        LED_RoundFunction0_MCInst1_MC3_n114), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n116) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U27 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n158), .B(SubCellOutput0[49]), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n115) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U26 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n120), .B(
        LED_RoundFunction0_MCInst1_MC3_n129), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n158) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U25 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n113), .B(
        LED_RoundFunction0_MCInst1_MC3_n112), .ZN(
        LED_RoundFunction0_Feedback_32_) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC3_U24 ( .A1(SubCellOutput0[46]), .A2(
        LED_RoundFunction0_MCInst1_MC3_n111), .B1(
        LED_RoundFunction0_MCInst1_MC3_n129), .B2(
        LED_RoundFunction0_MCInst1_MC3_n138), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n112) );
  INV_X1 LED_RoundFunction0_MCInst1_MC3_U23 ( .A(SubCellOutput0[46]), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n138) );
  INV_X1 LED_RoundFunction0_MCInst1_MC3_U22 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n111), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n129) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U21 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n145), .B(
        LED_RoundFunction0_MCInst1_MC3_n154), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n113) );
  AOI22_X1 LED_RoundFunction0_MCInst1_MC3_U20 ( .A1(SubCellOutput0[49]), .A2(
        SubCellOutput0[24]), .B1(LED_RoundFunction0_MCInst1_MC3_n110), .B2(
        LED_RoundFunction0_MCInst1_MC3_n132), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n154) );
  INV_X1 LED_RoundFunction0_MCInst1_MC3_U19 ( .A(SubCellOutput0[49]), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n132) );
  INV_X1 LED_RoundFunction0_MCInst1_MC3_U18 ( .A(SubCellOutput0[24]), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n110) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U17 ( .A(SubCellOutput0[7]), .B(
        SubCellOutput0[47]), .Z(LED_RoundFunction0_MCInst1_MC3_n145) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U16 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n111), .B(
        LED_RoundFunction0_MCInst1_MC3_n123), .ZN(
        LED_RoundFunction0_Feedback_51_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U15 ( .A(SubCellOutput0[49]), .B(
        SubCellOutput0[47]), .ZN(LED_RoundFunction0_MCInst1_MC3_n123) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U14 ( .A(SubCellOutput0[26]), .B(
        SubCellOutput0[6]), .Z(LED_RoundFunction0_MCInst1_MC3_n111) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U13 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n120), .B(
        LED_RoundFunction0_MCInst1_MC3_n121), .Z(
        LED_RoundFunction0_Feedback_50_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U12 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n147), .B(SubCellOutput0[48]), .Z(
        LED_RoundFunction0_MCInst1_MC3_n121) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U11 ( .A(SubCellOutput0[5]), .B(
        SubCellOutput0[51]), .Z(LED_RoundFunction0_MCInst1_MC3_n147) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U10 ( .A(SubCellOutput0[46]), .B(
        SubCellOutput0[25]), .Z(LED_RoundFunction0_MCInst1_MC3_n120) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U9 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n117), .B(
        LED_RoundFunction0_MCInst1_MC3_n109), .ZN(
        LED_RoundFunction0_Feedback_49_) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U8 ( .A(SubCellOutput0[50]), .B(
        LED_RoundFunction0_MCInst1_MC3_n133), .Z(
        LED_RoundFunction0_MCInst1_MC3_n109) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U7 ( .A(SubCellOutput0[7]), .B(
        SubCellOutput0[51]), .Z(LED_RoundFunction0_MCInst1_MC3_n133) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U6 ( .A(
        LED_RoundFunction0_MCInst1_MC3_n159), .B(
        LED_RoundFunction0_MCInst1_MC3_n125), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n117) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U5 ( .A(SubCellOutput0[27]), .B(
        SubCellOutput0[45]), .Z(LED_RoundFunction0_MCInst1_MC3_n125) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U4 ( .A(SubCellOutput0[4]), .B(
        SubCellOutput0[24]), .Z(LED_RoundFunction0_MCInst1_MC3_n159) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U3 ( .A(SubCellOutput0[7]), .B(
        LED_RoundFunction0_MCInst1_MC3_n114), .ZN(
        LED_RoundFunction0_Feedback_48_) );
  XNOR2_X1 LED_RoundFunction0_MCInst1_MC3_U2 ( .A(SubCellOutput0[27]), .B(
        LED_RoundFunction0_MCInst1_MC3_n126), .ZN(
        LED_RoundFunction0_MCInst1_MC3_n114) );
  XOR2_X1 LED_RoundFunction0_MCInst1_MC3_U1 ( .A(SubCellOutput0[50]), .B(
        SubCellOutput0[44]), .Z(LED_RoundFunction0_MCInst1_MC3_n126) );
  AOI22_X1 LED_RoundFunction1_U412 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n836), .B1(LED_RoundFunction1_n835), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U411 ( .A1(rst), .A2(Plaintext1[0]), .B1(
        LED_RoundFunction1_Feedback_0_), .B2(LED_RoundFunction1_n564), .ZN(
        LED_RoundFunction1_n835) );
  INV_X1 LED_RoundFunction1_U410 ( .A(Ciphertext1[0]), .ZN(
        LED_RoundFunction1_n836) );
  AOI22_X1 LED_RoundFunction1_U409 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n834), .B1(LED_RoundFunction1_n833), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U408 ( .A1(rst), .A2(Plaintext1[1]), .B1(
        LED_RoundFunction1_Feedback_1_), .B2(LED_RoundFunction1_n568), .ZN(
        LED_RoundFunction1_n833) );
  INV_X1 LED_RoundFunction1_U407 ( .A(Ciphertext1[1]), .ZN(
        LED_RoundFunction1_n834) );
  AOI22_X1 LED_RoundFunction1_U406 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n832), .B1(LED_RoundFunction1_n831), .B2(
        LED_RoundFunction1_n561), .ZN(SubCellInput1[2]) );
  AOI22_X1 LED_RoundFunction1_U405 ( .A1(rst), .A2(Plaintext1[2]), .B1(
        LED_RoundFunction1_Feedback_2_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n831) );
  INV_X1 LED_RoundFunction1_U404 ( .A(Ciphertext1[2]), .ZN(
        LED_RoundFunction1_n832) );
  AOI22_X1 LED_RoundFunction1_U403 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n830), .B1(LED_RoundFunction1_n829), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U402 ( .A1(rst), .A2(Plaintext1[3]), .B1(
        LED_RoundFunction1_Feedback_3_), .B2(LED_RoundFunction1_n568), .ZN(
        LED_RoundFunction1_n829) );
  INV_X1 LED_RoundFunction1_U401 ( .A(Ciphertext1[3]), .ZN(
        LED_RoundFunction1_n830) );
  AOI22_X1 LED_RoundFunction1_U400 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n828), .B1(LED_RoundFunction1_n827), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U399 ( .A1(rst), .A2(Plaintext1[4]), .B1(
        LED_RoundFunction1_Feedback_4_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n827) );
  INV_X1 LED_RoundFunction1_U398 ( .A(Ciphertext1[4]), .ZN(
        LED_RoundFunction1_n828) );
  AOI22_X1 LED_RoundFunction1_U397 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n826), .B1(LED_RoundFunction1_n825), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U396 ( .A1(rst), .A2(Plaintext1[5]), .B1(
        LED_RoundFunction1_Feedback_5_), .B2(LED_RoundFunction1_n568), .ZN(
        LED_RoundFunction1_n825) );
  INV_X1 LED_RoundFunction1_U395 ( .A(Ciphertext1[5]), .ZN(
        LED_RoundFunction1_n826) );
  AOI22_X1 LED_RoundFunction1_U394 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n824), .B1(LED_RoundFunction1_n823), .B2(
        LED_RoundFunction1_n560), .ZN(SubCellInput1[6]) );
  AOI22_X1 LED_RoundFunction1_U393 ( .A1(rst), .A2(Plaintext1[6]), .B1(
        LED_RoundFunction1_Feedback_6_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n823) );
  INV_X1 LED_RoundFunction1_U392 ( .A(Ciphertext1[6]), .ZN(
        LED_RoundFunction1_n824) );
  AOI22_X1 LED_RoundFunction1_U391 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n822), .B1(LED_RoundFunction1_n821), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U390 ( .A1(rst), .A2(Plaintext1[7]), .B1(
        LED_RoundFunction1_Feedback_7_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n821) );
  INV_X1 LED_RoundFunction1_U389 ( .A(Ciphertext1[7]), .ZN(
        LED_RoundFunction1_n822) );
  AOI22_X1 LED_RoundFunction1_U388 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n820), .B1(LED_RoundFunction1_n819), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U387 ( .A1(rst), .A2(Plaintext1[11]), .B1(
        LED_RoundFunction1_Feedback_11_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n819) );
  INV_X1 LED_RoundFunction1_U386 ( .A(Ciphertext1[11]), .ZN(
        LED_RoundFunction1_n820) );
  AOI22_X1 LED_RoundFunction1_U385 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n818), .B1(LED_RoundFunction1_n817), .B2(
        LED_RoundFunction1_n561), .ZN(SubCellInput1[14]) );
  AOI22_X1 LED_RoundFunction1_U384 ( .A1(rst), .A2(Plaintext1[14]), .B1(
        LED_RoundFunction1_Feedback_14_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n817) );
  INV_X1 LED_RoundFunction1_U383 ( .A(Ciphertext1[14]), .ZN(
        LED_RoundFunction1_n818) );
  AOI22_X1 LED_RoundFunction1_U382 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n816), .B1(LED_RoundFunction1_n815), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U381 ( .A1(rst), .A2(Plaintext1[15]), .B1(
        LED_RoundFunction1_Feedback_15_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n815) );
  INV_X1 LED_RoundFunction1_U380 ( .A(Ciphertext1[15]), .ZN(
        LED_RoundFunction1_n816) );
  AOI22_X1 LED_RoundFunction1_U379 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n814), .B1(LED_RoundFunction1_n813), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U378 ( .A1(rst), .A2(Plaintext1[16]), .B1(
        LED_RoundFunction1_Feedback_16_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n813) );
  INV_X1 LED_RoundFunction1_U377 ( .A(Ciphertext1[16]), .ZN(
        LED_RoundFunction1_n814) );
  AOI22_X1 LED_RoundFunction1_U376 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n812), .B1(LED_RoundFunction1_n811), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U375 ( .A1(rst), .A2(Plaintext1[17]), .B1(
        LED_RoundFunction1_Feedback_17_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n811) );
  INV_X1 LED_RoundFunction1_U374 ( .A(Ciphertext1[17]), .ZN(
        LED_RoundFunction1_n812) );
  AOI22_X1 LED_RoundFunction1_U373 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n810), .B1(LED_RoundFunction1_n809), .B2(
        LED_RoundFunction1_n560), .ZN(SubCellInput1[18]) );
  AOI22_X1 LED_RoundFunction1_U372 ( .A1(rst), .A2(Plaintext1[18]), .B1(
        LED_RoundFunction1_Feedback_18_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n809) );
  INV_X1 LED_RoundFunction1_U371 ( .A(Ciphertext1[18]), .ZN(
        LED_RoundFunction1_n810) );
  AOI22_X1 LED_RoundFunction1_U370 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n808), .B1(LED_RoundFunction1_n807), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U369 ( .A1(rst), .A2(Plaintext1[19]), .B1(
        LED_RoundFunction1_Feedback_19_), .B2(LED_RoundFunction1_n568), .ZN(
        LED_RoundFunction1_n807) );
  INV_X1 LED_RoundFunction1_U368 ( .A(Ciphertext1[19]), .ZN(
        LED_RoundFunction1_n808) );
  AOI22_X1 LED_RoundFunction1_U367 ( .A1(LED_RoundFunction1_n557), .A2(
        LED_RoundFunction1_n806), .B1(LED_RoundFunction1_n805), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U366 ( .A1(rst), .A2(Plaintext1[20]), .B1(
        LED_RoundFunction1_Feedback_20_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n805) );
  INV_X1 LED_RoundFunction1_U365 ( .A(Ciphertext1[20]), .ZN(
        LED_RoundFunction1_n806) );
  AOI22_X1 LED_RoundFunction1_U364 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n804), .B1(LED_RoundFunction1_n803), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U363 ( .A1(rst), .A2(Plaintext1[21]), .B1(
        LED_RoundFunction1_Feedback_21_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n803) );
  INV_X1 LED_RoundFunction1_U362 ( .A(Ciphertext1[21]), .ZN(
        LED_RoundFunction1_n804) );
  AOI22_X1 LED_RoundFunction1_U361 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n802), .B1(LED_RoundFunction1_n801), .B2(
        LED_RoundFunction1_n561), .ZN(SubCellInput1[22]) );
  AOI22_X1 LED_RoundFunction1_U360 ( .A1(rst), .A2(Plaintext1[22]), .B1(
        LED_RoundFunction1_Feedback_22_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n801) );
  INV_X1 LED_RoundFunction1_U359 ( .A(Ciphertext1[22]), .ZN(
        LED_RoundFunction1_n802) );
  AOI22_X1 LED_RoundFunction1_U358 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n800), .B1(LED_RoundFunction1_n799), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U357 ( .A1(rst), .A2(Plaintext1[23]), .B1(
        LED_RoundFunction1_Feedback_23_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n799) );
  INV_X1 LED_RoundFunction1_U356 ( .A(Ciphertext1[23]), .ZN(
        LED_RoundFunction1_n800) );
  AOI22_X1 LED_RoundFunction1_U355 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n798), .B1(LED_RoundFunction1_n797), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U354 ( .A1(rst), .A2(Plaintext1[27]), .B1(
        LED_RoundFunction1_Feedback_27_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n797) );
  INV_X1 LED_RoundFunction1_U353 ( .A(Ciphertext1[27]), .ZN(
        LED_RoundFunction1_n798) );
  AOI22_X1 LED_RoundFunction1_U352 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n796), .B1(LED_RoundFunction1_n795), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U351 ( .A1(rst), .A2(Plaintext1[28]), .B1(
        LED_RoundFunction1_Feedback_28_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n795) );
  INV_X1 LED_RoundFunction1_U350 ( .A(Ciphertext1[28]), .ZN(
        LED_RoundFunction1_n796) );
  AOI22_X1 LED_RoundFunction1_U349 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n794), .B1(LED_RoundFunction1_n793), .B2(
        LED_RoundFunction1_n560), .ZN(SubCellInput1[30]) );
  AOI22_X1 LED_RoundFunction1_U348 ( .A1(rst), .A2(Plaintext1[30]), .B1(
        LED_RoundFunction1_Feedback_30_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n793) );
  INV_X1 LED_RoundFunction1_U347 ( .A(Ciphertext1[30]), .ZN(
        LED_RoundFunction1_n794) );
  AOI22_X1 LED_RoundFunction1_U346 ( .A1(LED_RoundFunction1_n556), .A2(
        LED_RoundFunction1_n792), .B1(LED_RoundFunction1_n791), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U345 ( .A1(rst), .A2(Plaintext1[31]), .B1(
        LED_RoundFunction1_Feedback_31_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n791) );
  INV_X1 LED_RoundFunction1_U344 ( .A(Ciphertext1[31]), .ZN(
        LED_RoundFunction1_n792) );
  AOI22_X1 LED_RoundFunction1_U343 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n790), .B1(LED_RoundFunction1_n789), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U342 ( .A1(rst), .A2(Plaintext1[32]), .B1(
        LED_RoundFunction1_Feedback_32_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n789) );
  INV_X1 LED_RoundFunction1_U341 ( .A(Ciphertext1[32]), .ZN(
        LED_RoundFunction1_n790) );
  AOI22_X1 LED_RoundFunction1_U340 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n788), .B1(LED_RoundFunction1_n787), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U339 ( .A1(rst), .A2(Plaintext1[33]), .B1(
        LED_RoundFunction1_Feedback_33_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n787) );
  INV_X1 LED_RoundFunction1_U338 ( .A(Ciphertext1[33]), .ZN(
        LED_RoundFunction1_n788) );
  AOI22_X1 LED_RoundFunction1_U337 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n786), .B1(LED_RoundFunction1_n785), .B2(
        LED_RoundFunction1_n561), .ZN(SubCellInput1[34]) );
  AOI22_X1 LED_RoundFunction1_U336 ( .A1(rst), .A2(Plaintext1[34]), .B1(
        LED_RoundFunction1_Feedback_34_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n785) );
  INV_X1 LED_RoundFunction1_U335 ( .A(Ciphertext1[34]), .ZN(
        LED_RoundFunction1_n786) );
  AOI22_X1 LED_RoundFunction1_U334 ( .A1(LED_RoundFunction1_n557), .A2(
        LED_RoundFunction1_n784), .B1(LED_RoundFunction1_n783), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U333 ( .A1(rst), .A2(Plaintext1[35]), .B1(
        LED_RoundFunction1_Feedback_35_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n783) );
  INV_X1 LED_RoundFunction1_U332 ( .A(Ciphertext1[35]), .ZN(
        LED_RoundFunction1_n784) );
  AOI22_X1 LED_RoundFunction1_U331 ( .A1(LED_RoundFunction1_n556), .A2(
        LED_RoundFunction1_n782), .B1(LED_RoundFunction1_n781), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U330 ( .A1(rst), .A2(Plaintext1[36]), .B1(
        LED_RoundFunction1_Feedback_36_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n781) );
  INV_X1 LED_RoundFunction1_U329 ( .A(Ciphertext1[36]), .ZN(
        LED_RoundFunction1_n782) );
  AOI22_X1 LED_RoundFunction1_U328 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n780), .B1(LED_RoundFunction1_n779), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U327 ( .A1(rst), .A2(Plaintext1[37]), .B1(
        LED_RoundFunction1_Feedback_37_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n779) );
  INV_X1 LED_RoundFunction1_U326 ( .A(Ciphertext1[37]), .ZN(
        LED_RoundFunction1_n780) );
  AOI22_X1 LED_RoundFunction1_U325 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n778), .B1(LED_RoundFunction1_n777), .B2(
        LED_RoundFunction1_n561), .ZN(SubCellInput1[38]) );
  AOI22_X1 LED_RoundFunction1_U324 ( .A1(rst), .A2(Plaintext1[38]), .B1(
        LED_RoundFunction1_Feedback_38_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n777) );
  INV_X1 LED_RoundFunction1_U323 ( .A(Ciphertext1[38]), .ZN(
        LED_RoundFunction1_n778) );
  AOI22_X1 LED_RoundFunction1_U322 ( .A1(LED_RoundFunction1_n556), .A2(
        LED_RoundFunction1_n776), .B1(LED_RoundFunction1_n775), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U321 ( .A1(rst), .A2(Plaintext1[39]), .B1(
        LED_RoundFunction1_Feedback_39_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n775) );
  INV_X1 LED_RoundFunction1_U320 ( .A(Ciphertext1[39]), .ZN(
        LED_RoundFunction1_n776) );
  AOI22_X1 LED_RoundFunction1_U319 ( .A1(LED_RoundFunction1_n557), .A2(
        LED_RoundFunction1_n774), .B1(LED_RoundFunction1_n773), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U318 ( .A1(rst), .A2(Plaintext1[43]), .B1(
        LED_RoundFunction1_Feedback_43_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n773) );
  INV_X1 LED_RoundFunction1_U317 ( .A(Ciphertext1[43]), .ZN(
        LED_RoundFunction1_n774) );
  AOI22_X1 LED_RoundFunction1_U316 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n772), .B1(LED_RoundFunction1_n771), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U315 ( .A1(rst), .A2(Plaintext1[45]), .B1(
        LED_RoundFunction1_Feedback_45_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n771) );
  INV_X1 LED_RoundFunction1_U314 ( .A(Ciphertext1[45]), .ZN(
        LED_RoundFunction1_n772) );
  AOI22_X1 LED_RoundFunction1_U313 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n770), .B1(LED_RoundFunction1_n769), .B2(
        LED_RoundFunction1_n561), .ZN(SubCellInput1[46]) );
  AOI22_X1 LED_RoundFunction1_U312 ( .A1(rst), .A2(Plaintext1[46]), .B1(
        LED_RoundFunction1_Feedback_46_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n769) );
  INV_X1 LED_RoundFunction1_U311 ( .A(Ciphertext1[46]), .ZN(
        LED_RoundFunction1_n770) );
  AOI22_X1 LED_RoundFunction1_U310 ( .A1(LED_RoundFunction1_n557), .A2(
        LED_RoundFunction1_n768), .B1(LED_RoundFunction1_n767), .B2(
        LED_RoundFunction1_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U309 ( .A1(rst), .A2(Plaintext1[48]), .B1(
        LED_RoundFunction1_Feedback_48_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n767) );
  INV_X1 LED_RoundFunction1_U308 ( .A(Ciphertext1[48]), .ZN(
        LED_RoundFunction1_n768) );
  AOI22_X1 LED_RoundFunction1_U307 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n766), .B1(LED_RoundFunction1_n765), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U306 ( .A1(rst), .A2(Plaintext1[49]), .B1(
        LED_RoundFunction1_Feedback_49_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n765) );
  INV_X1 LED_RoundFunction1_U305 ( .A(Ciphertext1[49]), .ZN(
        LED_RoundFunction1_n766) );
  AOI22_X1 LED_RoundFunction1_U304 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n764), .B1(LED_RoundFunction1_n763), .B2(
        LED_RoundFunction1_n560), .ZN(SubCellInput1[50]) );
  AOI22_X1 LED_RoundFunction1_U303 ( .A1(rst), .A2(Plaintext1[50]), .B1(
        LED_RoundFunction1_Feedback_50_), .B2(LED_RoundFunction1_n562), .ZN(
        LED_RoundFunction1_n763) );
  INV_X1 LED_RoundFunction1_U302 ( .A(Ciphertext1[50]), .ZN(
        LED_RoundFunction1_n764) );
  AOI22_X1 LED_RoundFunction1_U301 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n762), .B1(LED_RoundFunction1_n761), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U300 ( .A1(rst), .A2(Plaintext1[51]), .B1(
        LED_RoundFunction1_Feedback_51_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n761) );
  INV_X1 LED_RoundFunction1_U299 ( .A(Ciphertext1[51]), .ZN(
        LED_RoundFunction1_n762) );
  AOI22_X1 LED_RoundFunction1_U298 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n760), .B1(LED_RoundFunction1_n759), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U297 ( .A1(rst), .A2(Plaintext1[52]), .B1(
        LED_RoundFunction1_Feedback_52_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n759) );
  INV_X1 LED_RoundFunction1_U296 ( .A(Ciphertext1[52]), .ZN(
        LED_RoundFunction1_n760) );
  AOI22_X1 LED_RoundFunction1_U295 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n758), .B1(LED_RoundFunction1_n757), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U294 ( .A1(rst), .A2(Plaintext1[53]), .B1(
        LED_RoundFunction1_Feedback_53_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n757) );
  INV_X1 LED_RoundFunction1_U293 ( .A(Ciphertext1[53]), .ZN(
        LED_RoundFunction1_n758) );
  AOI22_X1 LED_RoundFunction1_U292 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n756), .B1(LED_RoundFunction1_n755), .B2(
        LED_RoundFunction1_n560), .ZN(SubCellInput1[54]) );
  AOI22_X1 LED_RoundFunction1_U291 ( .A1(rst), .A2(Plaintext1[54]), .B1(
        LED_RoundFunction1_Feedback_54_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n755) );
  INV_X1 LED_RoundFunction1_U290 ( .A(Ciphertext1[54]), .ZN(
        LED_RoundFunction1_n756) );
  AOI22_X1 LED_RoundFunction1_U289 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n754), .B1(LED_RoundFunction1_n753), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U288 ( .A1(rst), .A2(Plaintext1[55]), .B1(
        LED_RoundFunction1_Feedback_55_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n753) );
  INV_X1 LED_RoundFunction1_U287 ( .A(Ciphertext1[55]), .ZN(
        LED_RoundFunction1_n754) );
  AOI22_X1 LED_RoundFunction1_U286 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n752), .B1(LED_RoundFunction1_n751), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[1]) );
  AOI22_X1 LED_RoundFunction1_U285 ( .A1(rst), .A2(Plaintext1[59]), .B1(
        LED_RoundFunction1_Feedback_59_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n751) );
  INV_X1 LED_RoundFunction1_U284 ( .A(Ciphertext1[59]), .ZN(
        LED_RoundFunction1_n752) );
  AOI22_X1 LED_RoundFunction1_U283 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n750), .B1(LED_RoundFunction1_n749), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[0]) );
  AOI22_X1 LED_RoundFunction1_U282 ( .A1(rst), .A2(Plaintext1[60]), .B1(
        LED_RoundFunction1_Feedback_60_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n749) );
  INV_X1 LED_RoundFunction1_U281 ( .A(Ciphertext1[60]), .ZN(
        LED_RoundFunction1_n750) );
  AOI22_X1 LED_RoundFunction1_U280 ( .A1(LED_RoundFunction1_n558), .A2(
        LED_RoundFunction1_n748), .B1(LED_RoundFunction1_n747), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[2]) );
  AOI22_X1 LED_RoundFunction1_U279 ( .A1(rst), .A2(Plaintext1[61]), .B1(
        LED_RoundFunction1_Feedback_61_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n747) );
  INV_X1 LED_RoundFunction1_U278 ( .A(Ciphertext1[61]), .ZN(
        LED_RoundFunction1_n748) );
  AOI22_X1 LED_RoundFunction1_U277 ( .A1(LED_RoundFunction1_n555), .A2(
        LED_RoundFunction1_n746), .B1(LED_RoundFunction1_n745), .B2(
        LED_RoundFunction1_n560), .ZN(SubCellInput1[62]) );
  AOI22_X1 LED_RoundFunction1_U276 ( .A1(rst), .A2(Plaintext1[62]), .B1(
        LED_RoundFunction1_Feedback_62_), .B2(LED_RoundFunction1_n563), .ZN(
        LED_RoundFunction1_n745) );
  INV_X1 LED_RoundFunction1_U275 ( .A(Ciphertext1[62]), .ZN(
        LED_RoundFunction1_n746) );
  XOR2_X1 LED_RoundFunction1_U274 ( .A(1'b0), .B(LED_RoundFunction1_n744), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[2]) );
  AOI21_X1 LED_RoundFunction1_U273 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n743), .A(LED_RoundFunction1_n742), .ZN(
        LED_RoundFunction1_n744) );
  AOI221_X1 LED_RoundFunction1_U272 ( .B1(Plaintext1[9]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_9_), .C2(LED_RoundFunction1_n568), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n742) );
  INV_X1 LED_RoundFunction1_U271 ( .A(Ciphertext1[9]), .ZN(
        LED_RoundFunction1_n743) );
  XOR2_X1 LED_RoundFunction1_U270 ( .A(1'b0), .B(LED_RoundFunction1_n741), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[0]) );
  AOI21_X1 LED_RoundFunction1_U269 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n740), .A(LED_RoundFunction1_n739), .ZN(
        LED_RoundFunction1_n741) );
  AOI221_X1 LED_RoundFunction1_U268 ( .B1(Plaintext1[8]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_8_), .C2(LED_RoundFunction1_n566), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n739) );
  INV_X1 LED_RoundFunction1_U267 ( .A(Ciphertext1[8]), .ZN(
        LED_RoundFunction1_n740) );
  AOI22_X1 LED_RoundFunction1_U266 ( .A1(LED_RoundFunction1_n555), .A2(
        Ciphertext1[63]), .B1(LED_RoundFunction1_n738), .B2(
        LED_RoundFunction1_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[1]) );
  INV_X1 LED_RoundFunction1_U265 ( .A(LED_RoundFunction1_n737), .ZN(
        LED_RoundFunction1_n738) );
  OAI22_X1 LED_RoundFunction1_U264 ( .A1(LED_RoundFunction1_n565), .A2(
        Plaintext1[63]), .B1(LED_RoundFunction1_Feedback_63_), .B2(rst), .ZN(
        LED_RoundFunction1_n737) );
  XOR2_X1 LED_RoundFunction1_U263 ( .A(1'b0), .B(LED_RoundFunction1_n736), .Z(
        SubCellInput1[58]) );
  AOI21_X1 LED_RoundFunction1_U262 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n735), .A(LED_RoundFunction1_n734), .ZN(
        LED_RoundFunction1_n736) );
  AOI221_X1 LED_RoundFunction1_U261 ( .B1(Plaintext1[58]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_58_), .C2(LED_RoundFunction1_n565), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n734) );
  INV_X1 LED_RoundFunction1_U260 ( .A(Ciphertext1[58]), .ZN(
        LED_RoundFunction1_n735) );
  XOR2_X1 LED_RoundFunction1_U259 ( .A(1'b0), .B(LED_RoundFunction1_n733), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[2]) );
  AOI21_X1 LED_RoundFunction1_U258 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n732), .A(LED_RoundFunction1_n731), .ZN(
        LED_RoundFunction1_n733) );
  AOI221_X1 LED_RoundFunction1_U257 ( .B1(Plaintext1[57]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_57_), .C2(LED_RoundFunction1_n566), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n731) );
  INV_X1 LED_RoundFunction1_U256 ( .A(Ciphertext1[57]), .ZN(
        LED_RoundFunction1_n732) );
  XOR2_X1 LED_RoundFunction1_U255 ( .A(1'b0), .B(LED_RoundFunction1_n730), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[0]) );
  AOI21_X1 LED_RoundFunction1_U254 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n729), .A(LED_RoundFunction1_n728), .ZN(
        LED_RoundFunction1_n730) );
  AOI221_X1 LED_RoundFunction1_U253 ( .B1(Plaintext1[56]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_56_), .C2(LED_RoundFunction1_n568), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n728) );
  INV_X1 LED_RoundFunction1_U252 ( .A(Ciphertext1[56]), .ZN(
        LED_RoundFunction1_n729) );
  AOI22_X1 LED_RoundFunction1_U251 ( .A1(LED_RoundFunction1_n556), .A2(
        Ciphertext1[47]), .B1(LED_RoundFunction1_n727), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[1]) );
  INV_X1 LED_RoundFunction1_U250 ( .A(LED_RoundFunction1_n726), .ZN(
        LED_RoundFunction1_n727) );
  OAI22_X1 LED_RoundFunction1_U249 ( .A1(LED_RoundFunction1_n568), .A2(
        Plaintext1[47]), .B1(LED_RoundFunction1_Feedback_47_), .B2(rst), .ZN(
        LED_RoundFunction1_n726) );
  AOI22_X1 LED_RoundFunction1_U248 ( .A1(LED_RoundFunction1_n556), .A2(
        Ciphertext1[44]), .B1(LED_RoundFunction1_n725), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[0]) );
  INV_X1 LED_RoundFunction1_U247 ( .A(LED_RoundFunction1_n724), .ZN(
        LED_RoundFunction1_n725) );
  OAI22_X1 LED_RoundFunction1_U246 ( .A1(LED_RoundFunction1_n568), .A2(
        Plaintext1[44]), .B1(LED_RoundFunction1_Feedback_44_), .B2(rst), .ZN(
        LED_RoundFunction1_n724) );
  XOR2_X1 LED_RoundFunction1_U245 ( .A(1'b0), .B(LED_RoundFunction1_n723), .Z(
        SubCellInput1[42]) );
  AOI21_X1 LED_RoundFunction1_U244 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n722), .A(LED_RoundFunction1_n721), .ZN(
        LED_RoundFunction1_n723) );
  AOI221_X1 LED_RoundFunction1_U243 ( .B1(Plaintext1[42]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_42_), .C2(LED_RoundFunction1_n568), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n721) );
  INV_X1 LED_RoundFunction1_U242 ( .A(Ciphertext1[42]), .ZN(
        LED_RoundFunction1_n722) );
  XOR2_X1 LED_RoundFunction1_U241 ( .A(1'b0), .B(LED_RoundFunction1_n720), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[2]) );
  AOI21_X1 LED_RoundFunction1_U240 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n719), .A(LED_RoundFunction1_n718), .ZN(
        LED_RoundFunction1_n720) );
  AOI221_X1 LED_RoundFunction1_U239 ( .B1(Plaintext1[41]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_41_), .C2(LED_RoundFunction1_n565), .A(
        LED_RoundFunction1_n557), .ZN(LED_RoundFunction1_n718) );
  INV_X1 LED_RoundFunction1_U238 ( .A(Ciphertext1[41]), .ZN(
        LED_RoundFunction1_n719) );
  XOR2_X1 LED_RoundFunction1_U237 ( .A(1'b0), .B(LED_RoundFunction1_n717), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[0]) );
  AOI21_X1 LED_RoundFunction1_U236 ( .B1(LED_RoundFunction1_n557), .B2(
        LED_RoundFunction1_n716), .A(LED_RoundFunction1_n715), .ZN(
        LED_RoundFunction1_n717) );
  AOI221_X1 LED_RoundFunction1_U235 ( .B1(Plaintext1[40]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_40_), .C2(LED_RoundFunction1_n568), .A(
        LED_RoundFunction1_n557), .ZN(LED_RoundFunction1_n715) );
  INV_X1 LED_RoundFunction1_U234 ( .A(Ciphertext1[40]), .ZN(
        LED_RoundFunction1_n716) );
  AOI22_X1 LED_RoundFunction1_U233 ( .A1(LED_RoundFunction1_n556), .A2(
        Ciphertext1[29]), .B1(LED_RoundFunction1_n714), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[2]) );
  INV_X1 LED_RoundFunction1_U232 ( .A(LED_RoundFunction1_n713), .ZN(
        LED_RoundFunction1_n714) );
  OAI22_X1 LED_RoundFunction1_U231 ( .A1(LED_RoundFunction1_n565), .A2(
        Plaintext1[29]), .B1(LED_RoundFunction1_Feedback_29_), .B2(rst), .ZN(
        LED_RoundFunction1_n713) );
  XOR2_X1 LED_RoundFunction1_U230 ( .A(1'b0), .B(LED_RoundFunction1_n712), .Z(
        SubCellInput1[26]) );
  AOI21_X1 LED_RoundFunction1_U229 ( .B1(LED_RoundFunction1_n558), .B2(
        LED_RoundFunction1_n711), .A(LED_RoundFunction1_n710), .ZN(
        LED_RoundFunction1_n712) );
  AOI221_X1 LED_RoundFunction1_U228 ( .B1(Plaintext1[26]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_26_), .C2(LED_RoundFunction1_n568), .A(
        LED_RoundFunction1_n557), .ZN(LED_RoundFunction1_n710) );
  INV_X1 LED_RoundFunction1_U227 ( .A(Ciphertext1[26]), .ZN(
        LED_RoundFunction1_n711) );
  XOR2_X1 LED_RoundFunction1_U226 ( .A(1'b0), .B(LED_RoundFunction1_n709), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[2]) );
  AOI21_X1 LED_RoundFunction1_U225 ( .B1(LED_RoundFunction1_n558), .B2(
        LED_RoundFunction1_n708), .A(LED_RoundFunction1_n707), .ZN(
        LED_RoundFunction1_n709) );
  AOI221_X1 LED_RoundFunction1_U224 ( .B1(Plaintext1[25]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_25_), .C2(LED_RoundFunction1_n568), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n707) );
  INV_X1 LED_RoundFunction1_U223 ( .A(Ciphertext1[25]), .ZN(
        LED_RoundFunction1_n708) );
  XOR2_X1 LED_RoundFunction1_U222 ( .A(1'b0), .B(LED_RoundFunction1_n706), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[0]) );
  AOI21_X1 LED_RoundFunction1_U221 ( .B1(LED_RoundFunction1_n558), .B2(
        LED_RoundFunction1_n705), .A(LED_RoundFunction1_n704), .ZN(
        LED_RoundFunction1_n706) );
  AOI221_X1 LED_RoundFunction1_U220 ( .B1(Plaintext1[24]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_24_), .C2(LED_RoundFunction1_n566), .A(
        LED_RoundFunction1_n557), .ZN(LED_RoundFunction1_n704) );
  INV_X1 LED_RoundFunction1_U219 ( .A(Ciphertext1[24]), .ZN(
        LED_RoundFunction1_n705) );
  AOI22_X1 LED_RoundFunction1_U218 ( .A1(LED_RoundFunction1_n556), .A2(
        Ciphertext1[13]), .B1(LED_RoundFunction1_n703), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[2]) );
  INV_X1 LED_RoundFunction1_U217 ( .A(LED_RoundFunction1_n702), .ZN(
        LED_RoundFunction1_n703) );
  OAI22_X1 LED_RoundFunction1_U216 ( .A1(LED_RoundFunction1_n568), .A2(
        Plaintext1[13]), .B1(LED_RoundFunction1_Feedback_13_), .B2(rst), .ZN(
        LED_RoundFunction1_n702) );
  AOI22_X1 LED_RoundFunction1_U215 ( .A1(LED_RoundFunction1_n556), .A2(
        Ciphertext1[12]), .B1(LED_RoundFunction1_n701), .B2(
        LED_RoundFunction1_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[0]) );
  INV_X1 LED_RoundFunction1_U214 ( .A(LED_RoundFunction1_n700), .ZN(
        LED_RoundFunction1_n701) );
  OAI22_X1 LED_RoundFunction1_U213 ( .A1(LED_RoundFunction1_n565), .A2(
        Plaintext1[12]), .B1(LED_RoundFunction1_Feedback_12_), .B2(rst), .ZN(
        LED_RoundFunction1_n700) );
  XOR2_X1 LED_RoundFunction1_U212 ( .A(1'b0), .B(LED_RoundFunction1_n699), .Z(
        SubCellInput1[10]) );
  AOI21_X1 LED_RoundFunction1_U211 ( .B1(LED_RoundFunction1_n558), .B2(
        LED_RoundFunction1_n698), .A(LED_RoundFunction1_n697), .ZN(
        LED_RoundFunction1_n699) );
  AOI221_X1 LED_RoundFunction1_U210 ( .B1(Plaintext1[10]), .B2(rst), .C1(
        LED_RoundFunction1_Feedback_10_), .C2(LED_RoundFunction1_n565), .A(
        LED_RoundFunction1_n556), .ZN(LED_RoundFunction1_n697) );
  INV_X1 LED_RoundFunction1_U209 ( .A(Ciphertext1[10]), .ZN(
        LED_RoundFunction1_n698) );
  AOI22_X1 LED_RoundFunction1_U208 ( .A1(rst), .A2(LED_RoundFunction1_n696), 
        .B1(LED_RoundFunction1_n695), .B2(LED_RoundFunction1_n563), .ZN(
        Ciphertext1[9]) );
  XNOR2_X1 LED_RoundFunction1_U207 ( .A(LED_RoundFunction1_Feedback_9_), .B(
        Key1[73]), .ZN(LED_RoundFunction1_n695) );
  XNOR2_X1 LED_RoundFunction1_U206 ( .A(Plaintext1[9]), .B(Key1[9]), .ZN(
        LED_RoundFunction1_n696) );
  AOI22_X1 LED_RoundFunction1_U205 ( .A1(rst), .A2(LED_RoundFunction1_n694), 
        .B1(LED_RoundFunction1_n693), .B2(LED_RoundFunction1_n563), .ZN(
        Ciphertext1[8]) );
  XNOR2_X1 LED_RoundFunction1_U204 ( .A(LED_RoundFunction1_Feedback_8_), .B(
        Key1[72]), .ZN(LED_RoundFunction1_n693) );
  XNOR2_X1 LED_RoundFunction1_U203 ( .A(Plaintext1[8]), .B(Key1[8]), .ZN(
        LED_RoundFunction1_n694) );
  AOI22_X1 LED_RoundFunction1_U202 ( .A1(rst), .A2(LED_RoundFunction1_n692), 
        .B1(LED_RoundFunction1_n691), .B2(LED_RoundFunction1_n563), .ZN(
        Ciphertext1[7]) );
  XNOR2_X1 LED_RoundFunction1_U201 ( .A(LED_RoundFunction1_Feedback_7_), .B(
        Key1[71]), .ZN(LED_RoundFunction1_n691) );
  XNOR2_X1 LED_RoundFunction1_U200 ( .A(Plaintext1[7]), .B(Key1[7]), .ZN(
        LED_RoundFunction1_n692) );
  AOI22_X1 LED_RoundFunction1_U199 ( .A1(rst), .A2(LED_RoundFunction1_n690), 
        .B1(LED_RoundFunction1_n689), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[6]) );
  XNOR2_X1 LED_RoundFunction1_U198 ( .A(LED_RoundFunction1_Feedback_6_), .B(
        Key1[70]), .ZN(LED_RoundFunction1_n689) );
  XNOR2_X1 LED_RoundFunction1_U197 ( .A(Plaintext1[6]), .B(Key1[6]), .ZN(
        LED_RoundFunction1_n690) );
  AOI22_X1 LED_RoundFunction1_U196 ( .A1(rst), .A2(LED_RoundFunction1_n688), 
        .B1(LED_RoundFunction1_n687), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[63]) );
  XNOR2_X1 LED_RoundFunction1_U195 ( .A(LED_RoundFunction1_Feedback_63_), .B(
        Key1[127]), .ZN(LED_RoundFunction1_n687) );
  XNOR2_X1 LED_RoundFunction1_U194 ( .A(Plaintext1[63]), .B(Key1[63]), .ZN(
        LED_RoundFunction1_n688) );
  AOI22_X1 LED_RoundFunction1_U193 ( .A1(rst), .A2(LED_RoundFunction1_n686), 
        .B1(LED_RoundFunction1_n685), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[5]) );
  XNOR2_X1 LED_RoundFunction1_U192 ( .A(LED_RoundFunction1_Feedback_5_), .B(
        Key1[69]), .ZN(LED_RoundFunction1_n685) );
  XNOR2_X1 LED_RoundFunction1_U191 ( .A(Plaintext1[5]), .B(Key1[5]), .ZN(
        LED_RoundFunction1_n686) );
  AOI22_X1 LED_RoundFunction1_U190 ( .A1(rst), .A2(LED_RoundFunction1_n684), 
        .B1(LED_RoundFunction1_n683), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[58]) );
  XNOR2_X1 LED_RoundFunction1_U189 ( .A(LED_RoundFunction1_Feedback_58_), .B(
        Key1[122]), .ZN(LED_RoundFunction1_n683) );
  XNOR2_X1 LED_RoundFunction1_U188 ( .A(Plaintext1[58]), .B(Key1[58]), .ZN(
        LED_RoundFunction1_n684) );
  AOI22_X1 LED_RoundFunction1_U187 ( .A1(rst), .A2(LED_RoundFunction1_n682), 
        .B1(LED_RoundFunction1_n681), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[57]) );
  XNOR2_X1 LED_RoundFunction1_U186 ( .A(LED_RoundFunction1_Feedback_57_), .B(
        Key1[121]), .ZN(LED_RoundFunction1_n681) );
  XNOR2_X1 LED_RoundFunction1_U185 ( .A(Plaintext1[57]), .B(Key1[57]), .ZN(
        LED_RoundFunction1_n682) );
  AOI22_X1 LED_RoundFunction1_U184 ( .A1(rst), .A2(LED_RoundFunction1_n680), 
        .B1(LED_RoundFunction1_n679), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[56]) );
  XNOR2_X1 LED_RoundFunction1_U183 ( .A(LED_RoundFunction1_Feedback_56_), .B(
        Key1[120]), .ZN(LED_RoundFunction1_n679) );
  XNOR2_X1 LED_RoundFunction1_U182 ( .A(Plaintext1[56]), .B(Key1[56]), .ZN(
        LED_RoundFunction1_n680) );
  AOI22_X1 LED_RoundFunction1_U181 ( .A1(rst), .A2(LED_RoundFunction1_n678), 
        .B1(LED_RoundFunction1_n677), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[55]) );
  XNOR2_X1 LED_RoundFunction1_U180 ( .A(LED_RoundFunction1_Feedback_55_), .B(
        Key1[119]), .ZN(LED_RoundFunction1_n677) );
  XNOR2_X1 LED_RoundFunction1_U179 ( .A(Plaintext1[55]), .B(Key1[55]), .ZN(
        LED_RoundFunction1_n678) );
  AOI22_X1 LED_RoundFunction1_U178 ( .A1(rst), .A2(LED_RoundFunction1_n676), 
        .B1(LED_RoundFunction1_n675), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[54]) );
  XNOR2_X1 LED_RoundFunction1_U177 ( .A(LED_RoundFunction1_Feedback_54_), .B(
        Key1[118]), .ZN(LED_RoundFunction1_n675) );
  XNOR2_X1 LED_RoundFunction1_U176 ( .A(Plaintext1[54]), .B(Key1[54]), .ZN(
        LED_RoundFunction1_n676) );
  AOI22_X1 LED_RoundFunction1_U175 ( .A1(rst), .A2(LED_RoundFunction1_n674), 
        .B1(LED_RoundFunction1_n673), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[53]) );
  XNOR2_X1 LED_RoundFunction1_U174 ( .A(LED_RoundFunction1_Feedback_53_), .B(
        Key1[117]), .ZN(LED_RoundFunction1_n673) );
  XNOR2_X1 LED_RoundFunction1_U173 ( .A(Plaintext1[53]), .B(Key1[53]), .ZN(
        LED_RoundFunction1_n674) );
  AOI22_X1 LED_RoundFunction1_U172 ( .A1(rst), .A2(LED_RoundFunction1_n672), 
        .B1(LED_RoundFunction1_n671), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[52]) );
  XNOR2_X1 LED_RoundFunction1_U171 ( .A(LED_RoundFunction1_Feedback_52_), .B(
        Key1[116]), .ZN(LED_RoundFunction1_n671) );
  XNOR2_X1 LED_RoundFunction1_U170 ( .A(Plaintext1[52]), .B(Key1[52]), .ZN(
        LED_RoundFunction1_n672) );
  AOI22_X1 LED_RoundFunction1_U169 ( .A1(rst), .A2(LED_RoundFunction1_n670), 
        .B1(LED_RoundFunction1_n669), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[51]) );
  XNOR2_X1 LED_RoundFunction1_U168 ( .A(LED_RoundFunction1_Feedback_51_), .B(
        Key1[115]), .ZN(LED_RoundFunction1_n669) );
  XNOR2_X1 LED_RoundFunction1_U167 ( .A(Plaintext1[51]), .B(Key1[51]), .ZN(
        LED_RoundFunction1_n670) );
  AOI22_X1 LED_RoundFunction1_U166 ( .A1(rst), .A2(LED_RoundFunction1_n668), 
        .B1(LED_RoundFunction1_n667), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[50]) );
  XNOR2_X1 LED_RoundFunction1_U165 ( .A(LED_RoundFunction1_Feedback_50_), .B(
        Key1[114]), .ZN(LED_RoundFunction1_n667) );
  XNOR2_X1 LED_RoundFunction1_U164 ( .A(Plaintext1[50]), .B(Key1[50]), .ZN(
        LED_RoundFunction1_n668) );
  AOI22_X1 LED_RoundFunction1_U163 ( .A1(rst), .A2(LED_RoundFunction1_n666), 
        .B1(LED_RoundFunction1_n665), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[4]) );
  XNOR2_X1 LED_RoundFunction1_U162 ( .A(LED_RoundFunction1_Feedback_4_), .B(
        Key1[68]), .ZN(LED_RoundFunction1_n665) );
  XNOR2_X1 LED_RoundFunction1_U161 ( .A(Plaintext1[4]), .B(Key1[4]), .ZN(
        LED_RoundFunction1_n666) );
  AOI22_X1 LED_RoundFunction1_U160 ( .A1(rst), .A2(LED_RoundFunction1_n664), 
        .B1(LED_RoundFunction1_n663), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[49]) );
  XNOR2_X1 LED_RoundFunction1_U159 ( .A(LED_RoundFunction1_Feedback_49_), .B(
        Key1[113]), .ZN(LED_RoundFunction1_n663) );
  XNOR2_X1 LED_RoundFunction1_U158 ( .A(Plaintext1[49]), .B(Key1[49]), .ZN(
        LED_RoundFunction1_n664) );
  AOI22_X1 LED_RoundFunction1_U157 ( .A1(rst), .A2(LED_RoundFunction1_n662), 
        .B1(LED_RoundFunction1_n661), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[48]) );
  XNOR2_X1 LED_RoundFunction1_U156 ( .A(LED_RoundFunction1_Feedback_48_), .B(
        Key1[112]), .ZN(LED_RoundFunction1_n661) );
  XNOR2_X1 LED_RoundFunction1_U155 ( .A(Plaintext1[48]), .B(Key1[48]), .ZN(
        LED_RoundFunction1_n662) );
  AOI22_X1 LED_RoundFunction1_U154 ( .A1(rst), .A2(LED_RoundFunction1_n660), 
        .B1(LED_RoundFunction1_n659), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[47]) );
  XNOR2_X1 LED_RoundFunction1_U153 ( .A(LED_RoundFunction1_Feedback_47_), .B(
        Key1[111]), .ZN(LED_RoundFunction1_n659) );
  XNOR2_X1 LED_RoundFunction1_U152 ( .A(Plaintext1[47]), .B(Key1[47]), .ZN(
        LED_RoundFunction1_n660) );
  AOI22_X1 LED_RoundFunction1_U151 ( .A1(rst), .A2(LED_RoundFunction1_n658), 
        .B1(LED_RoundFunction1_n657), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[44]) );
  XNOR2_X1 LED_RoundFunction1_U150 ( .A(LED_RoundFunction1_Feedback_44_), .B(
        Key1[108]), .ZN(LED_RoundFunction1_n657) );
  XNOR2_X1 LED_RoundFunction1_U149 ( .A(Plaintext1[44]), .B(Key1[44]), .ZN(
        LED_RoundFunction1_n658) );
  AOI22_X1 LED_RoundFunction1_U148 ( .A1(rst), .A2(LED_RoundFunction1_n656), 
        .B1(LED_RoundFunction1_n655), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[42]) );
  XNOR2_X1 LED_RoundFunction1_U147 ( .A(LED_RoundFunction1_Feedback_42_), .B(
        Key1[106]), .ZN(LED_RoundFunction1_n655) );
  XNOR2_X1 LED_RoundFunction1_U146 ( .A(Plaintext1[42]), .B(Key1[42]), .ZN(
        LED_RoundFunction1_n656) );
  AOI22_X1 LED_RoundFunction1_U145 ( .A1(rst), .A2(LED_RoundFunction1_n654), 
        .B1(LED_RoundFunction1_n653), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[41]) );
  XNOR2_X1 LED_RoundFunction1_U144 ( .A(LED_RoundFunction1_Feedback_41_), .B(
        Key1[105]), .ZN(LED_RoundFunction1_n653) );
  XNOR2_X1 LED_RoundFunction1_U143 ( .A(Plaintext1[41]), .B(Key1[41]), .ZN(
        LED_RoundFunction1_n654) );
  AOI22_X1 LED_RoundFunction1_U142 ( .A1(rst), .A2(LED_RoundFunction1_n652), 
        .B1(LED_RoundFunction1_n651), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[40]) );
  XNOR2_X1 LED_RoundFunction1_U141 ( .A(LED_RoundFunction1_Feedback_40_), .B(
        Key1[104]), .ZN(LED_RoundFunction1_n651) );
  XNOR2_X1 LED_RoundFunction1_U140 ( .A(Plaintext1[40]), .B(Key1[40]), .ZN(
        LED_RoundFunction1_n652) );
  AOI22_X1 LED_RoundFunction1_U139 ( .A1(rst), .A2(LED_RoundFunction1_n650), 
        .B1(LED_RoundFunction1_n649), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[3]) );
  XNOR2_X1 LED_RoundFunction1_U138 ( .A(LED_RoundFunction1_Feedback_3_), .B(
        Key1[67]), .ZN(LED_RoundFunction1_n649) );
  XNOR2_X1 LED_RoundFunction1_U137 ( .A(Plaintext1[3]), .B(Key1[3]), .ZN(
        LED_RoundFunction1_n650) );
  AOI22_X1 LED_RoundFunction1_U136 ( .A1(rst), .A2(LED_RoundFunction1_n648), 
        .B1(LED_RoundFunction1_n647), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[39]) );
  XNOR2_X1 LED_RoundFunction1_U135 ( .A(LED_RoundFunction1_Feedback_39_), .B(
        Key1[103]), .ZN(LED_RoundFunction1_n647) );
  XNOR2_X1 LED_RoundFunction1_U134 ( .A(Plaintext1[39]), .B(Key1[39]), .ZN(
        LED_RoundFunction1_n648) );
  AOI22_X1 LED_RoundFunction1_U133 ( .A1(rst), .A2(LED_RoundFunction1_n646), 
        .B1(LED_RoundFunction1_n645), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[38]) );
  XNOR2_X1 LED_RoundFunction1_U132 ( .A(LED_RoundFunction1_Feedback_38_), .B(
        Key1[102]), .ZN(LED_RoundFunction1_n645) );
  XNOR2_X1 LED_RoundFunction1_U131 ( .A(Plaintext1[38]), .B(Key1[38]), .ZN(
        LED_RoundFunction1_n646) );
  AOI22_X1 LED_RoundFunction1_U130 ( .A1(rst), .A2(LED_RoundFunction1_n644), 
        .B1(LED_RoundFunction1_n643), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[37]) );
  XNOR2_X1 LED_RoundFunction1_U129 ( .A(LED_RoundFunction1_Feedback_37_), .B(
        Key1[101]), .ZN(LED_RoundFunction1_n643) );
  XNOR2_X1 LED_RoundFunction1_U128 ( .A(Plaintext1[37]), .B(Key1[37]), .ZN(
        LED_RoundFunction1_n644) );
  AOI22_X1 LED_RoundFunction1_U127 ( .A1(rst), .A2(LED_RoundFunction1_n642), 
        .B1(LED_RoundFunction1_n641), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[36]) );
  XNOR2_X1 LED_RoundFunction1_U126 ( .A(LED_RoundFunction1_Feedback_36_), .B(
        Key1[100]), .ZN(LED_RoundFunction1_n641) );
  XNOR2_X1 LED_RoundFunction1_U125 ( .A(Plaintext1[36]), .B(Key1[36]), .ZN(
        LED_RoundFunction1_n642) );
  AOI22_X1 LED_RoundFunction1_U124 ( .A1(rst), .A2(LED_RoundFunction1_n640), 
        .B1(LED_RoundFunction1_n639), .B2(LED_RoundFunction1_n568), .ZN(
        Ciphertext1[35]) );
  XNOR2_X1 LED_RoundFunction1_U123 ( .A(LED_RoundFunction1_Feedback_35_), .B(
        Key1[99]), .ZN(LED_RoundFunction1_n639) );
  XNOR2_X1 LED_RoundFunction1_U122 ( .A(Plaintext1[35]), .B(Key1[35]), .ZN(
        LED_RoundFunction1_n640) );
  AOI22_X1 LED_RoundFunction1_U121 ( .A1(rst), .A2(LED_RoundFunction1_n638), 
        .B1(LED_RoundFunction1_n637), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[34]) );
  XNOR2_X1 LED_RoundFunction1_U120 ( .A(LED_RoundFunction1_Feedback_34_), .B(
        Key1[98]), .ZN(LED_RoundFunction1_n637) );
  XNOR2_X1 LED_RoundFunction1_U119 ( .A(Plaintext1[34]), .B(Key1[34]), .ZN(
        LED_RoundFunction1_n638) );
  AOI22_X1 LED_RoundFunction1_U118 ( .A1(rst), .A2(LED_RoundFunction1_n636), 
        .B1(LED_RoundFunction1_n635), .B2(LED_RoundFunction1_n568), .ZN(
        Ciphertext1[33]) );
  XNOR2_X1 LED_RoundFunction1_U117 ( .A(LED_RoundFunction1_Feedback_33_), .B(
        Key1[97]), .ZN(LED_RoundFunction1_n635) );
  XNOR2_X1 LED_RoundFunction1_U116 ( .A(Plaintext1[33]), .B(Key1[33]), .ZN(
        LED_RoundFunction1_n636) );
  AOI22_X1 LED_RoundFunction1_U115 ( .A1(rst), .A2(LED_RoundFunction1_n634), 
        .B1(LED_RoundFunction1_n633), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[32]) );
  XNOR2_X1 LED_RoundFunction1_U114 ( .A(LED_RoundFunction1_Feedback_32_), .B(
        Key1[96]), .ZN(LED_RoundFunction1_n633) );
  XNOR2_X1 LED_RoundFunction1_U113 ( .A(Plaintext1[32]), .B(Key1[32]), .ZN(
        LED_RoundFunction1_n634) );
  AOI22_X1 LED_RoundFunction1_U112 ( .A1(rst), .A2(LED_RoundFunction1_n632), 
        .B1(LED_RoundFunction1_n631), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[2]) );
  XNOR2_X1 LED_RoundFunction1_U111 ( .A(LED_RoundFunction1_Feedback_2_), .B(
        Key1[66]), .ZN(LED_RoundFunction1_n631) );
  XNOR2_X1 LED_RoundFunction1_U110 ( .A(Plaintext1[2]), .B(Key1[2]), .ZN(
        LED_RoundFunction1_n632) );
  AOI22_X1 LED_RoundFunction1_U109 ( .A1(rst), .A2(LED_RoundFunction1_n630), 
        .B1(LED_RoundFunction1_n629), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[29]) );
  XNOR2_X1 LED_RoundFunction1_U108 ( .A(LED_RoundFunction1_Feedback_29_), .B(
        Key1[93]), .ZN(LED_RoundFunction1_n629) );
  XNOR2_X1 LED_RoundFunction1_U107 ( .A(Plaintext1[29]), .B(Key1[29]), .ZN(
        LED_RoundFunction1_n630) );
  AOI22_X1 LED_RoundFunction1_U106 ( .A1(rst), .A2(LED_RoundFunction1_n628), 
        .B1(LED_RoundFunction1_n627), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[26]) );
  XNOR2_X1 LED_RoundFunction1_U105 ( .A(LED_RoundFunction1_Feedback_26_), .B(
        Key1[90]), .ZN(LED_RoundFunction1_n627) );
  XNOR2_X1 LED_RoundFunction1_U104 ( .A(Plaintext1[26]), .B(Key1[26]), .ZN(
        LED_RoundFunction1_n628) );
  AOI22_X1 LED_RoundFunction1_U103 ( .A1(rst), .A2(LED_RoundFunction1_n626), 
        .B1(LED_RoundFunction1_n625), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[25]) );
  XNOR2_X1 LED_RoundFunction1_U102 ( .A(LED_RoundFunction1_Feedback_25_), .B(
        Key1[89]), .ZN(LED_RoundFunction1_n625) );
  XNOR2_X1 LED_RoundFunction1_U101 ( .A(Plaintext1[25]), .B(Key1[25]), .ZN(
        LED_RoundFunction1_n626) );
  AOI22_X1 LED_RoundFunction1_U100 ( .A1(rst), .A2(LED_RoundFunction1_n624), 
        .B1(LED_RoundFunction1_n623), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[24]) );
  XNOR2_X1 LED_RoundFunction1_U99 ( .A(LED_RoundFunction1_Feedback_24_), .B(
        Key1[88]), .ZN(LED_RoundFunction1_n623) );
  XNOR2_X1 LED_RoundFunction1_U98 ( .A(Plaintext1[24]), .B(Key1[24]), .ZN(
        LED_RoundFunction1_n624) );
  AOI22_X1 LED_RoundFunction1_U97 ( .A1(rst), .A2(LED_RoundFunction1_n622), 
        .B1(LED_RoundFunction1_n621), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[23]) );
  XNOR2_X1 LED_RoundFunction1_U96 ( .A(LED_RoundFunction1_Feedback_23_), .B(
        Key1[87]), .ZN(LED_RoundFunction1_n621) );
  XNOR2_X1 LED_RoundFunction1_U95 ( .A(Plaintext1[23]), .B(Key1[23]), .ZN(
        LED_RoundFunction1_n622) );
  AOI22_X1 LED_RoundFunction1_U94 ( .A1(rst), .A2(LED_RoundFunction1_n620), 
        .B1(LED_RoundFunction1_n619), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[22]) );
  XNOR2_X1 LED_RoundFunction1_U93 ( .A(LED_RoundFunction1_Feedback_22_), .B(
        Key1[86]), .ZN(LED_RoundFunction1_n619) );
  XNOR2_X1 LED_RoundFunction1_U92 ( .A(Plaintext1[22]), .B(Key1[22]), .ZN(
        LED_RoundFunction1_n620) );
  AOI22_X1 LED_RoundFunction1_U91 ( .A1(rst), .A2(LED_RoundFunction1_n618), 
        .B1(LED_RoundFunction1_n617), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[21]) );
  XNOR2_X1 LED_RoundFunction1_U90 ( .A(LED_RoundFunction1_Feedback_21_), .B(
        Key1[85]), .ZN(LED_RoundFunction1_n617) );
  XNOR2_X1 LED_RoundFunction1_U89 ( .A(Plaintext1[21]), .B(Key1[21]), .ZN(
        LED_RoundFunction1_n618) );
  AOI22_X1 LED_RoundFunction1_U88 ( .A1(rst), .A2(LED_RoundFunction1_n616), 
        .B1(LED_RoundFunction1_n615), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[20]) );
  XNOR2_X1 LED_RoundFunction1_U87 ( .A(LED_RoundFunction1_Feedback_20_), .B(
        Key1[84]), .ZN(LED_RoundFunction1_n615) );
  XNOR2_X1 LED_RoundFunction1_U86 ( .A(Plaintext1[20]), .B(Key1[20]), .ZN(
        LED_RoundFunction1_n616) );
  AOI22_X1 LED_RoundFunction1_U85 ( .A1(rst), .A2(LED_RoundFunction1_n614), 
        .B1(LED_RoundFunction1_n613), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[1]) );
  XNOR2_X1 LED_RoundFunction1_U84 ( .A(LED_RoundFunction1_Feedback_1_), .B(
        Key1[65]), .ZN(LED_RoundFunction1_n613) );
  XNOR2_X1 LED_RoundFunction1_U83 ( .A(Plaintext1[1]), .B(Key1[1]), .ZN(
        LED_RoundFunction1_n614) );
  AOI22_X1 LED_RoundFunction1_U82 ( .A1(rst), .A2(LED_RoundFunction1_n612), 
        .B1(LED_RoundFunction1_n611), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[19]) );
  XNOR2_X1 LED_RoundFunction1_U81 ( .A(LED_RoundFunction1_Feedback_19_), .B(
        Key1[83]), .ZN(LED_RoundFunction1_n611) );
  XNOR2_X1 LED_RoundFunction1_U80 ( .A(Plaintext1[19]), .B(Key1[19]), .ZN(
        LED_RoundFunction1_n612) );
  AOI22_X1 LED_RoundFunction1_U79 ( .A1(rst), .A2(LED_RoundFunction1_n610), 
        .B1(LED_RoundFunction1_n609), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[18]) );
  XNOR2_X1 LED_RoundFunction1_U78 ( .A(LED_RoundFunction1_Feedback_18_), .B(
        Key1[82]), .ZN(LED_RoundFunction1_n609) );
  XNOR2_X1 LED_RoundFunction1_U77 ( .A(Plaintext1[18]), .B(Key1[18]), .ZN(
        LED_RoundFunction1_n610) );
  AOI22_X1 LED_RoundFunction1_U76 ( .A1(rst), .A2(LED_RoundFunction1_n608), 
        .B1(LED_RoundFunction1_n607), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[17]) );
  XNOR2_X1 LED_RoundFunction1_U75 ( .A(LED_RoundFunction1_Feedback_17_), .B(
        Key1[81]), .ZN(LED_RoundFunction1_n607) );
  XNOR2_X1 LED_RoundFunction1_U74 ( .A(Plaintext1[17]), .B(Key1[17]), .ZN(
        LED_RoundFunction1_n608) );
  AOI22_X1 LED_RoundFunction1_U73 ( .A1(rst), .A2(LED_RoundFunction1_n606), 
        .B1(LED_RoundFunction1_n605), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[16]) );
  XNOR2_X1 LED_RoundFunction1_U72 ( .A(LED_RoundFunction1_Feedback_16_), .B(
        Key1[80]), .ZN(LED_RoundFunction1_n605) );
  XNOR2_X1 LED_RoundFunction1_U71 ( .A(Plaintext1[16]), .B(Key1[16]), .ZN(
        LED_RoundFunction1_n606) );
  AOI22_X1 LED_RoundFunction1_U70 ( .A1(rst), .A2(LED_RoundFunction1_n604), 
        .B1(LED_RoundFunction1_n603), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[13]) );
  XNOR2_X1 LED_RoundFunction1_U69 ( .A(LED_RoundFunction1_Feedback_13_), .B(
        Key1[77]), .ZN(LED_RoundFunction1_n603) );
  XNOR2_X1 LED_RoundFunction1_U68 ( .A(Plaintext1[13]), .B(Key1[13]), .ZN(
        LED_RoundFunction1_n604) );
  AOI22_X1 LED_RoundFunction1_U67 ( .A1(rst), .A2(LED_RoundFunction1_n602), 
        .B1(LED_RoundFunction1_n601), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[12]) );
  XNOR2_X1 LED_RoundFunction1_U66 ( .A(LED_RoundFunction1_Feedback_12_), .B(
        Key1[76]), .ZN(LED_RoundFunction1_n601) );
  XNOR2_X1 LED_RoundFunction1_U65 ( .A(Plaintext1[12]), .B(Key1[12]), .ZN(
        LED_RoundFunction1_n602) );
  AOI22_X1 LED_RoundFunction1_U64 ( .A1(rst), .A2(LED_RoundFunction1_n600), 
        .B1(LED_RoundFunction1_n599), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[10]) );
  XNOR2_X1 LED_RoundFunction1_U63 ( .A(LED_RoundFunction1_Feedback_10_), .B(
        Key1[74]), .ZN(LED_RoundFunction1_n599) );
  XNOR2_X1 LED_RoundFunction1_U62 ( .A(Plaintext1[10]), .B(Key1[10]), .ZN(
        LED_RoundFunction1_n600) );
  AOI22_X1 LED_RoundFunction1_U61 ( .A1(rst), .A2(LED_RoundFunction1_n598), 
        .B1(LED_RoundFunction1_n597), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[0]) );
  XNOR2_X1 LED_RoundFunction1_U60 ( .A(LED_RoundFunction1_Feedback_0_), .B(
        Key1[64]), .ZN(LED_RoundFunction1_n597) );
  XNOR2_X1 LED_RoundFunction1_U59 ( .A(Plaintext1[0]), .B(Key1[0]), .ZN(
        LED_RoundFunction1_n598) );
  AOI22_X1 LED_RoundFunction1_U58 ( .A1(rst), .A2(LED_RoundFunction1_n596), 
        .B1(LED_RoundFunction1_n595), .B2(LED_RoundFunction1_n568), .ZN(
        Ciphertext1[46]) );
  XNOR2_X1 LED_RoundFunction1_U57 ( .A(LED_RoundFunction1_Feedback_46_), .B(
        Key1[110]), .ZN(LED_RoundFunction1_n595) );
  XNOR2_X1 LED_RoundFunction1_U56 ( .A(Plaintext1[46]), .B(Key1[46]), .ZN(
        LED_RoundFunction1_n596) );
  AOI22_X1 LED_RoundFunction1_U55 ( .A1(rst), .A2(LED_RoundFunction1_n594), 
        .B1(LED_RoundFunction1_n593), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[45]) );
  XNOR2_X1 LED_RoundFunction1_U54 ( .A(LED_RoundFunction1_Feedback_45_), .B(
        Key1[109]), .ZN(LED_RoundFunction1_n593) );
  XNOR2_X1 LED_RoundFunction1_U53 ( .A(Plaintext1[45]), .B(Key1[45]), .ZN(
        LED_RoundFunction1_n594) );
  AOI22_X1 LED_RoundFunction1_U52 ( .A1(rst), .A2(LED_RoundFunction1_n592), 
        .B1(LED_RoundFunction1_n591), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[43]) );
  XNOR2_X1 LED_RoundFunction1_U51 ( .A(LED_RoundFunction1_Feedback_43_), .B(
        Key1[107]), .ZN(LED_RoundFunction1_n591) );
  XNOR2_X1 LED_RoundFunction1_U50 ( .A(Plaintext1[43]), .B(Key1[43]), .ZN(
        LED_RoundFunction1_n592) );
  AOI22_X1 LED_RoundFunction1_U49 ( .A1(rst), .A2(LED_RoundFunction1_n590), 
        .B1(LED_RoundFunction1_n589), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[31]) );
  XNOR2_X1 LED_RoundFunction1_U48 ( .A(LED_RoundFunction1_Feedback_31_), .B(
        Key1[95]), .ZN(LED_RoundFunction1_n589) );
  XNOR2_X1 LED_RoundFunction1_U47 ( .A(Plaintext1[31]), .B(Key1[31]), .ZN(
        LED_RoundFunction1_n590) );
  AOI22_X1 LED_RoundFunction1_U46 ( .A1(rst), .A2(LED_RoundFunction1_n588), 
        .B1(LED_RoundFunction1_n587), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[30]) );
  XNOR2_X1 LED_RoundFunction1_U45 ( .A(LED_RoundFunction1_Feedback_30_), .B(
        Key1[94]), .ZN(LED_RoundFunction1_n587) );
  XNOR2_X1 LED_RoundFunction1_U44 ( .A(Plaintext1[30]), .B(Key1[30]), .ZN(
        LED_RoundFunction1_n588) );
  AOI22_X1 LED_RoundFunction1_U43 ( .A1(rst), .A2(LED_RoundFunction1_n586), 
        .B1(LED_RoundFunction1_n585), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[28]) );
  XNOR2_X1 LED_RoundFunction1_U42 ( .A(LED_RoundFunction1_Feedback_28_), .B(
        Key1[92]), .ZN(LED_RoundFunction1_n585) );
  XNOR2_X1 LED_RoundFunction1_U41 ( .A(Plaintext1[28]), .B(Key1[28]), .ZN(
        LED_RoundFunction1_n586) );
  AOI22_X1 LED_RoundFunction1_U40 ( .A1(rst), .A2(LED_RoundFunction1_n584), 
        .B1(LED_RoundFunction1_n583), .B2(LED_RoundFunction1_n564), .ZN(
        Ciphertext1[27]) );
  XNOR2_X1 LED_RoundFunction1_U39 ( .A(LED_RoundFunction1_Feedback_27_), .B(
        Key1[91]), .ZN(LED_RoundFunction1_n583) );
  XNOR2_X1 LED_RoundFunction1_U38 ( .A(Plaintext1[27]), .B(Key1[27]), .ZN(
        LED_RoundFunction1_n584) );
  AOI22_X1 LED_RoundFunction1_U37 ( .A1(rst), .A2(LED_RoundFunction1_n582), 
        .B1(LED_RoundFunction1_n581), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[15]) );
  XNOR2_X1 LED_RoundFunction1_U36 ( .A(LED_RoundFunction1_Feedback_15_), .B(
        Key1[79]), .ZN(LED_RoundFunction1_n581) );
  XNOR2_X1 LED_RoundFunction1_U35 ( .A(Plaintext1[15]), .B(Key1[15]), .ZN(
        LED_RoundFunction1_n582) );
  AOI22_X1 LED_RoundFunction1_U34 ( .A1(rst), .A2(LED_RoundFunction1_n580), 
        .B1(LED_RoundFunction1_n579), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[14]) );
  XNOR2_X1 LED_RoundFunction1_U33 ( .A(LED_RoundFunction1_Feedback_14_), .B(
        Key1[78]), .ZN(LED_RoundFunction1_n579) );
  XNOR2_X1 LED_RoundFunction1_U32 ( .A(Plaintext1[14]), .B(Key1[14]), .ZN(
        LED_RoundFunction1_n580) );
  AOI22_X1 LED_RoundFunction1_U31 ( .A1(rst), .A2(LED_RoundFunction1_n578), 
        .B1(LED_RoundFunction1_n577), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[11]) );
  XNOR2_X1 LED_RoundFunction1_U30 ( .A(LED_RoundFunction1_Feedback_11_), .B(
        Key1[75]), .ZN(LED_RoundFunction1_n577) );
  XNOR2_X1 LED_RoundFunction1_U29 ( .A(Plaintext1[11]), .B(Key1[11]), .ZN(
        LED_RoundFunction1_n578) );
  AOI22_X1 LED_RoundFunction1_U28 ( .A1(rst), .A2(LED_RoundFunction1_n576), 
        .B1(LED_RoundFunction1_n575), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[62]) );
  XNOR2_X1 LED_RoundFunction1_U27 ( .A(LED_RoundFunction1_Feedback_62_), .B(
        Key1[126]), .ZN(LED_RoundFunction1_n575) );
  XNOR2_X1 LED_RoundFunction1_U26 ( .A(Plaintext1[62]), .B(Key1[62]), .ZN(
        LED_RoundFunction1_n576) );
  AOI22_X1 LED_RoundFunction1_U25 ( .A1(rst), .A2(LED_RoundFunction1_n574), 
        .B1(LED_RoundFunction1_n573), .B2(LED_RoundFunction1_n565), .ZN(
        Ciphertext1[61]) );
  XNOR2_X1 LED_RoundFunction1_U24 ( .A(LED_RoundFunction1_Feedback_61_), .B(
        Key1[125]), .ZN(LED_RoundFunction1_n573) );
  XNOR2_X1 LED_RoundFunction1_U23 ( .A(Plaintext1[61]), .B(Key1[61]), .ZN(
        LED_RoundFunction1_n574) );
  AOI22_X1 LED_RoundFunction1_U22 ( .A1(rst), .A2(LED_RoundFunction1_n572), 
        .B1(LED_RoundFunction1_n571), .B2(LED_RoundFunction1_n566), .ZN(
        Ciphertext1[60]) );
  XNOR2_X1 LED_RoundFunction1_U21 ( .A(LED_RoundFunction1_Feedback_60_), .B(
        Key1[124]), .ZN(LED_RoundFunction1_n571) );
  XNOR2_X1 LED_RoundFunction1_U20 ( .A(Plaintext1[60]), .B(Key1[60]), .ZN(
        LED_RoundFunction1_n572) );
  AOI22_X1 LED_RoundFunction1_U19 ( .A1(rst), .A2(LED_RoundFunction1_n570), 
        .B1(LED_RoundFunction1_n569), .B2(LED_RoundFunction1_n567), .ZN(
        Ciphertext1[59]) );
  XNOR2_X1 LED_RoundFunction1_U18 ( .A(LED_RoundFunction1_Feedback_59_), .B(
        Key1[123]), .ZN(LED_RoundFunction1_n569) );
  XNOR2_X1 LED_RoundFunction1_U17 ( .A(Plaintext1[59]), .B(Key1[59]), .ZN(
        LED_RoundFunction1_n570) );
  INV_X1 LED_RoundFunction1_U16 ( .A(LED_RoundFunction1_n559), .ZN(
        LED_RoundFunction1_n557) );
  INV_X1 LED_RoundFunction1_U15 ( .A(rst), .ZN(LED_RoundFunction1_n568) );
  BUF_X1 LED_RoundFunction1_U14 ( .A(LED_RoundFunction1_n568), .Z(
        LED_RoundFunction1_n564) );
  BUF_X1 LED_RoundFunction1_U13 ( .A(LED_RoundFunction1_n568), .Z(
        LED_RoundFunction1_n566) );
  INV_X1 LED_RoundFunction1_U12 ( .A(LED_RoundFunction1_n559), .ZN(
        LED_RoundFunction1_n556) );
  BUF_X1 LED_RoundFunction1_U11 ( .A(LED_RoundFunction1_n568), .Z(
        LED_RoundFunction1_n565) );
  INV_X1 LED_RoundFunction1_U10 ( .A(LED_RoundFunction1_n559), .ZN(
        LED_RoundFunction1_n558) );
  BUF_X1 LED_RoundFunction1_U9 ( .A(LED_RoundFunction1_n568), .Z(
        LED_RoundFunction1_n563) );
  INV_X1 LED_RoundFunction1_U8 ( .A(LED_RoundFunction1_n559), .ZN(
        LED_RoundFunction1_n555) );
  BUF_X1 LED_RoundFunction1_U7 ( .A(LED_RoundFunction1_n568), .Z(
        LED_RoundFunction1_n562) );
  BUF_X1 LED_RoundFunction1_U6 ( .A(LED_RoundFunction1_n561), .Z(
        LED_RoundFunction1_n560) );
  BUF_X1 LED_RoundFunction1_U5 ( .A(LED_RoundFunction1_n568), .Z(
        LED_RoundFunction1_n567) );
  INV_X1 LED_RoundFunction1_U4 ( .A(AddKey), .ZN(LED_RoundFunction1_n561) );
  BUF_X1 LED_RoundFunction1_U3 ( .A(LED_RoundFunction1_n561), .Z(
        LED_RoundFunction1_n559) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U68 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n160), .B(
        LED_RoundFunction1_MCInst1_MC0_n159), .ZN(
        LED_RoundFunction1_Feedback_15_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U67 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n158), .B(SubCellOutput1[62]), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n160) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U66 ( .A(SubCellOutput1[3]), .B(
        LED_RoundFunction1_MCInst1_MC0_n157), .Z(
        LED_RoundFunction1_Feedback_14_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U65 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n156), .B(
        LED_RoundFunction1_MCInst1_MC0_n155), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n157) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U64 ( .A(SubCellOutput1[21]), .B(
        SubCellOutput1[1]), .ZN(LED_RoundFunction1_MCInst1_MC0_n155) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U63 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n154), .B(SubCellOutput1[41]), .Z(
        LED_RoundFunction1_MCInst1_MC0_n156) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U62 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n153), .B(
        LED_RoundFunction1_MCInst1_MC0_n152), .ZN(
        LED_RoundFunction1_Feedback_13_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U61 ( .A(SubCellOutput1[2]), .B(
        SubCellOutput1[40]), .ZN(LED_RoundFunction1_MCInst1_MC0_n152) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U60 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n151), .B(
        LED_RoundFunction1_MCInst1_MC0_n150), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n153) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U59 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n149), .B(
        LED_RoundFunction1_MCInst1_MC0_n148), .ZN(
        LED_RoundFunction1_Feedback_12_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U58 ( .A(SubCellOutput1[23]), .B(
        LED_RoundFunction1_MCInst1_MC0_n147), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n148) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U57 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n146), .B(
        LED_RoundFunction1_MCInst1_MC0_n150), .Z(
        LED_RoundFunction1_MCInst1_MC0_n149) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U56 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n145), .B(
        LED_RoundFunction1_MCInst1_MC0_n159), .Z(
        LED_RoundFunction1_MCInst1_MC0_n150) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC0_U55 ( .A1(SubCellOutput1[21]), .A2(
        SubCellOutput1[22]), .B1(LED_RoundFunction1_MCInst1_MC0_n144), .B2(
        LED_RoundFunction1_MCInst1_MC0_n143), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n146) );
  INV_X1 LED_RoundFunction1_MCInst1_MC0_U54 ( .A(SubCellOutput1[21]), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n143) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U53 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n142), .B(
        LED_RoundFunction1_MCInst1_MC0_n141), .ZN(
        LED_RoundFunction1_Feedback_31_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U52 ( .A(SubCellOutput1[43]), .B(
        LED_RoundFunction1_MCInst1_MC0_n140), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n141) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U51 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n139), .B(SubCellOutput1[60]), .Z(
        LED_RoundFunction1_MCInst1_MC0_n142) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC0_U50 ( .A1(SubCellOutput1[42]), .A2(
        SubCellOutput1[22]), .B1(LED_RoundFunction1_MCInst1_MC0_n144), .B2(
        LED_RoundFunction1_MCInst1_MC0_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n139) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U49 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n137), .B(
        LED_RoundFunction1_MCInst1_MC0_n136), .ZN(
        LED_RoundFunction1_Feedback_30_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U48 ( .A(SubCellOutput1[40]), .B(
        LED_RoundFunction1_MCInst1_MC0_n135), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n136) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U47 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n134), .B(
        LED_RoundFunction1_MCInst1_MC0_n133), .Z(
        LED_RoundFunction1_MCInst1_MC0_n137) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC0_U46 ( .A1(SubCellOutput1[22]), .A2(
        SubCellOutput1[61]), .B1(LED_RoundFunction1_MCInst1_MC0_n132), .B2(
        LED_RoundFunction1_MCInst1_MC0_n144), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n134) );
  INV_X1 LED_RoundFunction1_MCInst1_MC0_U45 ( .A(SubCellOutput1[22]), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n144) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U44 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n131), .B(
        LED_RoundFunction1_MCInst1_MC0_n151), .ZN(
        LED_RoundFunction1_Feedback_29_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U43 ( .A(SubCellOutput1[63]), .B(
        SubCellOutput1[60]), .ZN(LED_RoundFunction1_MCInst1_MC0_n151) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U42 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n130), .B(
        LED_RoundFunction1_MCInst1_MC0_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n131) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U41 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n128), .B(
        LED_RoundFunction1_MCInst1_MC0_n127), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n130) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U40 ( .A(SubCellOutput1[21]), .B(
        LED_RoundFunction1_MCInst1_MC0_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n127) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U39 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n125), .B(SubCellOutput1[20]), .Z(
        LED_RoundFunction1_MCInst1_MC0_n128) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U38 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n124), .B(
        LED_RoundFunction1_MCInst1_MC0_n123), .ZN(
        LED_RoundFunction1_Feedback_28_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U37 ( .A(SubCellOutput1[0]), .B(
        LED_RoundFunction1_MCInst1_MC0_n122), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n124) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U36 ( .A(SubCellOutput1[2]), .B(
        LED_RoundFunction1_MCInst1_MC0_n122), .ZN(
        LED_RoundFunction1_Feedback_47_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U35 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n135), .B(
        LED_RoundFunction1_MCInst1_MC0_n121), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n122) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U34 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n120), .B(
        LED_RoundFunction1_MCInst1_MC0_n125), .Z(
        LED_RoundFunction1_MCInst1_MC0_n135) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U33 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n119), .B(
        LED_RoundFunction1_MCInst1_MC0_n118), .ZN(
        LED_RoundFunction1_Feedback_46_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U32 ( .A(SubCellOutput1[22]), .B(
        LED_RoundFunction1_MCInst1_MC0_n145), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n118) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U31 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n140), .B(
        LED_RoundFunction1_MCInst1_MC0_n147), .Z(
        LED_RoundFunction1_MCInst1_MC0_n119) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U30 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n126), .B(
        LED_RoundFunction1_MCInst1_MC0_n117), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n140) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U29 ( .A(SubCellOutput1[0]), .B(
        LED_RoundFunction1_MCInst1_MC0_n116), .ZN(
        LED_RoundFunction1_Feedback_45_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U28 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n115), .B(
        LED_RoundFunction1_MCInst1_MC0_n114), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n116) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U27 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n158), .B(SubCellOutput1[61]), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n115) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U26 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n120), .B(
        LED_RoundFunction1_MCInst1_MC0_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n158) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U25 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n113), .B(
        LED_RoundFunction1_MCInst1_MC0_n112), .ZN(
        LED_RoundFunction1_Feedback_44_) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC0_U24 ( .A1(SubCellOutput1[42]), .A2(
        LED_RoundFunction1_MCInst1_MC0_n111), .B1(
        LED_RoundFunction1_MCInst1_MC0_n129), .B2(
        LED_RoundFunction1_MCInst1_MC0_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n112) );
  INV_X1 LED_RoundFunction1_MCInst1_MC0_U23 ( .A(SubCellOutput1[42]), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n138) );
  INV_X1 LED_RoundFunction1_MCInst1_MC0_U22 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n111), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n129) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U21 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n145), .B(
        LED_RoundFunction1_MCInst1_MC0_n154), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n113) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC0_U20 ( .A1(SubCellOutput1[61]), .A2(
        SubCellOutput1[20]), .B1(LED_RoundFunction1_MCInst1_MC0_n110), .B2(
        LED_RoundFunction1_MCInst1_MC0_n132), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n154) );
  INV_X1 LED_RoundFunction1_MCInst1_MC0_U19 ( .A(SubCellOutput1[61]), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n132) );
  INV_X1 LED_RoundFunction1_MCInst1_MC0_U18 ( .A(SubCellOutput1[20]), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n110) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U17 ( .A(SubCellOutput1[3]), .B(
        SubCellOutput1[43]), .Z(LED_RoundFunction1_MCInst1_MC0_n145) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U16 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n111), .B(
        LED_RoundFunction1_MCInst1_MC0_n123), .ZN(
        LED_RoundFunction1_Feedback_63_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U15 ( .A(SubCellOutput1[61]), .B(
        SubCellOutput1[43]), .ZN(LED_RoundFunction1_MCInst1_MC0_n123) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U14 ( .A(SubCellOutput1[22]), .B(
        SubCellOutput1[2]), .Z(LED_RoundFunction1_MCInst1_MC0_n111) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U13 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n120), .B(
        LED_RoundFunction1_MCInst1_MC0_n121), .Z(
        LED_RoundFunction1_Feedback_62_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U12 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n147), .B(SubCellOutput1[60]), .Z(
        LED_RoundFunction1_MCInst1_MC0_n121) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U11 ( .A(SubCellOutput1[1]), .B(
        SubCellOutput1[63]), .Z(LED_RoundFunction1_MCInst1_MC0_n147) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U10 ( .A(SubCellOutput1[42]), .B(
        SubCellOutput1[21]), .Z(LED_RoundFunction1_MCInst1_MC0_n120) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U9 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n117), .B(
        LED_RoundFunction1_MCInst1_MC0_n109), .ZN(
        LED_RoundFunction1_Feedback_61_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U8 ( .A(SubCellOutput1[62]), .B(
        LED_RoundFunction1_MCInst1_MC0_n133), .Z(
        LED_RoundFunction1_MCInst1_MC0_n109) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U7 ( .A(SubCellOutput1[3]), .B(
        SubCellOutput1[63]), .Z(LED_RoundFunction1_MCInst1_MC0_n133) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U6 ( .A(
        LED_RoundFunction1_MCInst1_MC0_n159), .B(
        LED_RoundFunction1_MCInst1_MC0_n125), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n117) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U5 ( .A(SubCellOutput1[23]), .B(
        SubCellOutput1[41]), .Z(LED_RoundFunction1_MCInst1_MC0_n125) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U4 ( .A(SubCellOutput1[0]), .B(
        SubCellOutput1[20]), .Z(LED_RoundFunction1_MCInst1_MC0_n159) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U3 ( .A(SubCellOutput1[3]), .B(
        LED_RoundFunction1_MCInst1_MC0_n114), .ZN(
        LED_RoundFunction1_Feedback_60_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC0_U2 ( .A(SubCellOutput1[23]), .B(
        LED_RoundFunction1_MCInst1_MC0_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC0_n114) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC0_U1 ( .A(SubCellOutput1[62]), .B(
        SubCellOutput1[40]), .Z(LED_RoundFunction1_MCInst1_MC0_n126) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U68 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n160), .B(
        LED_RoundFunction1_MCInst1_MC1_n159), .ZN(
        LED_RoundFunction1_Feedback_11_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U67 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n158), .B(SubCellOutput1[58]), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n160) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U66 ( .A(SubCellOutput1[15]), .B(
        LED_RoundFunction1_MCInst1_MC1_n157), .Z(
        LED_RoundFunction1_Feedback_10_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U65 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n156), .B(
        LED_RoundFunction1_MCInst1_MC1_n155), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n157) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U64 ( .A(SubCellOutput1[17]), .B(
        SubCellOutput1[13]), .ZN(LED_RoundFunction1_MCInst1_MC1_n155) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U63 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n154), .B(SubCellOutput1[37]), .Z(
        LED_RoundFunction1_MCInst1_MC1_n156) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U62 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n153), .B(
        LED_RoundFunction1_MCInst1_MC1_n152), .ZN(
        LED_RoundFunction1_Feedback_9_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U61 ( .A(SubCellOutput1[14]), .B(
        SubCellOutput1[36]), .ZN(LED_RoundFunction1_MCInst1_MC1_n152) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U60 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n151), .B(
        LED_RoundFunction1_MCInst1_MC1_n150), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n153) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U59 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n149), .B(
        LED_RoundFunction1_MCInst1_MC1_n148), .ZN(
        LED_RoundFunction1_Feedback_8_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U58 ( .A(SubCellOutput1[19]), .B(
        LED_RoundFunction1_MCInst1_MC1_n147), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n148) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U57 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n146), .B(
        LED_RoundFunction1_MCInst1_MC1_n150), .Z(
        LED_RoundFunction1_MCInst1_MC1_n149) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U56 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n145), .B(
        LED_RoundFunction1_MCInst1_MC1_n159), .Z(
        LED_RoundFunction1_MCInst1_MC1_n150) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC1_U55 ( .A1(SubCellOutput1[17]), .A2(
        SubCellOutput1[18]), .B1(LED_RoundFunction1_MCInst1_MC1_n144), .B2(
        LED_RoundFunction1_MCInst1_MC1_n143), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n146) );
  INV_X1 LED_RoundFunction1_MCInst1_MC1_U54 ( .A(SubCellOutput1[17]), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n143) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U53 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n142), .B(
        LED_RoundFunction1_MCInst1_MC1_n141), .ZN(
        LED_RoundFunction1_Feedback_27_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U52 ( .A(SubCellOutput1[39]), .B(
        LED_RoundFunction1_MCInst1_MC1_n140), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n141) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U51 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n139), .B(SubCellOutput1[56]), .Z(
        LED_RoundFunction1_MCInst1_MC1_n142) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC1_U50 ( .A1(SubCellOutput1[38]), .A2(
        SubCellOutput1[18]), .B1(LED_RoundFunction1_MCInst1_MC1_n144), .B2(
        LED_RoundFunction1_MCInst1_MC1_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n139) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U49 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n137), .B(
        LED_RoundFunction1_MCInst1_MC1_n136), .ZN(
        LED_RoundFunction1_Feedback_26_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U48 ( .A(SubCellOutput1[36]), .B(
        LED_RoundFunction1_MCInst1_MC1_n135), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n136) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U47 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n134), .B(
        LED_RoundFunction1_MCInst1_MC1_n133), .Z(
        LED_RoundFunction1_MCInst1_MC1_n137) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC1_U46 ( .A1(SubCellOutput1[18]), .A2(
        SubCellOutput1[57]), .B1(LED_RoundFunction1_MCInst1_MC1_n132), .B2(
        LED_RoundFunction1_MCInst1_MC1_n144), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n134) );
  INV_X1 LED_RoundFunction1_MCInst1_MC1_U45 ( .A(SubCellOutput1[18]), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n144) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U44 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n131), .B(
        LED_RoundFunction1_MCInst1_MC1_n151), .ZN(
        LED_RoundFunction1_Feedback_25_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U43 ( .A(SubCellOutput1[59]), .B(
        SubCellOutput1[56]), .ZN(LED_RoundFunction1_MCInst1_MC1_n151) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U42 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n130), .B(
        LED_RoundFunction1_MCInst1_MC1_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n131) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U41 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n128), .B(
        LED_RoundFunction1_MCInst1_MC1_n127), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n130) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U40 ( .A(SubCellOutput1[17]), .B(
        LED_RoundFunction1_MCInst1_MC1_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n127) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U39 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n125), .B(SubCellOutput1[16]), .Z(
        LED_RoundFunction1_MCInst1_MC1_n128) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U38 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n124), .B(
        LED_RoundFunction1_MCInst1_MC1_n123), .ZN(
        LED_RoundFunction1_Feedback_24_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U37 ( .A(SubCellOutput1[12]), .B(
        LED_RoundFunction1_MCInst1_MC1_n122), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n124) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U36 ( .A(SubCellOutput1[14]), .B(
        LED_RoundFunction1_MCInst1_MC1_n122), .ZN(
        LED_RoundFunction1_Feedback_43_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U35 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n135), .B(
        LED_RoundFunction1_MCInst1_MC1_n121), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n122) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U34 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n120), .B(
        LED_RoundFunction1_MCInst1_MC1_n125), .Z(
        LED_RoundFunction1_MCInst1_MC1_n135) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U33 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n119), .B(
        LED_RoundFunction1_MCInst1_MC1_n118), .ZN(
        LED_RoundFunction1_Feedback_42_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U32 ( .A(SubCellOutput1[18]), .B(
        LED_RoundFunction1_MCInst1_MC1_n145), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n118) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U31 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n140), .B(
        LED_RoundFunction1_MCInst1_MC1_n147), .Z(
        LED_RoundFunction1_MCInst1_MC1_n119) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U30 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n126), .B(
        LED_RoundFunction1_MCInst1_MC1_n117), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n140) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U29 ( .A(SubCellOutput1[12]), .B(
        LED_RoundFunction1_MCInst1_MC1_n116), .ZN(
        LED_RoundFunction1_Feedback_41_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U28 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n115), .B(
        LED_RoundFunction1_MCInst1_MC1_n114), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n116) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U27 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n158), .B(SubCellOutput1[57]), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n115) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U26 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n120), .B(
        LED_RoundFunction1_MCInst1_MC1_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n158) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U25 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n113), .B(
        LED_RoundFunction1_MCInst1_MC1_n112), .ZN(
        LED_RoundFunction1_Feedback_40_) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC1_U24 ( .A1(SubCellOutput1[38]), .A2(
        LED_RoundFunction1_MCInst1_MC1_n111), .B1(
        LED_RoundFunction1_MCInst1_MC1_n129), .B2(
        LED_RoundFunction1_MCInst1_MC1_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n112) );
  INV_X1 LED_RoundFunction1_MCInst1_MC1_U23 ( .A(SubCellOutput1[38]), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n138) );
  INV_X1 LED_RoundFunction1_MCInst1_MC1_U22 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n111), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n129) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U21 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n145), .B(
        LED_RoundFunction1_MCInst1_MC1_n154), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n113) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC1_U20 ( .A1(SubCellOutput1[57]), .A2(
        SubCellOutput1[16]), .B1(LED_RoundFunction1_MCInst1_MC1_n110), .B2(
        LED_RoundFunction1_MCInst1_MC1_n132), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n154) );
  INV_X1 LED_RoundFunction1_MCInst1_MC1_U19 ( .A(SubCellOutput1[57]), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n132) );
  INV_X1 LED_RoundFunction1_MCInst1_MC1_U18 ( .A(SubCellOutput1[16]), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n110) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U17 ( .A(SubCellOutput1[15]), .B(
        SubCellOutput1[39]), .Z(LED_RoundFunction1_MCInst1_MC1_n145) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U16 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n111), .B(
        LED_RoundFunction1_MCInst1_MC1_n123), .ZN(
        LED_RoundFunction1_Feedback_59_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U15 ( .A(SubCellOutput1[57]), .B(
        SubCellOutput1[39]), .ZN(LED_RoundFunction1_MCInst1_MC1_n123) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U14 ( .A(SubCellOutput1[18]), .B(
        SubCellOutput1[14]), .Z(LED_RoundFunction1_MCInst1_MC1_n111) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U13 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n120), .B(
        LED_RoundFunction1_MCInst1_MC1_n121), .Z(
        LED_RoundFunction1_Feedback_58_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U12 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n147), .B(SubCellOutput1[56]), .Z(
        LED_RoundFunction1_MCInst1_MC1_n121) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U11 ( .A(SubCellOutput1[13]), .B(
        SubCellOutput1[59]), .Z(LED_RoundFunction1_MCInst1_MC1_n147) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U10 ( .A(SubCellOutput1[38]), .B(
        SubCellOutput1[17]), .Z(LED_RoundFunction1_MCInst1_MC1_n120) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U9 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n117), .B(
        LED_RoundFunction1_MCInst1_MC1_n109), .ZN(
        LED_RoundFunction1_Feedback_57_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U8 ( .A(SubCellOutput1[58]), .B(
        LED_RoundFunction1_MCInst1_MC1_n133), .Z(
        LED_RoundFunction1_MCInst1_MC1_n109) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U7 ( .A(SubCellOutput1[15]), .B(
        SubCellOutput1[59]), .Z(LED_RoundFunction1_MCInst1_MC1_n133) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U6 ( .A(
        LED_RoundFunction1_MCInst1_MC1_n159), .B(
        LED_RoundFunction1_MCInst1_MC1_n125), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n117) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U5 ( .A(SubCellOutput1[19]), .B(
        SubCellOutput1[37]), .Z(LED_RoundFunction1_MCInst1_MC1_n125) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U4 ( .A(SubCellOutput1[12]), .B(
        SubCellOutput1[16]), .Z(LED_RoundFunction1_MCInst1_MC1_n159) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U3 ( .A(SubCellOutput1[15]), .B(
        LED_RoundFunction1_MCInst1_MC1_n114), .ZN(
        LED_RoundFunction1_Feedback_56_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC1_U2 ( .A(SubCellOutput1[19]), .B(
        LED_RoundFunction1_MCInst1_MC1_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC1_n114) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC1_U1 ( .A(SubCellOutput1[58]), .B(
        SubCellOutput1[36]), .Z(LED_RoundFunction1_MCInst1_MC1_n126) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U68 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n160), .B(
        LED_RoundFunction1_MCInst1_MC2_n159), .ZN(
        LED_RoundFunction1_Feedback_7_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U67 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n158), .B(SubCellOutput1[54]), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n160) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U66 ( .A(SubCellOutput1[11]), .B(
        LED_RoundFunction1_MCInst1_MC2_n157), .Z(
        LED_RoundFunction1_Feedback_6_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U65 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n156), .B(
        LED_RoundFunction1_MCInst1_MC2_n155), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n157) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U64 ( .A(SubCellOutput1[29]), .B(
        SubCellOutput1[9]), .ZN(LED_RoundFunction1_MCInst1_MC2_n155) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U63 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n154), .B(SubCellOutput1[33]), .Z(
        LED_RoundFunction1_MCInst1_MC2_n156) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U62 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n153), .B(
        LED_RoundFunction1_MCInst1_MC2_n152), .ZN(
        LED_RoundFunction1_Feedback_5_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U61 ( .A(SubCellOutput1[10]), .B(
        SubCellOutput1[32]), .ZN(LED_RoundFunction1_MCInst1_MC2_n152) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U60 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n151), .B(
        LED_RoundFunction1_MCInst1_MC2_n150), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n153) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U59 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n149), .B(
        LED_RoundFunction1_MCInst1_MC2_n148), .ZN(
        LED_RoundFunction1_Feedback_4_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U58 ( .A(SubCellOutput1[31]), .B(
        LED_RoundFunction1_MCInst1_MC2_n147), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n148) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U57 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n146), .B(
        LED_RoundFunction1_MCInst1_MC2_n150), .Z(
        LED_RoundFunction1_MCInst1_MC2_n149) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U56 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n145), .B(
        LED_RoundFunction1_MCInst1_MC2_n159), .Z(
        LED_RoundFunction1_MCInst1_MC2_n150) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC2_U55 ( .A1(SubCellOutput1[29]), .A2(
        SubCellOutput1[30]), .B1(LED_RoundFunction1_MCInst1_MC2_n144), .B2(
        LED_RoundFunction1_MCInst1_MC2_n143), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n146) );
  INV_X1 LED_RoundFunction1_MCInst1_MC2_U54 ( .A(SubCellOutput1[29]), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n143) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U53 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n142), .B(
        LED_RoundFunction1_MCInst1_MC2_n141), .ZN(
        LED_RoundFunction1_Feedback_23_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U52 ( .A(SubCellOutput1[35]), .B(
        LED_RoundFunction1_MCInst1_MC2_n140), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n141) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U51 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n139), .B(SubCellOutput1[52]), .Z(
        LED_RoundFunction1_MCInst1_MC2_n142) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC2_U50 ( .A1(SubCellOutput1[34]), .A2(
        SubCellOutput1[30]), .B1(LED_RoundFunction1_MCInst1_MC2_n144), .B2(
        LED_RoundFunction1_MCInst1_MC2_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n139) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U49 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n137), .B(
        LED_RoundFunction1_MCInst1_MC2_n136), .ZN(
        LED_RoundFunction1_Feedback_22_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U48 ( .A(SubCellOutput1[32]), .B(
        LED_RoundFunction1_MCInst1_MC2_n135), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n136) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U47 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n134), .B(
        LED_RoundFunction1_MCInst1_MC2_n133), .Z(
        LED_RoundFunction1_MCInst1_MC2_n137) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC2_U46 ( .A1(SubCellOutput1[30]), .A2(
        SubCellOutput1[53]), .B1(LED_RoundFunction1_MCInst1_MC2_n132), .B2(
        LED_RoundFunction1_MCInst1_MC2_n144), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n134) );
  INV_X1 LED_RoundFunction1_MCInst1_MC2_U45 ( .A(SubCellOutput1[30]), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n144) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U44 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n131), .B(
        LED_RoundFunction1_MCInst1_MC2_n151), .ZN(
        LED_RoundFunction1_Feedback_21_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U43 ( .A(SubCellOutput1[55]), .B(
        SubCellOutput1[52]), .ZN(LED_RoundFunction1_MCInst1_MC2_n151) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U42 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n130), .B(
        LED_RoundFunction1_MCInst1_MC2_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n131) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U41 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n128), .B(
        LED_RoundFunction1_MCInst1_MC2_n127), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n130) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U40 ( .A(SubCellOutput1[29]), .B(
        LED_RoundFunction1_MCInst1_MC2_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n127) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U39 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n125), .B(SubCellOutput1[28]), .Z(
        LED_RoundFunction1_MCInst1_MC2_n128) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U38 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n124), .B(
        LED_RoundFunction1_MCInst1_MC2_n123), .ZN(
        LED_RoundFunction1_Feedback_20_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U37 ( .A(SubCellOutput1[8]), .B(
        LED_RoundFunction1_MCInst1_MC2_n122), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n124) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U36 ( .A(SubCellOutput1[10]), .B(
        LED_RoundFunction1_MCInst1_MC2_n122), .ZN(
        LED_RoundFunction1_Feedback_39_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U35 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n135), .B(
        LED_RoundFunction1_MCInst1_MC2_n121), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n122) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U34 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n120), .B(
        LED_RoundFunction1_MCInst1_MC2_n125), .Z(
        LED_RoundFunction1_MCInst1_MC2_n135) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U33 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n119), .B(
        LED_RoundFunction1_MCInst1_MC2_n118), .ZN(
        LED_RoundFunction1_Feedback_38_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U32 ( .A(SubCellOutput1[30]), .B(
        LED_RoundFunction1_MCInst1_MC2_n145), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n118) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U31 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n140), .B(
        LED_RoundFunction1_MCInst1_MC2_n147), .Z(
        LED_RoundFunction1_MCInst1_MC2_n119) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U30 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n126), .B(
        LED_RoundFunction1_MCInst1_MC2_n117), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n140) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U29 ( .A(SubCellOutput1[8]), .B(
        LED_RoundFunction1_MCInst1_MC2_n116), .ZN(
        LED_RoundFunction1_Feedback_37_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U28 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n115), .B(
        LED_RoundFunction1_MCInst1_MC2_n114), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n116) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U27 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n158), .B(SubCellOutput1[53]), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n115) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U26 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n120), .B(
        LED_RoundFunction1_MCInst1_MC2_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n158) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U25 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n113), .B(
        LED_RoundFunction1_MCInst1_MC2_n112), .ZN(
        LED_RoundFunction1_Feedback_36_) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC2_U24 ( .A1(SubCellOutput1[34]), .A2(
        LED_RoundFunction1_MCInst1_MC2_n111), .B1(
        LED_RoundFunction1_MCInst1_MC2_n129), .B2(
        LED_RoundFunction1_MCInst1_MC2_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n112) );
  INV_X1 LED_RoundFunction1_MCInst1_MC2_U23 ( .A(SubCellOutput1[34]), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n138) );
  INV_X1 LED_RoundFunction1_MCInst1_MC2_U22 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n111), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n129) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U21 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n145), .B(
        LED_RoundFunction1_MCInst1_MC2_n154), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n113) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC2_U20 ( .A1(SubCellOutput1[53]), .A2(
        SubCellOutput1[28]), .B1(LED_RoundFunction1_MCInst1_MC2_n110), .B2(
        LED_RoundFunction1_MCInst1_MC2_n132), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n154) );
  INV_X1 LED_RoundFunction1_MCInst1_MC2_U19 ( .A(SubCellOutput1[53]), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n132) );
  INV_X1 LED_RoundFunction1_MCInst1_MC2_U18 ( .A(SubCellOutput1[28]), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n110) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U17 ( .A(SubCellOutput1[11]), .B(
        SubCellOutput1[35]), .Z(LED_RoundFunction1_MCInst1_MC2_n145) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U16 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n111), .B(
        LED_RoundFunction1_MCInst1_MC2_n123), .ZN(
        LED_RoundFunction1_Feedback_55_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U15 ( .A(SubCellOutput1[53]), .B(
        SubCellOutput1[35]), .ZN(LED_RoundFunction1_MCInst1_MC2_n123) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U14 ( .A(SubCellOutput1[30]), .B(
        SubCellOutput1[10]), .Z(LED_RoundFunction1_MCInst1_MC2_n111) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U13 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n120), .B(
        LED_RoundFunction1_MCInst1_MC2_n121), .Z(
        LED_RoundFunction1_Feedback_54_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U12 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n147), .B(SubCellOutput1[52]), .Z(
        LED_RoundFunction1_MCInst1_MC2_n121) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U11 ( .A(SubCellOutput1[9]), .B(
        SubCellOutput1[55]), .Z(LED_RoundFunction1_MCInst1_MC2_n147) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U10 ( .A(SubCellOutput1[34]), .B(
        SubCellOutput1[29]), .Z(LED_RoundFunction1_MCInst1_MC2_n120) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U9 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n117), .B(
        LED_RoundFunction1_MCInst1_MC2_n109), .ZN(
        LED_RoundFunction1_Feedback_53_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U8 ( .A(SubCellOutput1[54]), .B(
        LED_RoundFunction1_MCInst1_MC2_n133), .Z(
        LED_RoundFunction1_MCInst1_MC2_n109) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U7 ( .A(SubCellOutput1[11]), .B(
        SubCellOutput1[55]), .Z(LED_RoundFunction1_MCInst1_MC2_n133) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U6 ( .A(
        LED_RoundFunction1_MCInst1_MC2_n159), .B(
        LED_RoundFunction1_MCInst1_MC2_n125), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n117) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U5 ( .A(SubCellOutput1[31]), .B(
        SubCellOutput1[33]), .Z(LED_RoundFunction1_MCInst1_MC2_n125) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U4 ( .A(SubCellOutput1[8]), .B(
        SubCellOutput1[28]), .Z(LED_RoundFunction1_MCInst1_MC2_n159) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U3 ( .A(SubCellOutput1[11]), .B(
        LED_RoundFunction1_MCInst1_MC2_n114), .ZN(
        LED_RoundFunction1_Feedback_52_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC2_U2 ( .A(SubCellOutput1[31]), .B(
        LED_RoundFunction1_MCInst1_MC2_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC2_n114) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC2_U1 ( .A(SubCellOutput1[54]), .B(
        SubCellOutput1[32]), .Z(LED_RoundFunction1_MCInst1_MC2_n126) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U68 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n160), .B(
        LED_RoundFunction1_MCInst1_MC3_n159), .ZN(
        LED_RoundFunction1_Feedback_3_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U67 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n158), .B(SubCellOutput1[50]), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n160) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U66 ( .A(SubCellOutput1[7]), .B(
        LED_RoundFunction1_MCInst1_MC3_n157), .Z(
        LED_RoundFunction1_Feedback_2_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U65 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n156), .B(
        LED_RoundFunction1_MCInst1_MC3_n155), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n157) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U64 ( .A(SubCellOutput1[25]), .B(
        SubCellOutput1[5]), .ZN(LED_RoundFunction1_MCInst1_MC3_n155) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U63 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n154), .B(SubCellOutput1[45]), .Z(
        LED_RoundFunction1_MCInst1_MC3_n156) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U62 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n153), .B(
        LED_RoundFunction1_MCInst1_MC3_n152), .ZN(
        LED_RoundFunction1_Feedback_1_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U61 ( .A(SubCellOutput1[6]), .B(
        SubCellOutput1[44]), .ZN(LED_RoundFunction1_MCInst1_MC3_n152) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U60 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n151), .B(
        LED_RoundFunction1_MCInst1_MC3_n150), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n153) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U59 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n149), .B(
        LED_RoundFunction1_MCInst1_MC3_n148), .ZN(
        LED_RoundFunction1_Feedback_0_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U58 ( .A(SubCellOutput1[27]), .B(
        LED_RoundFunction1_MCInst1_MC3_n147), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n148) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U57 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n146), .B(
        LED_RoundFunction1_MCInst1_MC3_n150), .Z(
        LED_RoundFunction1_MCInst1_MC3_n149) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U56 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n145), .B(
        LED_RoundFunction1_MCInst1_MC3_n159), .Z(
        LED_RoundFunction1_MCInst1_MC3_n150) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC3_U55 ( .A1(SubCellOutput1[25]), .A2(
        SubCellOutput1[26]), .B1(LED_RoundFunction1_MCInst1_MC3_n144), .B2(
        LED_RoundFunction1_MCInst1_MC3_n143), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n146) );
  INV_X1 LED_RoundFunction1_MCInst1_MC3_U54 ( .A(SubCellOutput1[25]), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n143) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U53 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n142), .B(
        LED_RoundFunction1_MCInst1_MC3_n141), .ZN(
        LED_RoundFunction1_Feedback_19_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U52 ( .A(SubCellOutput1[47]), .B(
        LED_RoundFunction1_MCInst1_MC3_n140), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n141) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U51 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n139), .B(SubCellOutput1[48]), .Z(
        LED_RoundFunction1_MCInst1_MC3_n142) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC3_U50 ( .A1(SubCellOutput1[46]), .A2(
        SubCellOutput1[26]), .B1(LED_RoundFunction1_MCInst1_MC3_n144), .B2(
        LED_RoundFunction1_MCInst1_MC3_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n139) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U49 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n137), .B(
        LED_RoundFunction1_MCInst1_MC3_n136), .ZN(
        LED_RoundFunction1_Feedback_18_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U48 ( .A(SubCellOutput1[44]), .B(
        LED_RoundFunction1_MCInst1_MC3_n135), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n136) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U47 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n134), .B(
        LED_RoundFunction1_MCInst1_MC3_n133), .Z(
        LED_RoundFunction1_MCInst1_MC3_n137) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC3_U46 ( .A1(SubCellOutput1[26]), .A2(
        SubCellOutput1[49]), .B1(LED_RoundFunction1_MCInst1_MC3_n132), .B2(
        LED_RoundFunction1_MCInst1_MC3_n144), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n134) );
  INV_X1 LED_RoundFunction1_MCInst1_MC3_U45 ( .A(SubCellOutput1[26]), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n144) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U44 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n131), .B(
        LED_RoundFunction1_MCInst1_MC3_n151), .ZN(
        LED_RoundFunction1_Feedback_17_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U43 ( .A(SubCellOutput1[51]), .B(
        SubCellOutput1[48]), .ZN(LED_RoundFunction1_MCInst1_MC3_n151) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U42 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n130), .B(
        LED_RoundFunction1_MCInst1_MC3_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n131) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U41 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n128), .B(
        LED_RoundFunction1_MCInst1_MC3_n127), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n130) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U40 ( .A(SubCellOutput1[25]), .B(
        LED_RoundFunction1_MCInst1_MC3_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n127) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U39 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n125), .B(SubCellOutput1[24]), .Z(
        LED_RoundFunction1_MCInst1_MC3_n128) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U38 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n124), .B(
        LED_RoundFunction1_MCInst1_MC3_n123), .ZN(
        LED_RoundFunction1_Feedback_16_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U37 ( .A(SubCellOutput1[4]), .B(
        LED_RoundFunction1_MCInst1_MC3_n122), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n124) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U36 ( .A(SubCellOutput1[6]), .B(
        LED_RoundFunction1_MCInst1_MC3_n122), .ZN(
        LED_RoundFunction1_Feedback_35_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U35 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n135), .B(
        LED_RoundFunction1_MCInst1_MC3_n121), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n122) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U34 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n120), .B(
        LED_RoundFunction1_MCInst1_MC3_n125), .Z(
        LED_RoundFunction1_MCInst1_MC3_n135) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U33 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n119), .B(
        LED_RoundFunction1_MCInst1_MC3_n118), .ZN(
        LED_RoundFunction1_Feedback_34_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U32 ( .A(SubCellOutput1[26]), .B(
        LED_RoundFunction1_MCInst1_MC3_n145), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n118) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U31 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n140), .B(
        LED_RoundFunction1_MCInst1_MC3_n147), .Z(
        LED_RoundFunction1_MCInst1_MC3_n119) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U30 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n126), .B(
        LED_RoundFunction1_MCInst1_MC3_n117), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n140) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U29 ( .A(SubCellOutput1[4]), .B(
        LED_RoundFunction1_MCInst1_MC3_n116), .ZN(
        LED_RoundFunction1_Feedback_33_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U28 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n115), .B(
        LED_RoundFunction1_MCInst1_MC3_n114), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n116) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U27 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n158), .B(SubCellOutput1[49]), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n115) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U26 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n120), .B(
        LED_RoundFunction1_MCInst1_MC3_n129), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n158) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U25 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n113), .B(
        LED_RoundFunction1_MCInst1_MC3_n112), .ZN(
        LED_RoundFunction1_Feedback_32_) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC3_U24 ( .A1(SubCellOutput1[46]), .A2(
        LED_RoundFunction1_MCInst1_MC3_n111), .B1(
        LED_RoundFunction1_MCInst1_MC3_n129), .B2(
        LED_RoundFunction1_MCInst1_MC3_n138), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n112) );
  INV_X1 LED_RoundFunction1_MCInst1_MC3_U23 ( .A(SubCellOutput1[46]), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n138) );
  INV_X1 LED_RoundFunction1_MCInst1_MC3_U22 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n111), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n129) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U21 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n145), .B(
        LED_RoundFunction1_MCInst1_MC3_n154), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n113) );
  AOI22_X1 LED_RoundFunction1_MCInst1_MC3_U20 ( .A1(SubCellOutput1[49]), .A2(
        SubCellOutput1[24]), .B1(LED_RoundFunction1_MCInst1_MC3_n110), .B2(
        LED_RoundFunction1_MCInst1_MC3_n132), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n154) );
  INV_X1 LED_RoundFunction1_MCInst1_MC3_U19 ( .A(SubCellOutput1[49]), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n132) );
  INV_X1 LED_RoundFunction1_MCInst1_MC3_U18 ( .A(SubCellOutput1[24]), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n110) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U17 ( .A(SubCellOutput1[7]), .B(
        SubCellOutput1[47]), .Z(LED_RoundFunction1_MCInst1_MC3_n145) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U16 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n111), .B(
        LED_RoundFunction1_MCInst1_MC3_n123), .ZN(
        LED_RoundFunction1_Feedback_51_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U15 ( .A(SubCellOutput1[49]), .B(
        SubCellOutput1[47]), .ZN(LED_RoundFunction1_MCInst1_MC3_n123) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U14 ( .A(SubCellOutput1[26]), .B(
        SubCellOutput1[6]), .Z(LED_RoundFunction1_MCInst1_MC3_n111) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U13 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n120), .B(
        LED_RoundFunction1_MCInst1_MC3_n121), .Z(
        LED_RoundFunction1_Feedback_50_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U12 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n147), .B(SubCellOutput1[48]), .Z(
        LED_RoundFunction1_MCInst1_MC3_n121) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U11 ( .A(SubCellOutput1[5]), .B(
        SubCellOutput1[51]), .Z(LED_RoundFunction1_MCInst1_MC3_n147) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U10 ( .A(SubCellOutput1[46]), .B(
        SubCellOutput1[25]), .Z(LED_RoundFunction1_MCInst1_MC3_n120) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U9 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n117), .B(
        LED_RoundFunction1_MCInst1_MC3_n109), .ZN(
        LED_RoundFunction1_Feedback_49_) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U8 ( .A(SubCellOutput1[50]), .B(
        LED_RoundFunction1_MCInst1_MC3_n133), .Z(
        LED_RoundFunction1_MCInst1_MC3_n109) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U7 ( .A(SubCellOutput1[7]), .B(
        SubCellOutput1[51]), .Z(LED_RoundFunction1_MCInst1_MC3_n133) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U6 ( .A(
        LED_RoundFunction1_MCInst1_MC3_n159), .B(
        LED_RoundFunction1_MCInst1_MC3_n125), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n117) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U5 ( .A(SubCellOutput1[27]), .B(
        SubCellOutput1[45]), .Z(LED_RoundFunction1_MCInst1_MC3_n125) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U4 ( .A(SubCellOutput1[4]), .B(
        SubCellOutput1[24]), .Z(LED_RoundFunction1_MCInst1_MC3_n159) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U3 ( .A(SubCellOutput1[7]), .B(
        LED_RoundFunction1_MCInst1_MC3_n114), .ZN(
        LED_RoundFunction1_Feedback_48_) );
  XNOR2_X1 LED_RoundFunction1_MCInst1_MC3_U2 ( .A(SubCellOutput1[27]), .B(
        LED_RoundFunction1_MCInst1_MC3_n126), .ZN(
        LED_RoundFunction1_MCInst1_MC3_n114) );
  XOR2_X1 LED_RoundFunction1_MCInst1_MC3_U1 ( .A(SubCellOutput1[50]), .B(
        SubCellOutput1[44]), .Z(LED_RoundFunction1_MCInst1_MC3_n126) );
  AOI22_X1 LED_RoundFunction2_U412 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n836), .B1(LED_RoundFunction2_n835), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U411 ( .A1(rst), .A2(Plaintext2[0]), .B1(
        LED_RoundFunction2_Feedback_0_), .B2(LED_RoundFunction2_n564), .ZN(
        LED_RoundFunction2_n835) );
  INV_X1 LED_RoundFunction2_U410 ( .A(Ciphertext2[0]), .ZN(
        LED_RoundFunction2_n836) );
  AOI22_X1 LED_RoundFunction2_U409 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n834), .B1(LED_RoundFunction2_n833), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U408 ( .A1(rst), .A2(Plaintext2[1]), .B1(
        LED_RoundFunction2_Feedback_1_), .B2(LED_RoundFunction2_n568), .ZN(
        LED_RoundFunction2_n833) );
  INV_X1 LED_RoundFunction2_U407 ( .A(Ciphertext2[1]), .ZN(
        LED_RoundFunction2_n834) );
  AOI22_X1 LED_RoundFunction2_U406 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n832), .B1(LED_RoundFunction2_n831), .B2(
        LED_RoundFunction2_n561), .ZN(SubCellInput2[2]) );
  AOI22_X1 LED_RoundFunction2_U405 ( .A1(rst), .A2(Plaintext2[2]), .B1(
        LED_RoundFunction2_Feedback_2_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n831) );
  INV_X1 LED_RoundFunction2_U404 ( .A(Ciphertext2[2]), .ZN(
        LED_RoundFunction2_n832) );
  AOI22_X1 LED_RoundFunction2_U403 ( .A1(LED_RoundFunction2_n556), .A2(
        LED_RoundFunction2_n830), .B1(LED_RoundFunction2_n829), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U402 ( .A1(rst), .A2(Plaintext2[3]), .B1(
        LED_RoundFunction2_Feedback_3_), .B2(LED_RoundFunction2_n568), .ZN(
        LED_RoundFunction2_n829) );
  INV_X1 LED_RoundFunction2_U401 ( .A(Ciphertext2[3]), .ZN(
        LED_RoundFunction2_n830) );
  AOI22_X1 LED_RoundFunction2_U400 ( .A1(LED_RoundFunction2_n557), .A2(
        LED_RoundFunction2_n828), .B1(LED_RoundFunction2_n827), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U399 ( .A1(rst), .A2(Plaintext2[4]), .B1(
        LED_RoundFunction2_Feedback_4_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n827) );
  INV_X1 LED_RoundFunction2_U398 ( .A(Ciphertext2[4]), .ZN(
        LED_RoundFunction2_n828) );
  AOI22_X1 LED_RoundFunction2_U397 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n826), .B1(LED_RoundFunction2_n825), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U396 ( .A1(rst), .A2(Plaintext2[5]), .B1(
        LED_RoundFunction2_Feedback_5_), .B2(LED_RoundFunction2_n568), .ZN(
        LED_RoundFunction2_n825) );
  INV_X1 LED_RoundFunction2_U395 ( .A(Ciphertext2[5]), .ZN(
        LED_RoundFunction2_n826) );
  AOI22_X1 LED_RoundFunction2_U394 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n824), .B1(LED_RoundFunction2_n823), .B2(
        LED_RoundFunction2_n560), .ZN(SubCellInput2[6]) );
  AOI22_X1 LED_RoundFunction2_U393 ( .A1(rst), .A2(Plaintext2[6]), .B1(
        LED_RoundFunction2_Feedback_6_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n823) );
  INV_X1 LED_RoundFunction2_U392 ( .A(Ciphertext2[6]), .ZN(
        LED_RoundFunction2_n824) );
  AOI22_X1 LED_RoundFunction2_U391 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n822), .B1(LED_RoundFunction2_n821), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U390 ( .A1(rst), .A2(Plaintext2[7]), .B1(
        LED_RoundFunction2_Feedback_7_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n821) );
  INV_X1 LED_RoundFunction2_U389 ( .A(Ciphertext2[7]), .ZN(
        LED_RoundFunction2_n822) );
  AOI22_X1 LED_RoundFunction2_U388 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n820), .B1(LED_RoundFunction2_n819), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U387 ( .A1(rst), .A2(Plaintext2[11]), .B1(
        LED_RoundFunction2_Feedback_11_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n819) );
  INV_X1 LED_RoundFunction2_U386 ( .A(Ciphertext2[11]), .ZN(
        LED_RoundFunction2_n820) );
  AOI22_X1 LED_RoundFunction2_U385 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n818), .B1(LED_RoundFunction2_n817), .B2(
        LED_RoundFunction2_n561), .ZN(SubCellInput2[14]) );
  AOI22_X1 LED_RoundFunction2_U384 ( .A1(rst), .A2(Plaintext2[14]), .B1(
        LED_RoundFunction2_Feedback_14_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n817) );
  INV_X1 LED_RoundFunction2_U383 ( .A(Ciphertext2[14]), .ZN(
        LED_RoundFunction2_n818) );
  AOI22_X1 LED_RoundFunction2_U382 ( .A1(LED_RoundFunction2_n556), .A2(
        LED_RoundFunction2_n816), .B1(LED_RoundFunction2_n815), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U381 ( .A1(rst), .A2(Plaintext2[15]), .B1(
        LED_RoundFunction2_Feedback_15_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n815) );
  INV_X1 LED_RoundFunction2_U380 ( .A(Ciphertext2[15]), .ZN(
        LED_RoundFunction2_n816) );
  AOI22_X1 LED_RoundFunction2_U379 ( .A1(LED_RoundFunction2_n557), .A2(
        LED_RoundFunction2_n814), .B1(LED_RoundFunction2_n813), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U378 ( .A1(rst), .A2(Plaintext2[16]), .B1(
        LED_RoundFunction2_Feedback_16_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n813) );
  INV_X1 LED_RoundFunction2_U377 ( .A(Ciphertext2[16]), .ZN(
        LED_RoundFunction2_n814) );
  AOI22_X1 LED_RoundFunction2_U376 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n812), .B1(LED_RoundFunction2_n811), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U375 ( .A1(rst), .A2(Plaintext2[17]), .B1(
        LED_RoundFunction2_Feedback_17_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n811) );
  INV_X1 LED_RoundFunction2_U374 ( .A(Ciphertext2[17]), .ZN(
        LED_RoundFunction2_n812) );
  AOI22_X1 LED_RoundFunction2_U373 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n810), .B1(LED_RoundFunction2_n809), .B2(
        LED_RoundFunction2_n560), .ZN(SubCellInput2[18]) );
  AOI22_X1 LED_RoundFunction2_U372 ( .A1(rst), .A2(Plaintext2[18]), .B1(
        LED_RoundFunction2_Feedback_18_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n809) );
  INV_X1 LED_RoundFunction2_U371 ( .A(Ciphertext2[18]), .ZN(
        LED_RoundFunction2_n810) );
  AOI22_X1 LED_RoundFunction2_U370 ( .A1(LED_RoundFunction2_n556), .A2(
        LED_RoundFunction2_n808), .B1(LED_RoundFunction2_n807), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U369 ( .A1(rst), .A2(Plaintext2[19]), .B1(
        LED_RoundFunction2_Feedback_19_), .B2(LED_RoundFunction2_n568), .ZN(
        LED_RoundFunction2_n807) );
  INV_X1 LED_RoundFunction2_U368 ( .A(Ciphertext2[19]), .ZN(
        LED_RoundFunction2_n808) );
  AOI22_X1 LED_RoundFunction2_U367 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n806), .B1(LED_RoundFunction2_n805), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U366 ( .A1(rst), .A2(Plaintext2[20]), .B1(
        LED_RoundFunction2_Feedback_20_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n805) );
  INV_X1 LED_RoundFunction2_U365 ( .A(Ciphertext2[20]), .ZN(
        LED_RoundFunction2_n806) );
  AOI22_X1 LED_RoundFunction2_U364 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n804), .B1(LED_RoundFunction2_n803), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U363 ( .A1(rst), .A2(Plaintext2[21]), .B1(
        LED_RoundFunction2_Feedback_21_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n803) );
  INV_X1 LED_RoundFunction2_U362 ( .A(Ciphertext2[21]), .ZN(
        LED_RoundFunction2_n804) );
  AOI22_X1 LED_RoundFunction2_U361 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n802), .B1(LED_RoundFunction2_n801), .B2(
        LED_RoundFunction2_n561), .ZN(SubCellInput2[22]) );
  AOI22_X1 LED_RoundFunction2_U360 ( .A1(rst), .A2(Plaintext2[22]), .B1(
        LED_RoundFunction2_Feedback_22_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n801) );
  INV_X1 LED_RoundFunction2_U359 ( .A(Ciphertext2[22]), .ZN(
        LED_RoundFunction2_n802) );
  AOI22_X1 LED_RoundFunction2_U358 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n800), .B1(LED_RoundFunction2_n799), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U357 ( .A1(rst), .A2(Plaintext2[23]), .B1(
        LED_RoundFunction2_Feedback_23_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n799) );
  INV_X1 LED_RoundFunction2_U356 ( .A(Ciphertext2[23]), .ZN(
        LED_RoundFunction2_n800) );
  AOI22_X1 LED_RoundFunction2_U355 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n798), .B1(LED_RoundFunction2_n797), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U354 ( .A1(rst), .A2(Plaintext2[27]), .B1(
        LED_RoundFunction2_Feedback_27_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n797) );
  INV_X1 LED_RoundFunction2_U353 ( .A(Ciphertext2[27]), .ZN(
        LED_RoundFunction2_n798) );
  AOI22_X1 LED_RoundFunction2_U352 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n796), .B1(LED_RoundFunction2_n795), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U351 ( .A1(rst), .A2(Plaintext2[28]), .B1(
        LED_RoundFunction2_Feedback_28_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n795) );
  INV_X1 LED_RoundFunction2_U350 ( .A(Ciphertext2[28]), .ZN(
        LED_RoundFunction2_n796) );
  AOI22_X1 LED_RoundFunction2_U349 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n794), .B1(LED_RoundFunction2_n793), .B2(
        LED_RoundFunction2_n560), .ZN(SubCellInput2[30]) );
  AOI22_X1 LED_RoundFunction2_U348 ( .A1(rst), .A2(Plaintext2[30]), .B1(
        LED_RoundFunction2_Feedback_30_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n793) );
  INV_X1 LED_RoundFunction2_U347 ( .A(Ciphertext2[30]), .ZN(
        LED_RoundFunction2_n794) );
  AOI22_X1 LED_RoundFunction2_U346 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n792), .B1(LED_RoundFunction2_n791), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U345 ( .A1(rst), .A2(Plaintext2[31]), .B1(
        LED_RoundFunction2_Feedback_31_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n791) );
  INV_X1 LED_RoundFunction2_U344 ( .A(Ciphertext2[31]), .ZN(
        LED_RoundFunction2_n792) );
  AOI22_X1 LED_RoundFunction2_U343 ( .A1(LED_RoundFunction2_n556), .A2(
        LED_RoundFunction2_n790), .B1(LED_RoundFunction2_n789), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U342 ( .A1(rst), .A2(Plaintext2[32]), .B1(
        LED_RoundFunction2_Feedback_32_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n789) );
  INV_X1 LED_RoundFunction2_U341 ( .A(Ciphertext2[32]), .ZN(
        LED_RoundFunction2_n790) );
  AOI22_X1 LED_RoundFunction2_U340 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n788), .B1(LED_RoundFunction2_n787), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U339 ( .A1(rst), .A2(Plaintext2[33]), .B1(
        LED_RoundFunction2_Feedback_33_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n787) );
  INV_X1 LED_RoundFunction2_U338 ( .A(Ciphertext2[33]), .ZN(
        LED_RoundFunction2_n788) );
  AOI22_X1 LED_RoundFunction2_U337 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n786), .B1(LED_RoundFunction2_n785), .B2(
        LED_RoundFunction2_n561), .ZN(SubCellInput2[34]) );
  AOI22_X1 LED_RoundFunction2_U336 ( .A1(rst), .A2(Plaintext2[34]), .B1(
        LED_RoundFunction2_Feedback_34_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n785) );
  INV_X1 LED_RoundFunction2_U335 ( .A(Ciphertext2[34]), .ZN(
        LED_RoundFunction2_n786) );
  AOI22_X1 LED_RoundFunction2_U334 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n784), .B1(LED_RoundFunction2_n783), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U333 ( .A1(rst), .A2(Plaintext2[35]), .B1(
        LED_RoundFunction2_Feedback_35_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n783) );
  INV_X1 LED_RoundFunction2_U332 ( .A(Ciphertext2[35]), .ZN(
        LED_RoundFunction2_n784) );
  AOI22_X1 LED_RoundFunction2_U331 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n782), .B1(LED_RoundFunction2_n781), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U330 ( .A1(rst), .A2(Plaintext2[36]), .B1(
        LED_RoundFunction2_Feedback_36_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n781) );
  INV_X1 LED_RoundFunction2_U329 ( .A(Ciphertext2[36]), .ZN(
        LED_RoundFunction2_n782) );
  AOI22_X1 LED_RoundFunction2_U328 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n780), .B1(LED_RoundFunction2_n779), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U327 ( .A1(rst), .A2(Plaintext2[37]), .B1(
        LED_RoundFunction2_Feedback_37_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n779) );
  INV_X1 LED_RoundFunction2_U326 ( .A(Ciphertext2[37]), .ZN(
        LED_RoundFunction2_n780) );
  AOI22_X1 LED_RoundFunction2_U325 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n778), .B1(LED_RoundFunction2_n777), .B2(
        LED_RoundFunction2_n561), .ZN(SubCellInput2[38]) );
  AOI22_X1 LED_RoundFunction2_U324 ( .A1(rst), .A2(Plaintext2[38]), .B1(
        LED_RoundFunction2_Feedback_38_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n777) );
  INV_X1 LED_RoundFunction2_U323 ( .A(Ciphertext2[38]), .ZN(
        LED_RoundFunction2_n778) );
  AOI22_X1 LED_RoundFunction2_U322 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n776), .B1(LED_RoundFunction2_n775), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U321 ( .A1(rst), .A2(Plaintext2[39]), .B1(
        LED_RoundFunction2_Feedback_39_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n775) );
  INV_X1 LED_RoundFunction2_U320 ( .A(Ciphertext2[39]), .ZN(
        LED_RoundFunction2_n776) );
  AOI22_X1 LED_RoundFunction2_U319 ( .A1(LED_RoundFunction2_n557), .A2(
        LED_RoundFunction2_n774), .B1(LED_RoundFunction2_n773), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U318 ( .A1(rst), .A2(Plaintext2[43]), .B1(
        LED_RoundFunction2_Feedback_43_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n773) );
  INV_X1 LED_RoundFunction2_U317 ( .A(Ciphertext2[43]), .ZN(
        LED_RoundFunction2_n774) );
  AOI22_X1 LED_RoundFunction2_U316 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n772), .B1(LED_RoundFunction2_n771), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U315 ( .A1(rst), .A2(Plaintext2[45]), .B1(
        LED_RoundFunction2_Feedback_45_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n771) );
  INV_X1 LED_RoundFunction2_U314 ( .A(Ciphertext2[45]), .ZN(
        LED_RoundFunction2_n772) );
  AOI22_X1 LED_RoundFunction2_U313 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n770), .B1(LED_RoundFunction2_n769), .B2(
        LED_RoundFunction2_n561), .ZN(SubCellInput2[46]) );
  AOI22_X1 LED_RoundFunction2_U312 ( .A1(rst), .A2(Plaintext2[46]), .B1(
        LED_RoundFunction2_Feedback_46_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n769) );
  INV_X1 LED_RoundFunction2_U311 ( .A(Ciphertext2[46]), .ZN(
        LED_RoundFunction2_n770) );
  AOI22_X1 LED_RoundFunction2_U310 ( .A1(LED_RoundFunction2_n557), .A2(
        LED_RoundFunction2_n768), .B1(LED_RoundFunction2_n767), .B2(
        LED_RoundFunction2_n561), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U309 ( .A1(rst), .A2(Plaintext2[48]), .B1(
        LED_RoundFunction2_Feedback_48_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n767) );
  INV_X1 LED_RoundFunction2_U308 ( .A(Ciphertext2[48]), .ZN(
        LED_RoundFunction2_n768) );
  AOI22_X1 LED_RoundFunction2_U307 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n766), .B1(LED_RoundFunction2_n765), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U306 ( .A1(rst), .A2(Plaintext2[49]), .B1(
        LED_RoundFunction2_Feedback_49_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n765) );
  INV_X1 LED_RoundFunction2_U305 ( .A(Ciphertext2[49]), .ZN(
        LED_RoundFunction2_n766) );
  AOI22_X1 LED_RoundFunction2_U304 ( .A1(LED_RoundFunction2_n558), .A2(
        LED_RoundFunction2_n764), .B1(LED_RoundFunction2_n763), .B2(
        LED_RoundFunction2_n560), .ZN(SubCellInput2[50]) );
  AOI22_X1 LED_RoundFunction2_U303 ( .A1(rst), .A2(Plaintext2[50]), .B1(
        LED_RoundFunction2_Feedback_50_), .B2(LED_RoundFunction2_n562), .ZN(
        LED_RoundFunction2_n763) );
  INV_X1 LED_RoundFunction2_U302 ( .A(Ciphertext2[50]), .ZN(
        LED_RoundFunction2_n764) );
  AOI22_X1 LED_RoundFunction2_U301 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n762), .B1(LED_RoundFunction2_n761), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U300 ( .A1(rst), .A2(Plaintext2[51]), .B1(
        LED_RoundFunction2_Feedback_51_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n761) );
  INV_X1 LED_RoundFunction2_U299 ( .A(Ciphertext2[51]), .ZN(
        LED_RoundFunction2_n762) );
  AOI22_X1 LED_RoundFunction2_U298 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n760), .B1(LED_RoundFunction2_n759), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U297 ( .A1(rst), .A2(Plaintext2[52]), .B1(
        LED_RoundFunction2_Feedback_52_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n759) );
  INV_X1 LED_RoundFunction2_U296 ( .A(Ciphertext2[52]), .ZN(
        LED_RoundFunction2_n760) );
  AOI22_X1 LED_RoundFunction2_U295 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n758), .B1(LED_RoundFunction2_n757), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U294 ( .A1(rst), .A2(Plaintext2[53]), .B1(
        LED_RoundFunction2_Feedback_53_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n757) );
  INV_X1 LED_RoundFunction2_U293 ( .A(Ciphertext2[53]), .ZN(
        LED_RoundFunction2_n758) );
  AOI22_X1 LED_RoundFunction2_U292 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n756), .B1(LED_RoundFunction2_n755), .B2(
        LED_RoundFunction2_n560), .ZN(SubCellInput2[54]) );
  AOI22_X1 LED_RoundFunction2_U291 ( .A1(rst), .A2(Plaintext2[54]), .B1(
        LED_RoundFunction2_Feedback_54_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n755) );
  INV_X1 LED_RoundFunction2_U290 ( .A(Ciphertext2[54]), .ZN(
        LED_RoundFunction2_n756) );
  AOI22_X1 LED_RoundFunction2_U289 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n754), .B1(LED_RoundFunction2_n753), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U288 ( .A1(rst), .A2(Plaintext2[55]), .B1(
        LED_RoundFunction2_Feedback_55_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n753) );
  INV_X1 LED_RoundFunction2_U287 ( .A(Ciphertext2[55]), .ZN(
        LED_RoundFunction2_n754) );
  AOI22_X1 LED_RoundFunction2_U286 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n752), .B1(LED_RoundFunction2_n751), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[1]) );
  AOI22_X1 LED_RoundFunction2_U285 ( .A1(rst), .A2(Plaintext2[59]), .B1(
        LED_RoundFunction2_Feedback_59_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n751) );
  INV_X1 LED_RoundFunction2_U284 ( .A(Ciphertext2[59]), .ZN(
        LED_RoundFunction2_n752) );
  AOI22_X1 LED_RoundFunction2_U283 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n750), .B1(LED_RoundFunction2_n749), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[0]) );
  AOI22_X1 LED_RoundFunction2_U282 ( .A1(rst), .A2(Plaintext2[60]), .B1(
        LED_RoundFunction2_Feedback_60_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n749) );
  INV_X1 LED_RoundFunction2_U281 ( .A(Ciphertext2[60]), .ZN(
        LED_RoundFunction2_n750) );
  AOI22_X1 LED_RoundFunction2_U280 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n748), .B1(LED_RoundFunction2_n747), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[2]) );
  AOI22_X1 LED_RoundFunction2_U279 ( .A1(rst), .A2(Plaintext2[61]), .B1(
        LED_RoundFunction2_Feedback_61_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n747) );
  INV_X1 LED_RoundFunction2_U278 ( .A(Ciphertext2[61]), .ZN(
        LED_RoundFunction2_n748) );
  AOI22_X1 LED_RoundFunction2_U277 ( .A1(LED_RoundFunction2_n555), .A2(
        LED_RoundFunction2_n746), .B1(LED_RoundFunction2_n745), .B2(
        LED_RoundFunction2_n560), .ZN(SubCellInput2[62]) );
  AOI22_X1 LED_RoundFunction2_U276 ( .A1(rst), .A2(Plaintext2[62]), .B1(
        LED_RoundFunction2_Feedback_62_), .B2(LED_RoundFunction2_n563), .ZN(
        LED_RoundFunction2_n745) );
  INV_X1 LED_RoundFunction2_U275 ( .A(Ciphertext2[62]), .ZN(
        LED_RoundFunction2_n746) );
  XOR2_X1 LED_RoundFunction2_U274 ( .A(1'b0), .B(LED_RoundFunction2_n744), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[2]) );
  AOI21_X1 LED_RoundFunction2_U273 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n743), .A(LED_RoundFunction2_n742), .ZN(
        LED_RoundFunction2_n744) );
  AOI221_X1 LED_RoundFunction2_U272 ( .B1(Plaintext2[9]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_9_), .C2(LED_RoundFunction2_n568), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n742) );
  INV_X1 LED_RoundFunction2_U271 ( .A(Ciphertext2[9]), .ZN(
        LED_RoundFunction2_n743) );
  XOR2_X1 LED_RoundFunction2_U270 ( .A(1'b0), .B(LED_RoundFunction2_n741), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[0]) );
  AOI21_X1 LED_RoundFunction2_U269 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n740), .A(LED_RoundFunction2_n739), .ZN(
        LED_RoundFunction2_n741) );
  AOI221_X1 LED_RoundFunction2_U268 ( .B1(Plaintext2[8]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_8_), .C2(LED_RoundFunction2_n566), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n739) );
  INV_X1 LED_RoundFunction2_U267 ( .A(Ciphertext2[8]), .ZN(
        LED_RoundFunction2_n740) );
  AOI22_X1 LED_RoundFunction2_U266 ( .A1(LED_RoundFunction2_n555), .A2(
        Ciphertext2[63]), .B1(LED_RoundFunction2_n738), .B2(
        LED_RoundFunction2_n560), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[1]) );
  INV_X1 LED_RoundFunction2_U265 ( .A(LED_RoundFunction2_n737), .ZN(
        LED_RoundFunction2_n738) );
  OAI22_X1 LED_RoundFunction2_U264 ( .A1(LED_RoundFunction2_n565), .A2(
        Plaintext2[63]), .B1(LED_RoundFunction2_Feedback_63_), .B2(rst), .ZN(
        LED_RoundFunction2_n737) );
  XOR2_X1 LED_RoundFunction2_U263 ( .A(1'b0), .B(LED_RoundFunction2_n736), .Z(
        SubCellInput2[58]) );
  AOI21_X1 LED_RoundFunction2_U262 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n735), .A(LED_RoundFunction2_n734), .ZN(
        LED_RoundFunction2_n736) );
  AOI221_X1 LED_RoundFunction2_U261 ( .B1(Plaintext2[58]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_58_), .C2(LED_RoundFunction2_n565), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n734) );
  INV_X1 LED_RoundFunction2_U260 ( .A(Ciphertext2[58]), .ZN(
        LED_RoundFunction2_n735) );
  XOR2_X1 LED_RoundFunction2_U259 ( .A(1'b0), .B(LED_RoundFunction2_n733), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[2]) );
  AOI21_X1 LED_RoundFunction2_U258 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n732), .A(LED_RoundFunction2_n731), .ZN(
        LED_RoundFunction2_n733) );
  AOI221_X1 LED_RoundFunction2_U257 ( .B1(Plaintext2[57]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_57_), .C2(LED_RoundFunction2_n566), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n731) );
  INV_X1 LED_RoundFunction2_U256 ( .A(Ciphertext2[57]), .ZN(
        LED_RoundFunction2_n732) );
  XOR2_X1 LED_RoundFunction2_U255 ( .A(1'b0), .B(LED_RoundFunction2_n730), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[0]) );
  AOI21_X1 LED_RoundFunction2_U254 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n729), .A(LED_RoundFunction2_n728), .ZN(
        LED_RoundFunction2_n730) );
  AOI221_X1 LED_RoundFunction2_U253 ( .B1(Plaintext2[56]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_56_), .C2(LED_RoundFunction2_n568), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n728) );
  INV_X1 LED_RoundFunction2_U252 ( .A(Ciphertext2[56]), .ZN(
        LED_RoundFunction2_n729) );
  AOI22_X1 LED_RoundFunction2_U251 ( .A1(LED_RoundFunction2_n555), .A2(
        Ciphertext2[47]), .B1(LED_RoundFunction2_n727), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[1]) );
  INV_X1 LED_RoundFunction2_U250 ( .A(LED_RoundFunction2_n726), .ZN(
        LED_RoundFunction2_n727) );
  OAI22_X1 LED_RoundFunction2_U249 ( .A1(LED_RoundFunction2_n568), .A2(
        Plaintext2[47]), .B1(LED_RoundFunction2_Feedback_47_), .B2(rst), .ZN(
        LED_RoundFunction2_n726) );
  AOI22_X1 LED_RoundFunction2_U248 ( .A1(LED_RoundFunction2_n556), .A2(
        Ciphertext2[44]), .B1(LED_RoundFunction2_n725), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[0]) );
  INV_X1 LED_RoundFunction2_U247 ( .A(LED_RoundFunction2_n724), .ZN(
        LED_RoundFunction2_n725) );
  OAI22_X1 LED_RoundFunction2_U246 ( .A1(LED_RoundFunction2_n568), .A2(
        Plaintext2[44]), .B1(LED_RoundFunction2_Feedback_44_), .B2(rst), .ZN(
        LED_RoundFunction2_n724) );
  XOR2_X1 LED_RoundFunction2_U245 ( .A(1'b0), .B(LED_RoundFunction2_n723), .Z(
        SubCellInput2[42]) );
  AOI21_X1 LED_RoundFunction2_U244 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n722), .A(LED_RoundFunction2_n721), .ZN(
        LED_RoundFunction2_n723) );
  AOI221_X1 LED_RoundFunction2_U243 ( .B1(Plaintext2[42]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_42_), .C2(LED_RoundFunction2_n568), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n721) );
  INV_X1 LED_RoundFunction2_U242 ( .A(Ciphertext2[42]), .ZN(
        LED_RoundFunction2_n722) );
  XOR2_X1 LED_RoundFunction2_U241 ( .A(1'b0), .B(LED_RoundFunction2_n720), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[2]) );
  AOI21_X1 LED_RoundFunction2_U240 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n719), .A(LED_RoundFunction2_n718), .ZN(
        LED_RoundFunction2_n720) );
  AOI221_X1 LED_RoundFunction2_U239 ( .B1(Plaintext2[41]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_41_), .C2(LED_RoundFunction2_n565), .A(
        LED_RoundFunction2_n557), .ZN(LED_RoundFunction2_n718) );
  INV_X1 LED_RoundFunction2_U238 ( .A(Ciphertext2[41]), .ZN(
        LED_RoundFunction2_n719) );
  XOR2_X1 LED_RoundFunction2_U237 ( .A(1'b0), .B(LED_RoundFunction2_n717), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[0]) );
  AOI21_X1 LED_RoundFunction2_U236 ( .B1(LED_RoundFunction2_n557), .B2(
        LED_RoundFunction2_n716), .A(LED_RoundFunction2_n715), .ZN(
        LED_RoundFunction2_n717) );
  AOI221_X1 LED_RoundFunction2_U235 ( .B1(Plaintext2[40]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_40_), .C2(LED_RoundFunction2_n568), .A(
        LED_RoundFunction2_n557), .ZN(LED_RoundFunction2_n715) );
  INV_X1 LED_RoundFunction2_U234 ( .A(Ciphertext2[40]), .ZN(
        LED_RoundFunction2_n716) );
  AOI22_X1 LED_RoundFunction2_U233 ( .A1(LED_RoundFunction2_n556), .A2(
        Ciphertext2[29]), .B1(LED_RoundFunction2_n714), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[2]) );
  INV_X1 LED_RoundFunction2_U232 ( .A(LED_RoundFunction2_n713), .ZN(
        LED_RoundFunction2_n714) );
  OAI22_X1 LED_RoundFunction2_U231 ( .A1(LED_RoundFunction2_n565), .A2(
        Plaintext2[29]), .B1(LED_RoundFunction2_Feedback_29_), .B2(rst), .ZN(
        LED_RoundFunction2_n713) );
  XOR2_X1 LED_RoundFunction2_U230 ( .A(1'b0), .B(LED_RoundFunction2_n712), .Z(
        SubCellInput2[26]) );
  AOI21_X1 LED_RoundFunction2_U229 ( .B1(LED_RoundFunction2_n558), .B2(
        LED_RoundFunction2_n711), .A(LED_RoundFunction2_n710), .ZN(
        LED_RoundFunction2_n712) );
  AOI221_X1 LED_RoundFunction2_U228 ( .B1(Plaintext2[26]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_26_), .C2(LED_RoundFunction2_n568), .A(
        LED_RoundFunction2_n557), .ZN(LED_RoundFunction2_n710) );
  INV_X1 LED_RoundFunction2_U227 ( .A(Ciphertext2[26]), .ZN(
        LED_RoundFunction2_n711) );
  XOR2_X1 LED_RoundFunction2_U226 ( .A(1'b0), .B(LED_RoundFunction2_n709), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[2]) );
  AOI21_X1 LED_RoundFunction2_U225 ( .B1(LED_RoundFunction2_n558), .B2(
        LED_RoundFunction2_n708), .A(LED_RoundFunction2_n707), .ZN(
        LED_RoundFunction2_n709) );
  AOI221_X1 LED_RoundFunction2_U224 ( .B1(Plaintext2[25]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_25_), .C2(LED_RoundFunction2_n568), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n707) );
  INV_X1 LED_RoundFunction2_U223 ( .A(Ciphertext2[25]), .ZN(
        LED_RoundFunction2_n708) );
  XOR2_X1 LED_RoundFunction2_U222 ( .A(1'b0), .B(LED_RoundFunction2_n706), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[0]) );
  AOI21_X1 LED_RoundFunction2_U221 ( .B1(LED_RoundFunction2_n558), .B2(
        LED_RoundFunction2_n705), .A(LED_RoundFunction2_n704), .ZN(
        LED_RoundFunction2_n706) );
  AOI221_X1 LED_RoundFunction2_U220 ( .B1(Plaintext2[24]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_24_), .C2(LED_RoundFunction2_n566), .A(
        LED_RoundFunction2_n557), .ZN(LED_RoundFunction2_n704) );
  INV_X1 LED_RoundFunction2_U219 ( .A(Ciphertext2[24]), .ZN(
        LED_RoundFunction2_n705) );
  AOI22_X1 LED_RoundFunction2_U218 ( .A1(LED_RoundFunction2_n556), .A2(
        Ciphertext2[13]), .B1(LED_RoundFunction2_n703), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[2]) );
  INV_X1 LED_RoundFunction2_U217 ( .A(LED_RoundFunction2_n702), .ZN(
        LED_RoundFunction2_n703) );
  OAI22_X1 LED_RoundFunction2_U216 ( .A1(LED_RoundFunction2_n568), .A2(
        Plaintext2[13]), .B1(LED_RoundFunction2_Feedback_13_), .B2(rst), .ZN(
        LED_RoundFunction2_n702) );
  AOI22_X1 LED_RoundFunction2_U215 ( .A1(LED_RoundFunction2_n556), .A2(
        Ciphertext2[12]), .B1(LED_RoundFunction2_n701), .B2(
        LED_RoundFunction2_n559), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[0]) );
  INV_X1 LED_RoundFunction2_U214 ( .A(LED_RoundFunction2_n700), .ZN(
        LED_RoundFunction2_n701) );
  OAI22_X1 LED_RoundFunction2_U213 ( .A1(LED_RoundFunction2_n565), .A2(
        Plaintext2[12]), .B1(LED_RoundFunction2_Feedback_12_), .B2(rst), .ZN(
        LED_RoundFunction2_n700) );
  XOR2_X1 LED_RoundFunction2_U212 ( .A(1'b0), .B(LED_RoundFunction2_n699), .Z(
        SubCellInput2[10]) );
  AOI21_X1 LED_RoundFunction2_U211 ( .B1(LED_RoundFunction2_n558), .B2(
        LED_RoundFunction2_n698), .A(LED_RoundFunction2_n697), .ZN(
        LED_RoundFunction2_n699) );
  AOI221_X1 LED_RoundFunction2_U210 ( .B1(Plaintext2[10]), .B2(rst), .C1(
        LED_RoundFunction2_Feedback_10_), .C2(LED_RoundFunction2_n565), .A(
        LED_RoundFunction2_n556), .ZN(LED_RoundFunction2_n697) );
  INV_X1 LED_RoundFunction2_U209 ( .A(Ciphertext2[10]), .ZN(
        LED_RoundFunction2_n698) );
  AOI22_X1 LED_RoundFunction2_U208 ( .A1(rst), .A2(LED_RoundFunction2_n696), 
        .B1(LED_RoundFunction2_n695), .B2(LED_RoundFunction2_n563), .ZN(
        Ciphertext2[9]) );
  XNOR2_X1 LED_RoundFunction2_U207 ( .A(LED_RoundFunction2_Feedback_9_), .B(
        Key2[73]), .ZN(LED_RoundFunction2_n695) );
  XNOR2_X1 LED_RoundFunction2_U206 ( .A(Plaintext2[9]), .B(Key2[9]), .ZN(
        LED_RoundFunction2_n696) );
  AOI22_X1 LED_RoundFunction2_U205 ( .A1(rst), .A2(LED_RoundFunction2_n694), 
        .B1(LED_RoundFunction2_n693), .B2(LED_RoundFunction2_n563), .ZN(
        Ciphertext2[8]) );
  XNOR2_X1 LED_RoundFunction2_U204 ( .A(LED_RoundFunction2_Feedback_8_), .B(
        Key2[72]), .ZN(LED_RoundFunction2_n693) );
  XNOR2_X1 LED_RoundFunction2_U203 ( .A(Plaintext2[8]), .B(Key2[8]), .ZN(
        LED_RoundFunction2_n694) );
  AOI22_X1 LED_RoundFunction2_U202 ( .A1(rst), .A2(LED_RoundFunction2_n692), 
        .B1(LED_RoundFunction2_n691), .B2(LED_RoundFunction2_n563), .ZN(
        Ciphertext2[7]) );
  XNOR2_X1 LED_RoundFunction2_U201 ( .A(LED_RoundFunction2_Feedback_7_), .B(
        Key2[71]), .ZN(LED_RoundFunction2_n691) );
  XNOR2_X1 LED_RoundFunction2_U200 ( .A(Plaintext2[7]), .B(Key2[7]), .ZN(
        LED_RoundFunction2_n692) );
  AOI22_X1 LED_RoundFunction2_U199 ( .A1(rst), .A2(LED_RoundFunction2_n690), 
        .B1(LED_RoundFunction2_n689), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[6]) );
  XNOR2_X1 LED_RoundFunction2_U198 ( .A(LED_RoundFunction2_Feedback_6_), .B(
        Key2[70]), .ZN(LED_RoundFunction2_n689) );
  XNOR2_X1 LED_RoundFunction2_U197 ( .A(Plaintext2[6]), .B(Key2[6]), .ZN(
        LED_RoundFunction2_n690) );
  AOI22_X1 LED_RoundFunction2_U196 ( .A1(rst), .A2(LED_RoundFunction2_n688), 
        .B1(LED_RoundFunction2_n687), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[63]) );
  XNOR2_X1 LED_RoundFunction2_U195 ( .A(LED_RoundFunction2_Feedback_63_), .B(
        Key2[127]), .ZN(LED_RoundFunction2_n687) );
  XNOR2_X1 LED_RoundFunction2_U194 ( .A(Plaintext2[63]), .B(Key2[63]), .ZN(
        LED_RoundFunction2_n688) );
  AOI22_X1 LED_RoundFunction2_U193 ( .A1(rst), .A2(LED_RoundFunction2_n686), 
        .B1(LED_RoundFunction2_n685), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[5]) );
  XNOR2_X1 LED_RoundFunction2_U192 ( .A(LED_RoundFunction2_Feedback_5_), .B(
        Key2[69]), .ZN(LED_RoundFunction2_n685) );
  XNOR2_X1 LED_RoundFunction2_U191 ( .A(Plaintext2[5]), .B(Key2[5]), .ZN(
        LED_RoundFunction2_n686) );
  AOI22_X1 LED_RoundFunction2_U190 ( .A1(rst), .A2(LED_RoundFunction2_n684), 
        .B1(LED_RoundFunction2_n683), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[58]) );
  XNOR2_X1 LED_RoundFunction2_U189 ( .A(LED_RoundFunction2_Feedback_58_), .B(
        Key2[122]), .ZN(LED_RoundFunction2_n683) );
  XNOR2_X1 LED_RoundFunction2_U188 ( .A(Plaintext2[58]), .B(Key2[58]), .ZN(
        LED_RoundFunction2_n684) );
  AOI22_X1 LED_RoundFunction2_U187 ( .A1(rst), .A2(LED_RoundFunction2_n682), 
        .B1(LED_RoundFunction2_n681), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[57]) );
  XNOR2_X1 LED_RoundFunction2_U186 ( .A(LED_RoundFunction2_Feedback_57_), .B(
        Key2[121]), .ZN(LED_RoundFunction2_n681) );
  XNOR2_X1 LED_RoundFunction2_U185 ( .A(Plaintext2[57]), .B(Key2[57]), .ZN(
        LED_RoundFunction2_n682) );
  AOI22_X1 LED_RoundFunction2_U184 ( .A1(rst), .A2(LED_RoundFunction2_n680), 
        .B1(LED_RoundFunction2_n679), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[56]) );
  XNOR2_X1 LED_RoundFunction2_U183 ( .A(LED_RoundFunction2_Feedback_56_), .B(
        Key2[120]), .ZN(LED_RoundFunction2_n679) );
  XNOR2_X1 LED_RoundFunction2_U182 ( .A(Plaintext2[56]), .B(Key2[56]), .ZN(
        LED_RoundFunction2_n680) );
  AOI22_X1 LED_RoundFunction2_U181 ( .A1(rst), .A2(LED_RoundFunction2_n678), 
        .B1(LED_RoundFunction2_n677), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[55]) );
  XNOR2_X1 LED_RoundFunction2_U180 ( .A(LED_RoundFunction2_Feedback_55_), .B(
        Key2[119]), .ZN(LED_RoundFunction2_n677) );
  XNOR2_X1 LED_RoundFunction2_U179 ( .A(Plaintext2[55]), .B(Key2[55]), .ZN(
        LED_RoundFunction2_n678) );
  AOI22_X1 LED_RoundFunction2_U178 ( .A1(rst), .A2(LED_RoundFunction2_n676), 
        .B1(LED_RoundFunction2_n675), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[54]) );
  XNOR2_X1 LED_RoundFunction2_U177 ( .A(LED_RoundFunction2_Feedback_54_), .B(
        Key2[118]), .ZN(LED_RoundFunction2_n675) );
  XNOR2_X1 LED_RoundFunction2_U176 ( .A(Plaintext2[54]), .B(Key2[54]), .ZN(
        LED_RoundFunction2_n676) );
  AOI22_X1 LED_RoundFunction2_U175 ( .A1(rst), .A2(LED_RoundFunction2_n674), 
        .B1(LED_RoundFunction2_n673), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[53]) );
  XNOR2_X1 LED_RoundFunction2_U174 ( .A(LED_RoundFunction2_Feedback_53_), .B(
        Key2[117]), .ZN(LED_RoundFunction2_n673) );
  XNOR2_X1 LED_RoundFunction2_U173 ( .A(Plaintext2[53]), .B(Key2[53]), .ZN(
        LED_RoundFunction2_n674) );
  AOI22_X1 LED_RoundFunction2_U172 ( .A1(rst), .A2(LED_RoundFunction2_n672), 
        .B1(LED_RoundFunction2_n671), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[52]) );
  XNOR2_X1 LED_RoundFunction2_U171 ( .A(LED_RoundFunction2_Feedback_52_), .B(
        Key2[116]), .ZN(LED_RoundFunction2_n671) );
  XNOR2_X1 LED_RoundFunction2_U170 ( .A(Plaintext2[52]), .B(Key2[52]), .ZN(
        LED_RoundFunction2_n672) );
  AOI22_X1 LED_RoundFunction2_U169 ( .A1(rst), .A2(LED_RoundFunction2_n670), 
        .B1(LED_RoundFunction2_n669), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[51]) );
  XNOR2_X1 LED_RoundFunction2_U168 ( .A(LED_RoundFunction2_Feedback_51_), .B(
        Key2[115]), .ZN(LED_RoundFunction2_n669) );
  XNOR2_X1 LED_RoundFunction2_U167 ( .A(Plaintext2[51]), .B(Key2[51]), .ZN(
        LED_RoundFunction2_n670) );
  AOI22_X1 LED_RoundFunction2_U166 ( .A1(rst), .A2(LED_RoundFunction2_n668), 
        .B1(LED_RoundFunction2_n667), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[50]) );
  XNOR2_X1 LED_RoundFunction2_U165 ( .A(LED_RoundFunction2_Feedback_50_), .B(
        Key2[114]), .ZN(LED_RoundFunction2_n667) );
  XNOR2_X1 LED_RoundFunction2_U164 ( .A(Plaintext2[50]), .B(Key2[50]), .ZN(
        LED_RoundFunction2_n668) );
  AOI22_X1 LED_RoundFunction2_U163 ( .A1(rst), .A2(LED_RoundFunction2_n666), 
        .B1(LED_RoundFunction2_n665), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[4]) );
  XNOR2_X1 LED_RoundFunction2_U162 ( .A(LED_RoundFunction2_Feedback_4_), .B(
        Key2[68]), .ZN(LED_RoundFunction2_n665) );
  XNOR2_X1 LED_RoundFunction2_U161 ( .A(Plaintext2[4]), .B(Key2[4]), .ZN(
        LED_RoundFunction2_n666) );
  AOI22_X1 LED_RoundFunction2_U160 ( .A1(rst), .A2(LED_RoundFunction2_n664), 
        .B1(LED_RoundFunction2_n663), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[49]) );
  XNOR2_X1 LED_RoundFunction2_U159 ( .A(LED_RoundFunction2_Feedback_49_), .B(
        Key2[113]), .ZN(LED_RoundFunction2_n663) );
  XNOR2_X1 LED_RoundFunction2_U158 ( .A(Plaintext2[49]), .B(Key2[49]), .ZN(
        LED_RoundFunction2_n664) );
  AOI22_X1 LED_RoundFunction2_U157 ( .A1(rst), .A2(LED_RoundFunction2_n662), 
        .B1(LED_RoundFunction2_n661), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[48]) );
  XNOR2_X1 LED_RoundFunction2_U156 ( .A(LED_RoundFunction2_Feedback_48_), .B(
        Key2[112]), .ZN(LED_RoundFunction2_n661) );
  XNOR2_X1 LED_RoundFunction2_U155 ( .A(Plaintext2[48]), .B(Key2[48]), .ZN(
        LED_RoundFunction2_n662) );
  AOI22_X1 LED_RoundFunction2_U154 ( .A1(rst), .A2(LED_RoundFunction2_n660), 
        .B1(LED_RoundFunction2_n659), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[47]) );
  XNOR2_X1 LED_RoundFunction2_U153 ( .A(LED_RoundFunction2_Feedback_47_), .B(
        Key2[111]), .ZN(LED_RoundFunction2_n659) );
  XNOR2_X1 LED_RoundFunction2_U152 ( .A(Plaintext2[47]), .B(Key2[47]), .ZN(
        LED_RoundFunction2_n660) );
  AOI22_X1 LED_RoundFunction2_U151 ( .A1(rst), .A2(LED_RoundFunction2_n658), 
        .B1(LED_RoundFunction2_n657), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[44]) );
  XNOR2_X1 LED_RoundFunction2_U150 ( .A(LED_RoundFunction2_Feedback_44_), .B(
        Key2[108]), .ZN(LED_RoundFunction2_n657) );
  XNOR2_X1 LED_RoundFunction2_U149 ( .A(Plaintext2[44]), .B(Key2[44]), .ZN(
        LED_RoundFunction2_n658) );
  AOI22_X1 LED_RoundFunction2_U148 ( .A1(rst), .A2(LED_RoundFunction2_n656), 
        .B1(LED_RoundFunction2_n655), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[42]) );
  XNOR2_X1 LED_RoundFunction2_U147 ( .A(LED_RoundFunction2_Feedback_42_), .B(
        Key2[106]), .ZN(LED_RoundFunction2_n655) );
  XNOR2_X1 LED_RoundFunction2_U146 ( .A(Plaintext2[42]), .B(Key2[42]), .ZN(
        LED_RoundFunction2_n656) );
  AOI22_X1 LED_RoundFunction2_U145 ( .A1(rst), .A2(LED_RoundFunction2_n654), 
        .B1(LED_RoundFunction2_n653), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[41]) );
  XNOR2_X1 LED_RoundFunction2_U144 ( .A(LED_RoundFunction2_Feedback_41_), .B(
        Key2[105]), .ZN(LED_RoundFunction2_n653) );
  XNOR2_X1 LED_RoundFunction2_U143 ( .A(Plaintext2[41]), .B(Key2[41]), .ZN(
        LED_RoundFunction2_n654) );
  AOI22_X1 LED_RoundFunction2_U142 ( .A1(rst), .A2(LED_RoundFunction2_n652), 
        .B1(LED_RoundFunction2_n651), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[40]) );
  XNOR2_X1 LED_RoundFunction2_U141 ( .A(LED_RoundFunction2_Feedback_40_), .B(
        Key2[104]), .ZN(LED_RoundFunction2_n651) );
  XNOR2_X1 LED_RoundFunction2_U140 ( .A(Plaintext2[40]), .B(Key2[40]), .ZN(
        LED_RoundFunction2_n652) );
  AOI22_X1 LED_RoundFunction2_U139 ( .A1(rst), .A2(LED_RoundFunction2_n650), 
        .B1(LED_RoundFunction2_n649), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[3]) );
  XNOR2_X1 LED_RoundFunction2_U138 ( .A(LED_RoundFunction2_Feedback_3_), .B(
        Key2[67]), .ZN(LED_RoundFunction2_n649) );
  XNOR2_X1 LED_RoundFunction2_U137 ( .A(Plaintext2[3]), .B(Key2[3]), .ZN(
        LED_RoundFunction2_n650) );
  AOI22_X1 LED_RoundFunction2_U136 ( .A1(rst), .A2(LED_RoundFunction2_n648), 
        .B1(LED_RoundFunction2_n647), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[39]) );
  XNOR2_X1 LED_RoundFunction2_U135 ( .A(LED_RoundFunction2_Feedback_39_), .B(
        Key2[103]), .ZN(LED_RoundFunction2_n647) );
  XNOR2_X1 LED_RoundFunction2_U134 ( .A(Plaintext2[39]), .B(Key2[39]), .ZN(
        LED_RoundFunction2_n648) );
  AOI22_X1 LED_RoundFunction2_U133 ( .A1(rst), .A2(LED_RoundFunction2_n646), 
        .B1(LED_RoundFunction2_n645), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[38]) );
  XNOR2_X1 LED_RoundFunction2_U132 ( .A(LED_RoundFunction2_Feedback_38_), .B(
        Key2[102]), .ZN(LED_RoundFunction2_n645) );
  XNOR2_X1 LED_RoundFunction2_U131 ( .A(Plaintext2[38]), .B(Key2[38]), .ZN(
        LED_RoundFunction2_n646) );
  AOI22_X1 LED_RoundFunction2_U130 ( .A1(rst), .A2(LED_RoundFunction2_n644), 
        .B1(LED_RoundFunction2_n643), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[37]) );
  XNOR2_X1 LED_RoundFunction2_U129 ( .A(LED_RoundFunction2_Feedback_37_), .B(
        Key2[101]), .ZN(LED_RoundFunction2_n643) );
  XNOR2_X1 LED_RoundFunction2_U128 ( .A(Plaintext2[37]), .B(Key2[37]), .ZN(
        LED_RoundFunction2_n644) );
  AOI22_X1 LED_RoundFunction2_U127 ( .A1(rst), .A2(LED_RoundFunction2_n642), 
        .B1(LED_RoundFunction2_n641), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[36]) );
  XNOR2_X1 LED_RoundFunction2_U126 ( .A(LED_RoundFunction2_Feedback_36_), .B(
        Key2[100]), .ZN(LED_RoundFunction2_n641) );
  XNOR2_X1 LED_RoundFunction2_U125 ( .A(Plaintext2[36]), .B(Key2[36]), .ZN(
        LED_RoundFunction2_n642) );
  AOI22_X1 LED_RoundFunction2_U124 ( .A1(rst), .A2(LED_RoundFunction2_n640), 
        .B1(LED_RoundFunction2_n639), .B2(LED_RoundFunction2_n568), .ZN(
        Ciphertext2[35]) );
  XNOR2_X1 LED_RoundFunction2_U123 ( .A(LED_RoundFunction2_Feedback_35_), .B(
        Key2[99]), .ZN(LED_RoundFunction2_n639) );
  XNOR2_X1 LED_RoundFunction2_U122 ( .A(Plaintext2[35]), .B(Key2[35]), .ZN(
        LED_RoundFunction2_n640) );
  AOI22_X1 LED_RoundFunction2_U121 ( .A1(rst), .A2(LED_RoundFunction2_n638), 
        .B1(LED_RoundFunction2_n637), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[34]) );
  XNOR2_X1 LED_RoundFunction2_U120 ( .A(LED_RoundFunction2_Feedback_34_), .B(
        Key2[98]), .ZN(LED_RoundFunction2_n637) );
  XNOR2_X1 LED_RoundFunction2_U119 ( .A(Plaintext2[34]), .B(Key2[34]), .ZN(
        LED_RoundFunction2_n638) );
  AOI22_X1 LED_RoundFunction2_U118 ( .A1(rst), .A2(LED_RoundFunction2_n636), 
        .B1(LED_RoundFunction2_n635), .B2(LED_RoundFunction2_n568), .ZN(
        Ciphertext2[33]) );
  XNOR2_X1 LED_RoundFunction2_U117 ( .A(LED_RoundFunction2_Feedback_33_), .B(
        Key2[97]), .ZN(LED_RoundFunction2_n635) );
  XNOR2_X1 LED_RoundFunction2_U116 ( .A(Plaintext2[33]), .B(Key2[33]), .ZN(
        LED_RoundFunction2_n636) );
  AOI22_X1 LED_RoundFunction2_U115 ( .A1(rst), .A2(LED_RoundFunction2_n634), 
        .B1(LED_RoundFunction2_n633), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[32]) );
  XNOR2_X1 LED_RoundFunction2_U114 ( .A(LED_RoundFunction2_Feedback_32_), .B(
        Key2[96]), .ZN(LED_RoundFunction2_n633) );
  XNOR2_X1 LED_RoundFunction2_U113 ( .A(Plaintext2[32]), .B(Key2[32]), .ZN(
        LED_RoundFunction2_n634) );
  AOI22_X1 LED_RoundFunction2_U112 ( .A1(rst), .A2(LED_RoundFunction2_n632), 
        .B1(LED_RoundFunction2_n631), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[2]) );
  XNOR2_X1 LED_RoundFunction2_U111 ( .A(LED_RoundFunction2_Feedback_2_), .B(
        Key2[66]), .ZN(LED_RoundFunction2_n631) );
  XNOR2_X1 LED_RoundFunction2_U110 ( .A(Plaintext2[2]), .B(Key2[2]), .ZN(
        LED_RoundFunction2_n632) );
  AOI22_X1 LED_RoundFunction2_U109 ( .A1(rst), .A2(LED_RoundFunction2_n630), 
        .B1(LED_RoundFunction2_n629), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[29]) );
  XNOR2_X1 LED_RoundFunction2_U108 ( .A(LED_RoundFunction2_Feedback_29_), .B(
        Key2[93]), .ZN(LED_RoundFunction2_n629) );
  XNOR2_X1 LED_RoundFunction2_U107 ( .A(Plaintext2[29]), .B(Key2[29]), .ZN(
        LED_RoundFunction2_n630) );
  AOI22_X1 LED_RoundFunction2_U106 ( .A1(rst), .A2(LED_RoundFunction2_n628), 
        .B1(LED_RoundFunction2_n627), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[26]) );
  XNOR2_X1 LED_RoundFunction2_U105 ( .A(LED_RoundFunction2_Feedback_26_), .B(
        Key2[90]), .ZN(LED_RoundFunction2_n627) );
  XNOR2_X1 LED_RoundFunction2_U104 ( .A(Plaintext2[26]), .B(Key2[26]), .ZN(
        LED_RoundFunction2_n628) );
  AOI22_X1 LED_RoundFunction2_U103 ( .A1(rst), .A2(LED_RoundFunction2_n626), 
        .B1(LED_RoundFunction2_n625), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[25]) );
  XNOR2_X1 LED_RoundFunction2_U102 ( .A(LED_RoundFunction2_Feedback_25_), .B(
        Key2[89]), .ZN(LED_RoundFunction2_n625) );
  XNOR2_X1 LED_RoundFunction2_U101 ( .A(Plaintext2[25]), .B(Key2[25]), .ZN(
        LED_RoundFunction2_n626) );
  AOI22_X1 LED_RoundFunction2_U100 ( .A1(rst), .A2(LED_RoundFunction2_n624), 
        .B1(LED_RoundFunction2_n623), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[24]) );
  XNOR2_X1 LED_RoundFunction2_U99 ( .A(LED_RoundFunction2_Feedback_24_), .B(
        Key2[88]), .ZN(LED_RoundFunction2_n623) );
  XNOR2_X1 LED_RoundFunction2_U98 ( .A(Plaintext2[24]), .B(Key2[24]), .ZN(
        LED_RoundFunction2_n624) );
  AOI22_X1 LED_RoundFunction2_U97 ( .A1(rst), .A2(LED_RoundFunction2_n622), 
        .B1(LED_RoundFunction2_n621), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[23]) );
  XNOR2_X1 LED_RoundFunction2_U96 ( .A(LED_RoundFunction2_Feedback_23_), .B(
        Key2[87]), .ZN(LED_RoundFunction2_n621) );
  XNOR2_X1 LED_RoundFunction2_U95 ( .A(Plaintext2[23]), .B(Key2[23]), .ZN(
        LED_RoundFunction2_n622) );
  AOI22_X1 LED_RoundFunction2_U94 ( .A1(rst), .A2(LED_RoundFunction2_n620), 
        .B1(LED_RoundFunction2_n619), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[22]) );
  XNOR2_X1 LED_RoundFunction2_U93 ( .A(LED_RoundFunction2_Feedback_22_), .B(
        Key2[86]), .ZN(LED_RoundFunction2_n619) );
  XNOR2_X1 LED_RoundFunction2_U92 ( .A(Plaintext2[22]), .B(Key2[22]), .ZN(
        LED_RoundFunction2_n620) );
  AOI22_X1 LED_RoundFunction2_U91 ( .A1(rst), .A2(LED_RoundFunction2_n618), 
        .B1(LED_RoundFunction2_n617), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[21]) );
  XNOR2_X1 LED_RoundFunction2_U90 ( .A(LED_RoundFunction2_Feedback_21_), .B(
        Key2[85]), .ZN(LED_RoundFunction2_n617) );
  XNOR2_X1 LED_RoundFunction2_U89 ( .A(Plaintext2[21]), .B(Key2[21]), .ZN(
        LED_RoundFunction2_n618) );
  AOI22_X1 LED_RoundFunction2_U88 ( .A1(rst), .A2(LED_RoundFunction2_n616), 
        .B1(LED_RoundFunction2_n615), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[20]) );
  XNOR2_X1 LED_RoundFunction2_U87 ( .A(LED_RoundFunction2_Feedback_20_), .B(
        Key2[84]), .ZN(LED_RoundFunction2_n615) );
  XNOR2_X1 LED_RoundFunction2_U86 ( .A(Plaintext2[20]), .B(Key2[20]), .ZN(
        LED_RoundFunction2_n616) );
  AOI22_X1 LED_RoundFunction2_U85 ( .A1(rst), .A2(LED_RoundFunction2_n614), 
        .B1(LED_RoundFunction2_n613), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[1]) );
  XNOR2_X1 LED_RoundFunction2_U84 ( .A(LED_RoundFunction2_Feedback_1_), .B(
        Key2[65]), .ZN(LED_RoundFunction2_n613) );
  XNOR2_X1 LED_RoundFunction2_U83 ( .A(Plaintext2[1]), .B(Key2[1]), .ZN(
        LED_RoundFunction2_n614) );
  AOI22_X1 LED_RoundFunction2_U82 ( .A1(rst), .A2(LED_RoundFunction2_n612), 
        .B1(LED_RoundFunction2_n611), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[19]) );
  XNOR2_X1 LED_RoundFunction2_U81 ( .A(LED_RoundFunction2_Feedback_19_), .B(
        Key2[83]), .ZN(LED_RoundFunction2_n611) );
  XNOR2_X1 LED_RoundFunction2_U80 ( .A(Plaintext2[19]), .B(Key2[19]), .ZN(
        LED_RoundFunction2_n612) );
  AOI22_X1 LED_RoundFunction2_U79 ( .A1(rst), .A2(LED_RoundFunction2_n610), 
        .B1(LED_RoundFunction2_n609), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[18]) );
  XNOR2_X1 LED_RoundFunction2_U78 ( .A(LED_RoundFunction2_Feedback_18_), .B(
        Key2[82]), .ZN(LED_RoundFunction2_n609) );
  XNOR2_X1 LED_RoundFunction2_U77 ( .A(Plaintext2[18]), .B(Key2[18]), .ZN(
        LED_RoundFunction2_n610) );
  AOI22_X1 LED_RoundFunction2_U76 ( .A1(rst), .A2(LED_RoundFunction2_n608), 
        .B1(LED_RoundFunction2_n607), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[17]) );
  XNOR2_X1 LED_RoundFunction2_U75 ( .A(LED_RoundFunction2_Feedback_17_), .B(
        Key2[81]), .ZN(LED_RoundFunction2_n607) );
  XNOR2_X1 LED_RoundFunction2_U74 ( .A(Plaintext2[17]), .B(Key2[17]), .ZN(
        LED_RoundFunction2_n608) );
  AOI22_X1 LED_RoundFunction2_U73 ( .A1(rst), .A2(LED_RoundFunction2_n606), 
        .B1(LED_RoundFunction2_n605), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[16]) );
  XNOR2_X1 LED_RoundFunction2_U72 ( .A(LED_RoundFunction2_Feedback_16_), .B(
        Key2[80]), .ZN(LED_RoundFunction2_n605) );
  XNOR2_X1 LED_RoundFunction2_U71 ( .A(Plaintext2[16]), .B(Key2[16]), .ZN(
        LED_RoundFunction2_n606) );
  AOI22_X1 LED_RoundFunction2_U70 ( .A1(rst), .A2(LED_RoundFunction2_n604), 
        .B1(LED_RoundFunction2_n603), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[13]) );
  XNOR2_X1 LED_RoundFunction2_U69 ( .A(LED_RoundFunction2_Feedback_13_), .B(
        Key2[77]), .ZN(LED_RoundFunction2_n603) );
  XNOR2_X1 LED_RoundFunction2_U68 ( .A(Plaintext2[13]), .B(Key2[13]), .ZN(
        LED_RoundFunction2_n604) );
  AOI22_X1 LED_RoundFunction2_U67 ( .A1(rst), .A2(LED_RoundFunction2_n602), 
        .B1(LED_RoundFunction2_n601), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[12]) );
  XNOR2_X1 LED_RoundFunction2_U66 ( .A(LED_RoundFunction2_Feedback_12_), .B(
        Key2[76]), .ZN(LED_RoundFunction2_n601) );
  XNOR2_X1 LED_RoundFunction2_U65 ( .A(Plaintext2[12]), .B(Key2[12]), .ZN(
        LED_RoundFunction2_n602) );
  AOI22_X1 LED_RoundFunction2_U64 ( .A1(rst), .A2(LED_RoundFunction2_n600), 
        .B1(LED_RoundFunction2_n599), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[10]) );
  XNOR2_X1 LED_RoundFunction2_U63 ( .A(LED_RoundFunction2_Feedback_10_), .B(
        Key2[74]), .ZN(LED_RoundFunction2_n599) );
  XNOR2_X1 LED_RoundFunction2_U62 ( .A(Plaintext2[10]), .B(Key2[10]), .ZN(
        LED_RoundFunction2_n600) );
  AOI22_X1 LED_RoundFunction2_U61 ( .A1(rst), .A2(LED_RoundFunction2_n598), 
        .B1(LED_RoundFunction2_n597), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[0]) );
  XNOR2_X1 LED_RoundFunction2_U60 ( .A(LED_RoundFunction2_Feedback_0_), .B(
        Key2[64]), .ZN(LED_RoundFunction2_n597) );
  XNOR2_X1 LED_RoundFunction2_U59 ( .A(Plaintext2[0]), .B(Key2[0]), .ZN(
        LED_RoundFunction2_n598) );
  AOI22_X1 LED_RoundFunction2_U58 ( .A1(rst), .A2(LED_RoundFunction2_n596), 
        .B1(LED_RoundFunction2_n595), .B2(LED_RoundFunction2_n568), .ZN(
        Ciphertext2[46]) );
  XNOR2_X1 LED_RoundFunction2_U57 ( .A(LED_RoundFunction2_Feedback_46_), .B(
        Key2[110]), .ZN(LED_RoundFunction2_n595) );
  XNOR2_X1 LED_RoundFunction2_U56 ( .A(Plaintext2[46]), .B(Key2[46]), .ZN(
        LED_RoundFunction2_n596) );
  AOI22_X1 LED_RoundFunction2_U55 ( .A1(rst), .A2(LED_RoundFunction2_n594), 
        .B1(LED_RoundFunction2_n593), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[45]) );
  XNOR2_X1 LED_RoundFunction2_U54 ( .A(LED_RoundFunction2_Feedback_45_), .B(
        Key2[109]), .ZN(LED_RoundFunction2_n593) );
  XNOR2_X1 LED_RoundFunction2_U53 ( .A(Plaintext2[45]), .B(Key2[45]), .ZN(
        LED_RoundFunction2_n594) );
  AOI22_X1 LED_RoundFunction2_U52 ( .A1(rst), .A2(LED_RoundFunction2_n592), 
        .B1(LED_RoundFunction2_n591), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[43]) );
  XNOR2_X1 LED_RoundFunction2_U51 ( .A(LED_RoundFunction2_Feedback_43_), .B(
        Key2[107]), .ZN(LED_RoundFunction2_n591) );
  XNOR2_X1 LED_RoundFunction2_U50 ( .A(Plaintext2[43]), .B(Key2[43]), .ZN(
        LED_RoundFunction2_n592) );
  AOI22_X1 LED_RoundFunction2_U49 ( .A1(rst), .A2(LED_RoundFunction2_n590), 
        .B1(LED_RoundFunction2_n589), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[31]) );
  XNOR2_X1 LED_RoundFunction2_U48 ( .A(LED_RoundFunction2_Feedback_31_), .B(
        Key2[95]), .ZN(LED_RoundFunction2_n589) );
  XNOR2_X1 LED_RoundFunction2_U47 ( .A(Plaintext2[31]), .B(Key2[31]), .ZN(
        LED_RoundFunction2_n590) );
  AOI22_X1 LED_RoundFunction2_U46 ( .A1(rst), .A2(LED_RoundFunction2_n588), 
        .B1(LED_RoundFunction2_n587), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[30]) );
  XNOR2_X1 LED_RoundFunction2_U45 ( .A(LED_RoundFunction2_Feedback_30_), .B(
        Key2[94]), .ZN(LED_RoundFunction2_n587) );
  XNOR2_X1 LED_RoundFunction2_U44 ( .A(Plaintext2[30]), .B(Key2[30]), .ZN(
        LED_RoundFunction2_n588) );
  AOI22_X1 LED_RoundFunction2_U43 ( .A1(rst), .A2(LED_RoundFunction2_n586), 
        .B1(LED_RoundFunction2_n585), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[28]) );
  XNOR2_X1 LED_RoundFunction2_U42 ( .A(LED_RoundFunction2_Feedback_28_), .B(
        Key2[92]), .ZN(LED_RoundFunction2_n585) );
  XNOR2_X1 LED_RoundFunction2_U41 ( .A(Plaintext2[28]), .B(Key2[28]), .ZN(
        LED_RoundFunction2_n586) );
  AOI22_X1 LED_RoundFunction2_U40 ( .A1(rst), .A2(LED_RoundFunction2_n584), 
        .B1(LED_RoundFunction2_n583), .B2(LED_RoundFunction2_n564), .ZN(
        Ciphertext2[27]) );
  XNOR2_X1 LED_RoundFunction2_U39 ( .A(LED_RoundFunction2_Feedback_27_), .B(
        Key2[91]), .ZN(LED_RoundFunction2_n583) );
  XNOR2_X1 LED_RoundFunction2_U38 ( .A(Plaintext2[27]), .B(Key2[27]), .ZN(
        LED_RoundFunction2_n584) );
  AOI22_X1 LED_RoundFunction2_U37 ( .A1(rst), .A2(LED_RoundFunction2_n582), 
        .B1(LED_RoundFunction2_n581), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[15]) );
  XNOR2_X1 LED_RoundFunction2_U36 ( .A(LED_RoundFunction2_Feedback_15_), .B(
        Key2[79]), .ZN(LED_RoundFunction2_n581) );
  XNOR2_X1 LED_RoundFunction2_U35 ( .A(Plaintext2[15]), .B(Key2[15]), .ZN(
        LED_RoundFunction2_n582) );
  AOI22_X1 LED_RoundFunction2_U34 ( .A1(rst), .A2(LED_RoundFunction2_n580), 
        .B1(LED_RoundFunction2_n579), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[14]) );
  XNOR2_X1 LED_RoundFunction2_U33 ( .A(LED_RoundFunction2_Feedback_14_), .B(
        Key2[78]), .ZN(LED_RoundFunction2_n579) );
  XNOR2_X1 LED_RoundFunction2_U32 ( .A(Plaintext2[14]), .B(Key2[14]), .ZN(
        LED_RoundFunction2_n580) );
  AOI22_X1 LED_RoundFunction2_U31 ( .A1(rst), .A2(LED_RoundFunction2_n578), 
        .B1(LED_RoundFunction2_n577), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[11]) );
  XNOR2_X1 LED_RoundFunction2_U30 ( .A(LED_RoundFunction2_Feedback_11_), .B(
        Key2[75]), .ZN(LED_RoundFunction2_n577) );
  XNOR2_X1 LED_RoundFunction2_U29 ( .A(Plaintext2[11]), .B(Key2[11]), .ZN(
        LED_RoundFunction2_n578) );
  AOI22_X1 LED_RoundFunction2_U28 ( .A1(rst), .A2(LED_RoundFunction2_n576), 
        .B1(LED_RoundFunction2_n575), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[62]) );
  XNOR2_X1 LED_RoundFunction2_U27 ( .A(LED_RoundFunction2_Feedback_62_), .B(
        Key2[126]), .ZN(LED_RoundFunction2_n575) );
  XNOR2_X1 LED_RoundFunction2_U26 ( .A(Plaintext2[62]), .B(Key2[62]), .ZN(
        LED_RoundFunction2_n576) );
  AOI22_X1 LED_RoundFunction2_U25 ( .A1(rst), .A2(LED_RoundFunction2_n574), 
        .B1(LED_RoundFunction2_n573), .B2(LED_RoundFunction2_n565), .ZN(
        Ciphertext2[61]) );
  XNOR2_X1 LED_RoundFunction2_U24 ( .A(LED_RoundFunction2_Feedback_61_), .B(
        Key2[125]), .ZN(LED_RoundFunction2_n573) );
  XNOR2_X1 LED_RoundFunction2_U23 ( .A(Plaintext2[61]), .B(Key2[61]), .ZN(
        LED_RoundFunction2_n574) );
  AOI22_X1 LED_RoundFunction2_U22 ( .A1(rst), .A2(LED_RoundFunction2_n572), 
        .B1(LED_RoundFunction2_n571), .B2(LED_RoundFunction2_n566), .ZN(
        Ciphertext2[60]) );
  XNOR2_X1 LED_RoundFunction2_U21 ( .A(LED_RoundFunction2_Feedback_60_), .B(
        Key2[124]), .ZN(LED_RoundFunction2_n571) );
  XNOR2_X1 LED_RoundFunction2_U20 ( .A(Plaintext2[60]), .B(Key2[60]), .ZN(
        LED_RoundFunction2_n572) );
  AOI22_X1 LED_RoundFunction2_U19 ( .A1(rst), .A2(LED_RoundFunction2_n570), 
        .B1(LED_RoundFunction2_n569), .B2(LED_RoundFunction2_n567), .ZN(
        Ciphertext2[59]) );
  XNOR2_X1 LED_RoundFunction2_U18 ( .A(LED_RoundFunction2_Feedback_59_), .B(
        Key2[123]), .ZN(LED_RoundFunction2_n569) );
  XNOR2_X1 LED_RoundFunction2_U17 ( .A(Plaintext2[59]), .B(Key2[59]), .ZN(
        LED_RoundFunction2_n570) );
  BUF_X1 LED_RoundFunction2_U16 ( .A(LED_RoundFunction2_n568), .Z(
        LED_RoundFunction2_n562) );
  INV_X1 LED_RoundFunction2_U15 ( .A(AddKey), .ZN(LED_RoundFunction2_n561) );
  BUF_X1 LED_RoundFunction2_U14 ( .A(LED_RoundFunction2_n561), .Z(
        LED_RoundFunction2_n559) );
  INV_X1 LED_RoundFunction2_U13 ( .A(LED_RoundFunction2_n559), .ZN(
        LED_RoundFunction2_n557) );
  INV_X1 LED_RoundFunction2_U12 ( .A(rst), .ZN(LED_RoundFunction2_n568) );
  BUF_X1 LED_RoundFunction2_U11 ( .A(LED_RoundFunction2_n568), .Z(
        LED_RoundFunction2_n564) );
  BUF_X1 LED_RoundFunction2_U10 ( .A(LED_RoundFunction2_n568), .Z(
        LED_RoundFunction2_n566) );
  INV_X1 LED_RoundFunction2_U9 ( .A(LED_RoundFunction2_n559), .ZN(
        LED_RoundFunction2_n556) );
  BUF_X1 LED_RoundFunction2_U8 ( .A(LED_RoundFunction2_n568), .Z(
        LED_RoundFunction2_n565) );
  BUF_X1 LED_RoundFunction2_U7 ( .A(LED_RoundFunction2_n568), .Z(
        LED_RoundFunction2_n563) );
  INV_X1 LED_RoundFunction2_U6 ( .A(LED_RoundFunction2_n559), .ZN(
        LED_RoundFunction2_n558) );
  BUF_X1 LED_RoundFunction2_U5 ( .A(LED_RoundFunction2_n561), .Z(
        LED_RoundFunction2_n560) );
  BUF_X1 LED_RoundFunction2_U4 ( .A(LED_RoundFunction2_n568), .Z(
        LED_RoundFunction2_n567) );
  INV_X1 LED_RoundFunction2_U3 ( .A(LED_RoundFunction2_n559), .ZN(
        LED_RoundFunction2_n555) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U68 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n160), .B(
        LED_RoundFunction2_MCInst1_MC0_n159), .ZN(
        LED_RoundFunction2_Feedback_15_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U67 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n158), .B(SubCellOutput2[62]), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n160) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U66 ( .A(SubCellOutput2[3]), .B(
        LED_RoundFunction2_MCInst1_MC0_n157), .Z(
        LED_RoundFunction2_Feedback_14_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U65 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n156), .B(
        LED_RoundFunction2_MCInst1_MC0_n155), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n157) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U64 ( .A(SubCellOutput2[21]), .B(
        SubCellOutput2[1]), .ZN(LED_RoundFunction2_MCInst1_MC0_n155) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U63 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n154), .B(SubCellOutput2[41]), .Z(
        LED_RoundFunction2_MCInst1_MC0_n156) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U62 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n153), .B(
        LED_RoundFunction2_MCInst1_MC0_n152), .ZN(
        LED_RoundFunction2_Feedback_13_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U61 ( .A(SubCellOutput2[2]), .B(
        SubCellOutput2[40]), .ZN(LED_RoundFunction2_MCInst1_MC0_n152) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U60 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n151), .B(
        LED_RoundFunction2_MCInst1_MC0_n150), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n153) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U59 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n149), .B(
        LED_RoundFunction2_MCInst1_MC0_n148), .ZN(
        LED_RoundFunction2_Feedback_12_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U58 ( .A(SubCellOutput2[23]), .B(
        LED_RoundFunction2_MCInst1_MC0_n147), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n148) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U57 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n146), .B(
        LED_RoundFunction2_MCInst1_MC0_n150), .Z(
        LED_RoundFunction2_MCInst1_MC0_n149) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U56 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n145), .B(
        LED_RoundFunction2_MCInst1_MC0_n159), .Z(
        LED_RoundFunction2_MCInst1_MC0_n150) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC0_U55 ( .A1(SubCellOutput2[21]), .A2(
        SubCellOutput2[22]), .B1(LED_RoundFunction2_MCInst1_MC0_n144), .B2(
        LED_RoundFunction2_MCInst1_MC0_n143), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n146) );
  INV_X1 LED_RoundFunction2_MCInst1_MC0_U54 ( .A(SubCellOutput2[21]), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n143) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U53 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n142), .B(
        LED_RoundFunction2_MCInst1_MC0_n141), .ZN(
        LED_RoundFunction2_Feedback_31_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U52 ( .A(SubCellOutput2[43]), .B(
        LED_RoundFunction2_MCInst1_MC0_n140), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n141) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U51 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n139), .B(SubCellOutput2[60]), .Z(
        LED_RoundFunction2_MCInst1_MC0_n142) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC0_U50 ( .A1(SubCellOutput2[42]), .A2(
        SubCellOutput2[22]), .B1(LED_RoundFunction2_MCInst1_MC0_n144), .B2(
        LED_RoundFunction2_MCInst1_MC0_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n139) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U49 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n137), .B(
        LED_RoundFunction2_MCInst1_MC0_n136), .ZN(
        LED_RoundFunction2_Feedback_30_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U48 ( .A(SubCellOutput2[40]), .B(
        LED_RoundFunction2_MCInst1_MC0_n135), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n136) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U47 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n134), .B(
        LED_RoundFunction2_MCInst1_MC0_n133), .Z(
        LED_RoundFunction2_MCInst1_MC0_n137) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC0_U46 ( .A1(SubCellOutput2[22]), .A2(
        SubCellOutput2[61]), .B1(LED_RoundFunction2_MCInst1_MC0_n132), .B2(
        LED_RoundFunction2_MCInst1_MC0_n144), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n134) );
  INV_X1 LED_RoundFunction2_MCInst1_MC0_U45 ( .A(SubCellOutput2[22]), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n144) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U44 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n131), .B(
        LED_RoundFunction2_MCInst1_MC0_n151), .ZN(
        LED_RoundFunction2_Feedback_29_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U43 ( .A(SubCellOutput2[63]), .B(
        SubCellOutput2[60]), .ZN(LED_RoundFunction2_MCInst1_MC0_n151) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U42 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n130), .B(
        LED_RoundFunction2_MCInst1_MC0_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n131) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U41 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n128), .B(
        LED_RoundFunction2_MCInst1_MC0_n127), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n130) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U40 ( .A(SubCellOutput2[21]), .B(
        LED_RoundFunction2_MCInst1_MC0_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n127) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U39 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n125), .B(SubCellOutput2[20]), .Z(
        LED_RoundFunction2_MCInst1_MC0_n128) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U38 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n124), .B(
        LED_RoundFunction2_MCInst1_MC0_n123), .ZN(
        LED_RoundFunction2_Feedback_28_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U37 ( .A(SubCellOutput2[0]), .B(
        LED_RoundFunction2_MCInst1_MC0_n122), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n124) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U36 ( .A(SubCellOutput2[2]), .B(
        LED_RoundFunction2_MCInst1_MC0_n122), .ZN(
        LED_RoundFunction2_Feedback_47_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U35 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n135), .B(
        LED_RoundFunction2_MCInst1_MC0_n121), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n122) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U34 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n120), .B(
        LED_RoundFunction2_MCInst1_MC0_n125), .Z(
        LED_RoundFunction2_MCInst1_MC0_n135) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U33 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n119), .B(
        LED_RoundFunction2_MCInst1_MC0_n118), .ZN(
        LED_RoundFunction2_Feedback_46_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U32 ( .A(SubCellOutput2[22]), .B(
        LED_RoundFunction2_MCInst1_MC0_n145), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n118) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U31 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n140), .B(
        LED_RoundFunction2_MCInst1_MC0_n147), .Z(
        LED_RoundFunction2_MCInst1_MC0_n119) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U30 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n126), .B(
        LED_RoundFunction2_MCInst1_MC0_n117), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n140) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U29 ( .A(SubCellOutput2[0]), .B(
        LED_RoundFunction2_MCInst1_MC0_n116), .ZN(
        LED_RoundFunction2_Feedback_45_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U28 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n115), .B(
        LED_RoundFunction2_MCInst1_MC0_n114), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n116) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U27 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n158), .B(SubCellOutput2[61]), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n115) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U26 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n120), .B(
        LED_RoundFunction2_MCInst1_MC0_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n158) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U25 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n113), .B(
        LED_RoundFunction2_MCInst1_MC0_n112), .ZN(
        LED_RoundFunction2_Feedback_44_) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC0_U24 ( .A1(SubCellOutput2[42]), .A2(
        LED_RoundFunction2_MCInst1_MC0_n111), .B1(
        LED_RoundFunction2_MCInst1_MC0_n129), .B2(
        LED_RoundFunction2_MCInst1_MC0_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n112) );
  INV_X1 LED_RoundFunction2_MCInst1_MC0_U23 ( .A(SubCellOutput2[42]), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n138) );
  INV_X1 LED_RoundFunction2_MCInst1_MC0_U22 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n111), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n129) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U21 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n145), .B(
        LED_RoundFunction2_MCInst1_MC0_n154), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n113) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC0_U20 ( .A1(SubCellOutput2[61]), .A2(
        SubCellOutput2[20]), .B1(LED_RoundFunction2_MCInst1_MC0_n110), .B2(
        LED_RoundFunction2_MCInst1_MC0_n132), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n154) );
  INV_X1 LED_RoundFunction2_MCInst1_MC0_U19 ( .A(SubCellOutput2[61]), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n132) );
  INV_X1 LED_RoundFunction2_MCInst1_MC0_U18 ( .A(SubCellOutput2[20]), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n110) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U17 ( .A(SubCellOutput2[3]), .B(
        SubCellOutput2[43]), .Z(LED_RoundFunction2_MCInst1_MC0_n145) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U16 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n111), .B(
        LED_RoundFunction2_MCInst1_MC0_n123), .ZN(
        LED_RoundFunction2_Feedback_63_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U15 ( .A(SubCellOutput2[61]), .B(
        SubCellOutput2[43]), .ZN(LED_RoundFunction2_MCInst1_MC0_n123) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U14 ( .A(SubCellOutput2[22]), .B(
        SubCellOutput2[2]), .Z(LED_RoundFunction2_MCInst1_MC0_n111) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U13 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n120), .B(
        LED_RoundFunction2_MCInst1_MC0_n121), .Z(
        LED_RoundFunction2_Feedback_62_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U12 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n147), .B(SubCellOutput2[60]), .Z(
        LED_RoundFunction2_MCInst1_MC0_n121) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U11 ( .A(SubCellOutput2[1]), .B(
        SubCellOutput2[63]), .Z(LED_RoundFunction2_MCInst1_MC0_n147) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U10 ( .A(SubCellOutput2[42]), .B(
        SubCellOutput2[21]), .Z(LED_RoundFunction2_MCInst1_MC0_n120) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U9 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n117), .B(
        LED_RoundFunction2_MCInst1_MC0_n109), .ZN(
        LED_RoundFunction2_Feedback_61_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U8 ( .A(SubCellOutput2[62]), .B(
        LED_RoundFunction2_MCInst1_MC0_n133), .Z(
        LED_RoundFunction2_MCInst1_MC0_n109) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U7 ( .A(SubCellOutput2[3]), .B(
        SubCellOutput2[63]), .Z(LED_RoundFunction2_MCInst1_MC0_n133) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U6 ( .A(
        LED_RoundFunction2_MCInst1_MC0_n159), .B(
        LED_RoundFunction2_MCInst1_MC0_n125), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n117) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U5 ( .A(SubCellOutput2[23]), .B(
        SubCellOutput2[41]), .Z(LED_RoundFunction2_MCInst1_MC0_n125) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U4 ( .A(SubCellOutput2[0]), .B(
        SubCellOutput2[20]), .Z(LED_RoundFunction2_MCInst1_MC0_n159) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U3 ( .A(SubCellOutput2[3]), .B(
        LED_RoundFunction2_MCInst1_MC0_n114), .ZN(
        LED_RoundFunction2_Feedback_60_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC0_U2 ( .A(SubCellOutput2[23]), .B(
        LED_RoundFunction2_MCInst1_MC0_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC0_n114) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC0_U1 ( .A(SubCellOutput2[62]), .B(
        SubCellOutput2[40]), .Z(LED_RoundFunction2_MCInst1_MC0_n126) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U68 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n160), .B(
        LED_RoundFunction2_MCInst1_MC1_n159), .ZN(
        LED_RoundFunction2_Feedback_11_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U67 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n158), .B(SubCellOutput2[58]), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n160) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U66 ( .A(SubCellOutput2[15]), .B(
        LED_RoundFunction2_MCInst1_MC1_n157), .Z(
        LED_RoundFunction2_Feedback_10_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U65 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n156), .B(
        LED_RoundFunction2_MCInst1_MC1_n155), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n157) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U64 ( .A(SubCellOutput2[17]), .B(
        SubCellOutput2[13]), .ZN(LED_RoundFunction2_MCInst1_MC1_n155) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U63 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n154), .B(SubCellOutput2[37]), .Z(
        LED_RoundFunction2_MCInst1_MC1_n156) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U62 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n153), .B(
        LED_RoundFunction2_MCInst1_MC1_n152), .ZN(
        LED_RoundFunction2_Feedback_9_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U61 ( .A(SubCellOutput2[14]), .B(
        SubCellOutput2[36]), .ZN(LED_RoundFunction2_MCInst1_MC1_n152) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U60 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n151), .B(
        LED_RoundFunction2_MCInst1_MC1_n150), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n153) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U59 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n149), .B(
        LED_RoundFunction2_MCInst1_MC1_n148), .ZN(
        LED_RoundFunction2_Feedback_8_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U58 ( .A(SubCellOutput2[19]), .B(
        LED_RoundFunction2_MCInst1_MC1_n147), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n148) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U57 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n146), .B(
        LED_RoundFunction2_MCInst1_MC1_n150), .Z(
        LED_RoundFunction2_MCInst1_MC1_n149) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U56 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n145), .B(
        LED_RoundFunction2_MCInst1_MC1_n159), .Z(
        LED_RoundFunction2_MCInst1_MC1_n150) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC1_U55 ( .A1(SubCellOutput2[17]), .A2(
        SubCellOutput2[18]), .B1(LED_RoundFunction2_MCInst1_MC1_n144), .B2(
        LED_RoundFunction2_MCInst1_MC1_n143), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n146) );
  INV_X1 LED_RoundFunction2_MCInst1_MC1_U54 ( .A(SubCellOutput2[17]), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n143) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U53 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n142), .B(
        LED_RoundFunction2_MCInst1_MC1_n141), .ZN(
        LED_RoundFunction2_Feedback_27_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U52 ( .A(SubCellOutput2[39]), .B(
        LED_RoundFunction2_MCInst1_MC1_n140), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n141) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U51 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n139), .B(SubCellOutput2[56]), .Z(
        LED_RoundFunction2_MCInst1_MC1_n142) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC1_U50 ( .A1(SubCellOutput2[38]), .A2(
        SubCellOutput2[18]), .B1(LED_RoundFunction2_MCInst1_MC1_n144), .B2(
        LED_RoundFunction2_MCInst1_MC1_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n139) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U49 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n137), .B(
        LED_RoundFunction2_MCInst1_MC1_n136), .ZN(
        LED_RoundFunction2_Feedback_26_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U48 ( .A(SubCellOutput2[36]), .B(
        LED_RoundFunction2_MCInst1_MC1_n135), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n136) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U47 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n134), .B(
        LED_RoundFunction2_MCInst1_MC1_n133), .Z(
        LED_RoundFunction2_MCInst1_MC1_n137) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC1_U46 ( .A1(SubCellOutput2[18]), .A2(
        SubCellOutput2[57]), .B1(LED_RoundFunction2_MCInst1_MC1_n132), .B2(
        LED_RoundFunction2_MCInst1_MC1_n144), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n134) );
  INV_X1 LED_RoundFunction2_MCInst1_MC1_U45 ( .A(SubCellOutput2[18]), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n144) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U44 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n131), .B(
        LED_RoundFunction2_MCInst1_MC1_n151), .ZN(
        LED_RoundFunction2_Feedback_25_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U43 ( .A(SubCellOutput2[59]), .B(
        SubCellOutput2[56]), .ZN(LED_RoundFunction2_MCInst1_MC1_n151) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U42 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n130), .B(
        LED_RoundFunction2_MCInst1_MC1_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n131) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U41 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n128), .B(
        LED_RoundFunction2_MCInst1_MC1_n127), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n130) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U40 ( .A(SubCellOutput2[17]), .B(
        LED_RoundFunction2_MCInst1_MC1_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n127) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U39 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n125), .B(SubCellOutput2[16]), .Z(
        LED_RoundFunction2_MCInst1_MC1_n128) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U38 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n124), .B(
        LED_RoundFunction2_MCInst1_MC1_n123), .ZN(
        LED_RoundFunction2_Feedback_24_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U37 ( .A(SubCellOutput2[12]), .B(
        LED_RoundFunction2_MCInst1_MC1_n122), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n124) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U36 ( .A(SubCellOutput2[14]), .B(
        LED_RoundFunction2_MCInst1_MC1_n122), .ZN(
        LED_RoundFunction2_Feedback_43_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U35 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n135), .B(
        LED_RoundFunction2_MCInst1_MC1_n121), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n122) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U34 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n120), .B(
        LED_RoundFunction2_MCInst1_MC1_n125), .Z(
        LED_RoundFunction2_MCInst1_MC1_n135) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U33 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n119), .B(
        LED_RoundFunction2_MCInst1_MC1_n118), .ZN(
        LED_RoundFunction2_Feedback_42_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U32 ( .A(SubCellOutput2[18]), .B(
        LED_RoundFunction2_MCInst1_MC1_n145), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n118) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U31 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n140), .B(
        LED_RoundFunction2_MCInst1_MC1_n147), .Z(
        LED_RoundFunction2_MCInst1_MC1_n119) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U30 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n126), .B(
        LED_RoundFunction2_MCInst1_MC1_n117), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n140) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U29 ( .A(SubCellOutput2[12]), .B(
        LED_RoundFunction2_MCInst1_MC1_n116), .ZN(
        LED_RoundFunction2_Feedback_41_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U28 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n115), .B(
        LED_RoundFunction2_MCInst1_MC1_n114), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n116) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U27 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n158), .B(SubCellOutput2[57]), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n115) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U26 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n120), .B(
        LED_RoundFunction2_MCInst1_MC1_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n158) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U25 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n113), .B(
        LED_RoundFunction2_MCInst1_MC1_n112), .ZN(
        LED_RoundFunction2_Feedback_40_) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC1_U24 ( .A1(SubCellOutput2[38]), .A2(
        LED_RoundFunction2_MCInst1_MC1_n111), .B1(
        LED_RoundFunction2_MCInst1_MC1_n129), .B2(
        LED_RoundFunction2_MCInst1_MC1_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n112) );
  INV_X1 LED_RoundFunction2_MCInst1_MC1_U23 ( .A(SubCellOutput2[38]), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n138) );
  INV_X1 LED_RoundFunction2_MCInst1_MC1_U22 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n111), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n129) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U21 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n145), .B(
        LED_RoundFunction2_MCInst1_MC1_n154), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n113) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC1_U20 ( .A1(SubCellOutput2[57]), .A2(
        SubCellOutput2[16]), .B1(LED_RoundFunction2_MCInst1_MC1_n110), .B2(
        LED_RoundFunction2_MCInst1_MC1_n132), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n154) );
  INV_X1 LED_RoundFunction2_MCInst1_MC1_U19 ( .A(SubCellOutput2[57]), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n132) );
  INV_X1 LED_RoundFunction2_MCInst1_MC1_U18 ( .A(SubCellOutput2[16]), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n110) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U17 ( .A(SubCellOutput2[15]), .B(
        SubCellOutput2[39]), .Z(LED_RoundFunction2_MCInst1_MC1_n145) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U16 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n111), .B(
        LED_RoundFunction2_MCInst1_MC1_n123), .ZN(
        LED_RoundFunction2_Feedback_59_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U15 ( .A(SubCellOutput2[57]), .B(
        SubCellOutput2[39]), .ZN(LED_RoundFunction2_MCInst1_MC1_n123) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U14 ( .A(SubCellOutput2[18]), .B(
        SubCellOutput2[14]), .Z(LED_RoundFunction2_MCInst1_MC1_n111) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U13 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n120), .B(
        LED_RoundFunction2_MCInst1_MC1_n121), .Z(
        LED_RoundFunction2_Feedback_58_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U12 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n147), .B(SubCellOutput2[56]), .Z(
        LED_RoundFunction2_MCInst1_MC1_n121) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U11 ( .A(SubCellOutput2[13]), .B(
        SubCellOutput2[59]), .Z(LED_RoundFunction2_MCInst1_MC1_n147) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U10 ( .A(SubCellOutput2[38]), .B(
        SubCellOutput2[17]), .Z(LED_RoundFunction2_MCInst1_MC1_n120) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U9 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n117), .B(
        LED_RoundFunction2_MCInst1_MC1_n109), .ZN(
        LED_RoundFunction2_Feedback_57_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U8 ( .A(SubCellOutput2[58]), .B(
        LED_RoundFunction2_MCInst1_MC1_n133), .Z(
        LED_RoundFunction2_MCInst1_MC1_n109) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U7 ( .A(SubCellOutput2[15]), .B(
        SubCellOutput2[59]), .Z(LED_RoundFunction2_MCInst1_MC1_n133) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U6 ( .A(
        LED_RoundFunction2_MCInst1_MC1_n159), .B(
        LED_RoundFunction2_MCInst1_MC1_n125), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n117) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U5 ( .A(SubCellOutput2[19]), .B(
        SubCellOutput2[37]), .Z(LED_RoundFunction2_MCInst1_MC1_n125) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U4 ( .A(SubCellOutput2[12]), .B(
        SubCellOutput2[16]), .Z(LED_RoundFunction2_MCInst1_MC1_n159) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U3 ( .A(SubCellOutput2[15]), .B(
        LED_RoundFunction2_MCInst1_MC1_n114), .ZN(
        LED_RoundFunction2_Feedback_56_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC1_U2 ( .A(SubCellOutput2[19]), .B(
        LED_RoundFunction2_MCInst1_MC1_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC1_n114) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC1_U1 ( .A(SubCellOutput2[58]), .B(
        SubCellOutput2[36]), .Z(LED_RoundFunction2_MCInst1_MC1_n126) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U68 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n160), .B(
        LED_RoundFunction2_MCInst1_MC2_n159), .ZN(
        LED_RoundFunction2_Feedback_7_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U67 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n158), .B(SubCellOutput2[54]), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n160) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U66 ( .A(SubCellOutput2[11]), .B(
        LED_RoundFunction2_MCInst1_MC2_n157), .Z(
        LED_RoundFunction2_Feedback_6_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U65 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n156), .B(
        LED_RoundFunction2_MCInst1_MC2_n155), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n157) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U64 ( .A(SubCellOutput2[29]), .B(
        SubCellOutput2[9]), .ZN(LED_RoundFunction2_MCInst1_MC2_n155) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U63 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n154), .B(SubCellOutput2[33]), .Z(
        LED_RoundFunction2_MCInst1_MC2_n156) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U62 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n153), .B(
        LED_RoundFunction2_MCInst1_MC2_n152), .ZN(
        LED_RoundFunction2_Feedback_5_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U61 ( .A(SubCellOutput2[10]), .B(
        SubCellOutput2[32]), .ZN(LED_RoundFunction2_MCInst1_MC2_n152) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U60 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n151), .B(
        LED_RoundFunction2_MCInst1_MC2_n150), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n153) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U59 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n149), .B(
        LED_RoundFunction2_MCInst1_MC2_n148), .ZN(
        LED_RoundFunction2_Feedback_4_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U58 ( .A(SubCellOutput2[31]), .B(
        LED_RoundFunction2_MCInst1_MC2_n147), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n148) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U57 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n146), .B(
        LED_RoundFunction2_MCInst1_MC2_n150), .Z(
        LED_RoundFunction2_MCInst1_MC2_n149) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U56 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n145), .B(
        LED_RoundFunction2_MCInst1_MC2_n159), .Z(
        LED_RoundFunction2_MCInst1_MC2_n150) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC2_U55 ( .A1(SubCellOutput2[29]), .A2(
        SubCellOutput2[30]), .B1(LED_RoundFunction2_MCInst1_MC2_n144), .B2(
        LED_RoundFunction2_MCInst1_MC2_n143), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n146) );
  INV_X1 LED_RoundFunction2_MCInst1_MC2_U54 ( .A(SubCellOutput2[29]), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n143) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U53 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n142), .B(
        LED_RoundFunction2_MCInst1_MC2_n141), .ZN(
        LED_RoundFunction2_Feedback_23_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U52 ( .A(SubCellOutput2[35]), .B(
        LED_RoundFunction2_MCInst1_MC2_n140), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n141) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U51 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n139), .B(SubCellOutput2[52]), .Z(
        LED_RoundFunction2_MCInst1_MC2_n142) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC2_U50 ( .A1(SubCellOutput2[34]), .A2(
        SubCellOutput2[30]), .B1(LED_RoundFunction2_MCInst1_MC2_n144), .B2(
        LED_RoundFunction2_MCInst1_MC2_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n139) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U49 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n137), .B(
        LED_RoundFunction2_MCInst1_MC2_n136), .ZN(
        LED_RoundFunction2_Feedback_22_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U48 ( .A(SubCellOutput2[32]), .B(
        LED_RoundFunction2_MCInst1_MC2_n135), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n136) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U47 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n134), .B(
        LED_RoundFunction2_MCInst1_MC2_n133), .Z(
        LED_RoundFunction2_MCInst1_MC2_n137) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC2_U46 ( .A1(SubCellOutput2[30]), .A2(
        SubCellOutput2[53]), .B1(LED_RoundFunction2_MCInst1_MC2_n132), .B2(
        LED_RoundFunction2_MCInst1_MC2_n144), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n134) );
  INV_X1 LED_RoundFunction2_MCInst1_MC2_U45 ( .A(SubCellOutput2[30]), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n144) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U44 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n131), .B(
        LED_RoundFunction2_MCInst1_MC2_n151), .ZN(
        LED_RoundFunction2_Feedback_21_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U43 ( .A(SubCellOutput2[55]), .B(
        SubCellOutput2[52]), .ZN(LED_RoundFunction2_MCInst1_MC2_n151) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U42 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n130), .B(
        LED_RoundFunction2_MCInst1_MC2_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n131) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U41 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n128), .B(
        LED_RoundFunction2_MCInst1_MC2_n127), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n130) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U40 ( .A(SubCellOutput2[29]), .B(
        LED_RoundFunction2_MCInst1_MC2_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n127) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U39 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n125), .B(SubCellOutput2[28]), .Z(
        LED_RoundFunction2_MCInst1_MC2_n128) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U38 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n124), .B(
        LED_RoundFunction2_MCInst1_MC2_n123), .ZN(
        LED_RoundFunction2_Feedback_20_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U37 ( .A(SubCellOutput2[8]), .B(
        LED_RoundFunction2_MCInst1_MC2_n122), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n124) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U36 ( .A(SubCellOutput2[10]), .B(
        LED_RoundFunction2_MCInst1_MC2_n122), .ZN(
        LED_RoundFunction2_Feedback_39_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U35 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n135), .B(
        LED_RoundFunction2_MCInst1_MC2_n121), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n122) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U34 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n120), .B(
        LED_RoundFunction2_MCInst1_MC2_n125), .Z(
        LED_RoundFunction2_MCInst1_MC2_n135) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U33 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n119), .B(
        LED_RoundFunction2_MCInst1_MC2_n118), .ZN(
        LED_RoundFunction2_Feedback_38_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U32 ( .A(SubCellOutput2[30]), .B(
        LED_RoundFunction2_MCInst1_MC2_n145), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n118) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U31 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n140), .B(
        LED_RoundFunction2_MCInst1_MC2_n147), .Z(
        LED_RoundFunction2_MCInst1_MC2_n119) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U30 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n126), .B(
        LED_RoundFunction2_MCInst1_MC2_n117), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n140) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U29 ( .A(SubCellOutput2[8]), .B(
        LED_RoundFunction2_MCInst1_MC2_n116), .ZN(
        LED_RoundFunction2_Feedback_37_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U28 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n115), .B(
        LED_RoundFunction2_MCInst1_MC2_n114), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n116) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U27 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n158), .B(SubCellOutput2[53]), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n115) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U26 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n120), .B(
        LED_RoundFunction2_MCInst1_MC2_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n158) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U25 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n113), .B(
        LED_RoundFunction2_MCInst1_MC2_n112), .ZN(
        LED_RoundFunction2_Feedback_36_) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC2_U24 ( .A1(SubCellOutput2[34]), .A2(
        LED_RoundFunction2_MCInst1_MC2_n111), .B1(
        LED_RoundFunction2_MCInst1_MC2_n129), .B2(
        LED_RoundFunction2_MCInst1_MC2_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n112) );
  INV_X1 LED_RoundFunction2_MCInst1_MC2_U23 ( .A(SubCellOutput2[34]), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n138) );
  INV_X1 LED_RoundFunction2_MCInst1_MC2_U22 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n111), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n129) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U21 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n145), .B(
        LED_RoundFunction2_MCInst1_MC2_n154), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n113) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC2_U20 ( .A1(SubCellOutput2[53]), .A2(
        SubCellOutput2[28]), .B1(LED_RoundFunction2_MCInst1_MC2_n110), .B2(
        LED_RoundFunction2_MCInst1_MC2_n132), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n154) );
  INV_X1 LED_RoundFunction2_MCInst1_MC2_U19 ( .A(SubCellOutput2[53]), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n132) );
  INV_X1 LED_RoundFunction2_MCInst1_MC2_U18 ( .A(SubCellOutput2[28]), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n110) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U17 ( .A(SubCellOutput2[11]), .B(
        SubCellOutput2[35]), .Z(LED_RoundFunction2_MCInst1_MC2_n145) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U16 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n111), .B(
        LED_RoundFunction2_MCInst1_MC2_n123), .ZN(
        LED_RoundFunction2_Feedback_55_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U15 ( .A(SubCellOutput2[53]), .B(
        SubCellOutput2[35]), .ZN(LED_RoundFunction2_MCInst1_MC2_n123) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U14 ( .A(SubCellOutput2[30]), .B(
        SubCellOutput2[10]), .Z(LED_RoundFunction2_MCInst1_MC2_n111) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U13 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n120), .B(
        LED_RoundFunction2_MCInst1_MC2_n121), .Z(
        LED_RoundFunction2_Feedback_54_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U12 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n147), .B(SubCellOutput2[52]), .Z(
        LED_RoundFunction2_MCInst1_MC2_n121) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U11 ( .A(SubCellOutput2[9]), .B(
        SubCellOutput2[55]), .Z(LED_RoundFunction2_MCInst1_MC2_n147) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U10 ( .A(SubCellOutput2[34]), .B(
        SubCellOutput2[29]), .Z(LED_RoundFunction2_MCInst1_MC2_n120) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U9 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n117), .B(
        LED_RoundFunction2_MCInst1_MC2_n109), .ZN(
        LED_RoundFunction2_Feedback_53_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U8 ( .A(SubCellOutput2[54]), .B(
        LED_RoundFunction2_MCInst1_MC2_n133), .Z(
        LED_RoundFunction2_MCInst1_MC2_n109) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U7 ( .A(SubCellOutput2[11]), .B(
        SubCellOutput2[55]), .Z(LED_RoundFunction2_MCInst1_MC2_n133) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U6 ( .A(
        LED_RoundFunction2_MCInst1_MC2_n159), .B(
        LED_RoundFunction2_MCInst1_MC2_n125), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n117) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U5 ( .A(SubCellOutput2[31]), .B(
        SubCellOutput2[33]), .Z(LED_RoundFunction2_MCInst1_MC2_n125) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U4 ( .A(SubCellOutput2[8]), .B(
        SubCellOutput2[28]), .Z(LED_RoundFunction2_MCInst1_MC2_n159) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U3 ( .A(SubCellOutput2[11]), .B(
        LED_RoundFunction2_MCInst1_MC2_n114), .ZN(
        LED_RoundFunction2_Feedback_52_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC2_U2 ( .A(SubCellOutput2[31]), .B(
        LED_RoundFunction2_MCInst1_MC2_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC2_n114) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC2_U1 ( .A(SubCellOutput2[54]), .B(
        SubCellOutput2[32]), .Z(LED_RoundFunction2_MCInst1_MC2_n126) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U68 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n160), .B(
        LED_RoundFunction2_MCInst1_MC3_n159), .ZN(
        LED_RoundFunction2_Feedback_3_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U67 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n158), .B(SubCellOutput2[50]), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n160) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U66 ( .A(SubCellOutput2[7]), .B(
        LED_RoundFunction2_MCInst1_MC3_n157), .Z(
        LED_RoundFunction2_Feedback_2_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U65 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n156), .B(
        LED_RoundFunction2_MCInst1_MC3_n155), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n157) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U64 ( .A(SubCellOutput2[25]), .B(
        SubCellOutput2[5]), .ZN(LED_RoundFunction2_MCInst1_MC3_n155) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U63 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n154), .B(SubCellOutput2[45]), .Z(
        LED_RoundFunction2_MCInst1_MC3_n156) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U62 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n153), .B(
        LED_RoundFunction2_MCInst1_MC3_n152), .ZN(
        LED_RoundFunction2_Feedback_1_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U61 ( .A(SubCellOutput2[6]), .B(
        SubCellOutput2[44]), .ZN(LED_RoundFunction2_MCInst1_MC3_n152) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U60 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n151), .B(
        LED_RoundFunction2_MCInst1_MC3_n150), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n153) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U59 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n149), .B(
        LED_RoundFunction2_MCInst1_MC3_n148), .ZN(
        LED_RoundFunction2_Feedback_0_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U58 ( .A(SubCellOutput2[27]), .B(
        LED_RoundFunction2_MCInst1_MC3_n147), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n148) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U57 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n146), .B(
        LED_RoundFunction2_MCInst1_MC3_n150), .Z(
        LED_RoundFunction2_MCInst1_MC3_n149) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U56 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n145), .B(
        LED_RoundFunction2_MCInst1_MC3_n159), .Z(
        LED_RoundFunction2_MCInst1_MC3_n150) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC3_U55 ( .A1(SubCellOutput2[25]), .A2(
        SubCellOutput2[26]), .B1(LED_RoundFunction2_MCInst1_MC3_n144), .B2(
        LED_RoundFunction2_MCInst1_MC3_n143), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n146) );
  INV_X1 LED_RoundFunction2_MCInst1_MC3_U54 ( .A(SubCellOutput2[25]), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n143) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U53 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n142), .B(
        LED_RoundFunction2_MCInst1_MC3_n141), .ZN(
        LED_RoundFunction2_Feedback_19_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U52 ( .A(SubCellOutput2[47]), .B(
        LED_RoundFunction2_MCInst1_MC3_n140), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n141) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U51 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n139), .B(SubCellOutput2[48]), .Z(
        LED_RoundFunction2_MCInst1_MC3_n142) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC3_U50 ( .A1(SubCellOutput2[46]), .A2(
        SubCellOutput2[26]), .B1(LED_RoundFunction2_MCInst1_MC3_n144), .B2(
        LED_RoundFunction2_MCInst1_MC3_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n139) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U49 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n137), .B(
        LED_RoundFunction2_MCInst1_MC3_n136), .ZN(
        LED_RoundFunction2_Feedback_18_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U48 ( .A(SubCellOutput2[44]), .B(
        LED_RoundFunction2_MCInst1_MC3_n135), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n136) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U47 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n134), .B(
        LED_RoundFunction2_MCInst1_MC3_n133), .Z(
        LED_RoundFunction2_MCInst1_MC3_n137) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC3_U46 ( .A1(SubCellOutput2[26]), .A2(
        SubCellOutput2[49]), .B1(LED_RoundFunction2_MCInst1_MC3_n132), .B2(
        LED_RoundFunction2_MCInst1_MC3_n144), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n134) );
  INV_X1 LED_RoundFunction2_MCInst1_MC3_U45 ( .A(SubCellOutput2[26]), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n144) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U44 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n131), .B(
        LED_RoundFunction2_MCInst1_MC3_n151), .ZN(
        LED_RoundFunction2_Feedback_17_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U43 ( .A(SubCellOutput2[51]), .B(
        SubCellOutput2[48]), .ZN(LED_RoundFunction2_MCInst1_MC3_n151) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U42 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n130), .B(
        LED_RoundFunction2_MCInst1_MC3_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n131) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U41 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n128), .B(
        LED_RoundFunction2_MCInst1_MC3_n127), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n130) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U40 ( .A(SubCellOutput2[25]), .B(
        LED_RoundFunction2_MCInst1_MC3_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n127) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U39 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n125), .B(SubCellOutput2[24]), .Z(
        LED_RoundFunction2_MCInst1_MC3_n128) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U38 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n124), .B(
        LED_RoundFunction2_MCInst1_MC3_n123), .ZN(
        LED_RoundFunction2_Feedback_16_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U37 ( .A(SubCellOutput2[4]), .B(
        LED_RoundFunction2_MCInst1_MC3_n122), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n124) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U36 ( .A(SubCellOutput2[6]), .B(
        LED_RoundFunction2_MCInst1_MC3_n122), .ZN(
        LED_RoundFunction2_Feedback_35_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U35 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n135), .B(
        LED_RoundFunction2_MCInst1_MC3_n121), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n122) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U34 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n120), .B(
        LED_RoundFunction2_MCInst1_MC3_n125), .Z(
        LED_RoundFunction2_MCInst1_MC3_n135) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U33 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n119), .B(
        LED_RoundFunction2_MCInst1_MC3_n118), .ZN(
        LED_RoundFunction2_Feedback_34_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U32 ( .A(SubCellOutput2[26]), .B(
        LED_RoundFunction2_MCInst1_MC3_n145), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n118) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U31 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n140), .B(
        LED_RoundFunction2_MCInst1_MC3_n147), .Z(
        LED_RoundFunction2_MCInst1_MC3_n119) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U30 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n126), .B(
        LED_RoundFunction2_MCInst1_MC3_n117), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n140) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U29 ( .A(SubCellOutput2[4]), .B(
        LED_RoundFunction2_MCInst1_MC3_n116), .ZN(
        LED_RoundFunction2_Feedback_33_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U28 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n115), .B(
        LED_RoundFunction2_MCInst1_MC3_n114), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n116) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U27 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n158), .B(SubCellOutput2[49]), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n115) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U26 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n120), .B(
        LED_RoundFunction2_MCInst1_MC3_n129), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n158) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U25 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n113), .B(
        LED_RoundFunction2_MCInst1_MC3_n112), .ZN(
        LED_RoundFunction2_Feedback_32_) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC3_U24 ( .A1(SubCellOutput2[46]), .A2(
        LED_RoundFunction2_MCInst1_MC3_n111), .B1(
        LED_RoundFunction2_MCInst1_MC3_n129), .B2(
        LED_RoundFunction2_MCInst1_MC3_n138), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n112) );
  INV_X1 LED_RoundFunction2_MCInst1_MC3_U23 ( .A(SubCellOutput2[46]), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n138) );
  INV_X1 LED_RoundFunction2_MCInst1_MC3_U22 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n111), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n129) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U21 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n145), .B(
        LED_RoundFunction2_MCInst1_MC3_n154), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n113) );
  AOI22_X1 LED_RoundFunction2_MCInst1_MC3_U20 ( .A1(SubCellOutput2[49]), .A2(
        SubCellOutput2[24]), .B1(LED_RoundFunction2_MCInst1_MC3_n110), .B2(
        LED_RoundFunction2_MCInst1_MC3_n132), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n154) );
  INV_X1 LED_RoundFunction2_MCInst1_MC3_U19 ( .A(SubCellOutput2[49]), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n132) );
  INV_X1 LED_RoundFunction2_MCInst1_MC3_U18 ( .A(SubCellOutput2[24]), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n110) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U17 ( .A(SubCellOutput2[7]), .B(
        SubCellOutput2[47]), .Z(LED_RoundFunction2_MCInst1_MC3_n145) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U16 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n111), .B(
        LED_RoundFunction2_MCInst1_MC3_n123), .ZN(
        LED_RoundFunction2_Feedback_51_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U15 ( .A(SubCellOutput2[49]), .B(
        SubCellOutput2[47]), .ZN(LED_RoundFunction2_MCInst1_MC3_n123) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U14 ( .A(SubCellOutput2[26]), .B(
        SubCellOutput2[6]), .Z(LED_RoundFunction2_MCInst1_MC3_n111) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U13 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n120), .B(
        LED_RoundFunction2_MCInst1_MC3_n121), .Z(
        LED_RoundFunction2_Feedback_50_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U12 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n147), .B(SubCellOutput2[48]), .Z(
        LED_RoundFunction2_MCInst1_MC3_n121) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U11 ( .A(SubCellOutput2[5]), .B(
        SubCellOutput2[51]), .Z(LED_RoundFunction2_MCInst1_MC3_n147) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U10 ( .A(SubCellOutput2[46]), .B(
        SubCellOutput2[25]), .Z(LED_RoundFunction2_MCInst1_MC3_n120) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U9 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n117), .B(
        LED_RoundFunction2_MCInst1_MC3_n109), .ZN(
        LED_RoundFunction2_Feedback_49_) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U8 ( .A(SubCellOutput2[50]), .B(
        LED_RoundFunction2_MCInst1_MC3_n133), .Z(
        LED_RoundFunction2_MCInst1_MC3_n109) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U7 ( .A(SubCellOutput2[7]), .B(
        SubCellOutput2[51]), .Z(LED_RoundFunction2_MCInst1_MC3_n133) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U6 ( .A(
        LED_RoundFunction2_MCInst1_MC3_n159), .B(
        LED_RoundFunction2_MCInst1_MC3_n125), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n117) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U5 ( .A(SubCellOutput2[27]), .B(
        SubCellOutput2[45]), .Z(LED_RoundFunction2_MCInst1_MC3_n125) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U4 ( .A(SubCellOutput2[4]), .B(
        SubCellOutput2[24]), .Z(LED_RoundFunction2_MCInst1_MC3_n159) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U3 ( .A(SubCellOutput2[7]), .B(
        LED_RoundFunction2_MCInst1_MC3_n114), .ZN(
        LED_RoundFunction2_Feedback_48_) );
  XNOR2_X1 LED_RoundFunction2_MCInst1_MC3_U2 ( .A(SubCellOutput2[27]), .B(
        LED_RoundFunction2_MCInst1_MC3_n126), .ZN(
        LED_RoundFunction2_MCInst1_MC3_n114) );
  XOR2_X1 LED_RoundFunction2_MCInst1_MC3_U1 ( .A(SubCellOutput2[50]), .B(
        SubCellOutput2[44]), .Z(LED_RoundFunction2_MCInst1_MC3_n126) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_U1 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n36) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n35) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n34) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n33) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n16), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n43), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n32) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n43) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U12 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n15), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n42), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n31) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n42) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n14), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n41), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n30) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n41) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n13), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n40), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n29) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n28) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n27) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n26) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n25) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n39) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n25), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n26), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n27), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n28), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n29), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n13) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n30), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n14) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n31), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n15) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n32), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n16) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n33), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n34), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n35), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_n36), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[2]), .B(
        SubCellInput2[2]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[2]), .B(
        SubCellInput1[2]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[2]), .B(
        SubCellInput0[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_n1), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_n1) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_n1) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_n1), .CK(clk), .Q(
        SubCellOutput2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[2]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[2]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[2]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U14 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U13 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U12 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U11 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U10 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U9 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U8 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n76) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U7 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n75), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U6 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n75) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_0_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n39) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[2]), .B(
        SubCellInput2[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[2]), .B(
        SubCellInput1[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[2]), .B(
        SubCellInput0[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[5]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[5]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[5]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_0_S2_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U12 ( .B1(RoundFunctionEN), 
        .B2(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_U2 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[2]), .B(
        SubCellInput2[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[2]), .B(
        SubCellInput1[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[2]), .B(
        SubCellInput0[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[9]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[9]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[9]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U12 ( .B1(RoundFunctionEN), 
        .B2(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_U2 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[2]), .B(
        SubCellInput2[14]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[2]), .B(
        SubCellInput1[14]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[2]), .B(
        SubCellInput0[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[15]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[15]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[15]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_1_S2_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U12 ( .B1(RoundFunctionEN), 
        .B2(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_U2 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[2]), .B(
        SubCellInput2[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[2]), .B(
        SubCellInput1[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[2]), .B(
        SubCellInput0[18]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U12 ( .B1(RoundFunctionEN), 
        .B2(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_U2 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[2]), .B(
        SubCellInput2[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[2]), .B(
        SubCellInput1[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[2]), .B(
        SubCellInput0[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_2_S2_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U12 ( .B1(RoundFunctionEN), 
        .B2(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_U2 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[2]), .B(
        SubCellInput2[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[2]), .B(
        SubCellInput1[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[2]), .B(
        SubCellInput0[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[25]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[25]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[25]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[27]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[27]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[27]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U12 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_U2 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[2]), .B(
        SubCellInput2[30]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[2]), .B(
        SubCellInput1[30]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[2]), .B(
        SubCellInput0[30]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[28]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[28]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[28]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[29]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[29]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[29]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[30]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[30]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[30]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[31]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[31]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[31]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_3_S2_G_inst_InstXOR_2__Compression3_n3) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_U1 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U12 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[2]), .B(
        SubCellInput2[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[2]), .B(
        SubCellInput1[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[2]), .B(
        SubCellInput0[34]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[32]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[32]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[32]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[33]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[33]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[33]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[34]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[34]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[34]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[35]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[35]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[35]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U14 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U13 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U12 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U11 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U10 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U9 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U8 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n76) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U7 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n75), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U6 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n75) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_4_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n39) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[2]), .B(
        SubCellInput2[38]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[2]), .B(
        SubCellInput1[38]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[2]), .B(
        SubCellInput0[38]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[36]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[36]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[36]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[37]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[37]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[37]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[38]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[38]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[38]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[39]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[39]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[39]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_4_S2_G_inst_InstXOR_2__Compression3_n3) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_U1 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U14 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U13 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U12 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U11 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U10 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U9 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U8 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n76) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U7 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n75), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U6 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n75) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n39) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[2]), .B(
        SubCellInput2[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[2]), .B(
        SubCellInput1[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[2]), .B(
        SubCellInput0[42]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[40]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[40]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[40]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[41]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[41]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[41]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[42]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[42]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[42]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[43]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[43]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[43]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U12 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[2]), .B(
        SubCellInput2[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[2]), .B(
        SubCellInput1[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[2]), .B(
        SubCellInput0[46]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[44]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[44]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[44]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[45]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[45]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[45]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[46]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[46]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[46]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[47]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[47]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[47]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_5_S2_G_inst_InstXOR_2__Compression3_n3) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_U1 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U12 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[2]), .B(
        SubCellInput2[50]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[2]), .B(
        SubCellInput1[50]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[2]), .B(
        SubCellInput0[50]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[48]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[48]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[48]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[49]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[49]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[49]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[50]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[50]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[50]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[51]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[51]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[51]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U14 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U13 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U12 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U11 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U10 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U9 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U8 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n76) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U7 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n75), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U6 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n75) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_6_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n39) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[2]), .B(
        SubCellInput2[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[2]), .B(
        SubCellInput1[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[2]), .B(
        SubCellInput0[54]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[52]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[52]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[52]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[53]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[53]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[53]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[54]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[54]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[54]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[55]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[55]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[55]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_6_S2_G_inst_InstXOR_2__Compression3_n3) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_U1 ( .A(RoundFunctionEN), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U14 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U13 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U12 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U11 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U10 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U9 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U8 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n76) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U7 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n75), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U6 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n75) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n39) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[2]), .B(
        SubCellInput2[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[2]), .B(
        SubCellInput1[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[2]), .B(
        SubCellInput0[58]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[0]), .B(r[1]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[2]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[2]), .B(r[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[4]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[5]), .B(r[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[5]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[0]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[8]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[10]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[11]), .B(r[10]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .B(r[6]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .B(r[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[12]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[14]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[0]), .B(r[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[14]), .B(r[15]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[16]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_InAff_out3_reg[0]), .B(r[15]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .B(r[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .B(r[16]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[12]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[17]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[56]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[56]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[56]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[19]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[1]), .B(r[18]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[19]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[1]), .B(r[20]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[21]), .B(r[22]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[22]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[1]), .B(r[23]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[25]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[0]), .B(r[24]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[26]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .B(r[25]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[27]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[0]), .B(r[26]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[28]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .B(r[27]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[29]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .B(r[28]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[0]), .B(r[29]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[31]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[1]), .B(r[30]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[31]), .B(r[32]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[33]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[1]), .B(r[32]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[33]), .B(r[34]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[34]), .B(r[35]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[30]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_Q12_1_out2[1]), .B(r[35]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[57]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[57]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[57]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[58]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[58]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[58]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[59]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[59]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[59]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S1_G_inst_InstXOR_2__Compression3_n3) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U18 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n50) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U17 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n49) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U16 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n48) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U15 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n47) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U14 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n62), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n79), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n46) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U13 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n79) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U12 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n61), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n78), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n45) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U11 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n78) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U10 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n60), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n77), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n44) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U9 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n77) );
  OAI21_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U8 ( .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n59), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n76), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n43) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U7 ( .A1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n76) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[0]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n42) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[1]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n41) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[2]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n40) );
  MUX2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[3]), .S(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n39) );
  BUF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_n1), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n75) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n50), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n49), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n48), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n47), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n46), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[0]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n62) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n45), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n61) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n44), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n60) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n43), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .QN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n59) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2_reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n42), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2_reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n41), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2_reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n40), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2_reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_n39), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .QN() );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InputAffine_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[2]), .B(
        SubCellInput2[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InputAffine_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[2]), .B(
        SubCellInput1[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InputAffine_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[2]), .B(
        SubCellInput0[62]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out1[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_U6 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N2) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_n3), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N0) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[1]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_n3) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[26]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N2), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N1), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_N0), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .QN() );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_0__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_0__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[0]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_0__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_0__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_U1 ( .A(
        r[36]), .B(r[37]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_U4 ( .A(
        r[37]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_U2 ( 
        .A(r[38]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_3__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_3__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[3]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_3__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_3__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_U1 ( .A(
        r[38]), .B(r[39]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_U4 ( .A(
        r[39]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_U2 ( 
        .A(r[40]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_6__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_6__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[6]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_6__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_6__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[7]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        r[41]), .B(r[40]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n14)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n11), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n12) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        r[41]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[3]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_U1 ( 
        .A(r[36]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_9__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_9__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[9]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_9__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_U1 ( 
        .A(r[42]), .B(r[43]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_10__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[11]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_U4 ( 
        .A(r[43]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_U2 ( 
        .A(r[44]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n11)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_11__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_12__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_12__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[12]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_12__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_U1 ( 
        .A(r[44]), .B(r[45]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_13__CF_Inst_n8) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[14]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_U5 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_U4 ( 
        .A(r[45]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n13), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n13)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_U2 ( 
        .A(r[46]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_14__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_15__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_15__CF_Inst_n3), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[15]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_15__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_U2 ( 
        .A(r[47]), .B(r[46]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n10), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n9), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n11)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[4]), .B(r[42]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n10) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[5]), .B(r[47]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_17__CF_Inst_n12) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[18]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_U3 ( 
        .A(r[48]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_19__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_U7 ( 
        .A(r[50]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[20]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[0]), .B(r[49]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n15) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_20__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[21]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n12), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_U3 ( 
        .A(r[50]), .B(r[51]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n12) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n14)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_22__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_U7 ( 
        .A(r[52]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n20), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[23]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n19), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n18), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n20)
         );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n17), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n18)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n17) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n16), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n19)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_InAff_out3_reg[0]), .B(r[51]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n15)
         );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_23__CF_Inst_n16) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_n6), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[24]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_U2 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_n5), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_U1 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n17), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n16), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[25]) );
  OAI211_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_U5 ( 
        .C1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .C2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n15), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n16)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[5]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n15) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_U3 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n14), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n13), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n17)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .B(r[53]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n13) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[4]), .B(r[52]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_25__CF_Inst_n14) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_U6 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n15), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n14), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n13), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n12), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n14)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_U4 ( 
        .A(r[48]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[6]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n12) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_U3 ( 
        .A(r[53]), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_rs1[7]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n13) );
  AOI22_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[2]), .B1(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[1]), .B2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n11), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n15)
         );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_rs2[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_Inst_26__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[5]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[8]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[0]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[11]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[14]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[17]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[20]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[23]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[26]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_F_inst_InstXOR_2__Compression3_n3) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_U5 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_N0) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_U4 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[0]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_N1) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[0]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_n2) );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_areg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_n2), .CK(clk), .Q(
        SubCellOutput2[60]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_areg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_N1), .CK(clk), .Q(
        SubCellOutput0[60]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_areg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_N0), .CK(clk), .Q(
        SubCellOutput1[60]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[26]), .QN() );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_0__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[0]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_U6 ( .A(
        r[55]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[1]), .B(r[54]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_1__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[2]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(
        r[55]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_2__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_3__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[3]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_U6 ( .A(
        r[57]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[1]), .B(r[56]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_4__CF_Inst_n11) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[5]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(
        r[57]), .B(r[58]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_5__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_6__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[6]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[7]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_U2 ( .A(
        r[58]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_7__CF_Inst_n6) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        r[54]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[8]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[1]), .B(r[59]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_8__CF_Inst_n11) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_9__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[9]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_U6 ( 
        .A(r[61]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[0]), .B(r[60]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_10__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_U5 ( 
        .A(r[62]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[11]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .B(r[61]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_11__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_12__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[12]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_U6 ( 
        .A(r[63]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[0]), .B(r[62]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_13__CF_Inst_n11) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_U5 ( 
        .A(r[64]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[14]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .B(r[63]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_14__CF_Inst_n8) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_15__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[15]) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_U5 ( 
        .A(r[65]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n9), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n9)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[1]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n7) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .B(r[64]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_16__CF_Inst_n8) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_U6 ( 
        .A(r[60]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n12), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_U5 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n11), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n10), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n12)
         );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_U4 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n10) );
  INV_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n9) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[0]), .B(r[65]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_17__CF_Inst_n11) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_18__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[18]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_U5 ( 
        .A(r[67]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[1]), .B(r[66]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_19__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[20]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_U2 ( 
        .A(r[67]), .B(r[68]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_20__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_21__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[21]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_U5 ( 
        .A(r[69]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[1]), .B(r[68]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_22__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[23]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out3[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_U2 ( 
        .A(r[69]), .B(r[70]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_23__CF_Inst_n6) );
  AND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_24__CF_Inst_U2 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[24]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_n6), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_n5), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[25]) );
  NAND2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[2]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[3]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_n5) );
  XOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_U2 ( 
        .A(r[70]), .B(r[71]), .Z(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_25__CF_Inst_n6) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_U5 ( 
        .A(r[66]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n9), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_U4 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n8), 
        .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n7), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n9)
         );
  NOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_U3 ( 
        .A1(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out1[3]), .A2(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[2]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n7) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_U2 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_Q12_1_out2[1]), .B(r[71]), 
        .ZN(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_Inst_26__CF_Inst_n8)
         );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[2]), .ZN(
        SubCellOutput0[61]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[0]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[1]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[5]), .ZN(
        SubCellOutput1[61]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[3]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[4]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[8]), .ZN(
        SubCellOutput2[61]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[6]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[7]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[11]), .ZN(
        SubCellOutput0[62]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[9]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[10]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[14]), .ZN(
        SubCellOutput1[62]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[12]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[13]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[17]), .ZN(
        SubCellOutput2[62]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[15]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[16]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression1_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression1_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[20]), .ZN(
        SubCellOutput0[63]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression1_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[18]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[19]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression2_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression2_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[23]), .ZN(
        SubCellOutput1[63]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression2_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[21]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[22]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression3_U2 ( 
        .A(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression3_n3), .B(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[26]), .ZN(
        SubCellOutput2[63]) );
  XNOR2_X1 Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression3_U1 ( 
        .A(Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[24]), .B(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_CF_Reg[25]), .ZN(
        Inst_SubCell_Multi_Inst_TwoSbox_7_S2_G_inst_InstXOR_2__Compression3_n3) );
  AOI22_X1 LED128_Controller_Inst_U48 ( .A1(LED128_Controller_Inst_n48), .A2(
        LED128_Controller_Inst_n3), .B1(LED128_Controller_Inst_n38), .B2(
        LED128_Controller_Inst_n19), .ZN(LED128_Controller_Inst_n46) );
  INV_X1 LED128_Controller_Inst_U47 ( .A(FSM[5]), .ZN(
        LED128_Controller_Inst_n38) );
  AOI22_X1 LED128_Controller_Inst_U46 ( .A1(LED128_Controller_Inst_n48), .A2(
        LED128_Controller_Inst_n15), .B1(LED128_Controller_Inst_n37), .B2(
        LED128_Controller_Inst_n19), .ZN(LED128_Controller_Inst_n45) );
  AOI22_X1 LED128_Controller_Inst_U45 ( .A1(LED128_Controller_Inst_n48), .A2(
        LED128_Controller_Inst_n12), .B1(LED128_Controller_Inst_n36), .B2(
        LED128_Controller_Inst_n19), .ZN(LED128_Controller_Inst_n44) );
  AOI22_X1 LED128_Controller_Inst_U44 ( .A1(LED128_Controller_Inst_n48), .A2(
        LED128_Controller_Inst_n9), .B1(LED128_Controller_Inst_n35), .B2(
        LED128_Controller_Inst_n19), .ZN(LED128_Controller_Inst_n43) );
  AOI22_X1 LED128_Controller_Inst_U43 ( .A1(LED128_Controller_Inst_n48), .A2(
        LED128_Controller_Inst_n7), .B1(LED128_Controller_Inst_n34), .B2(
        LED128_Controller_Inst_n19), .ZN(LED128_Controller_Inst_n42) );
  AOI22_X1 LED128_Controller_Inst_U42 ( .A1(LED128_Controller_Inst_n48), .A2(
        LED128_Controller_Inst_n6), .B1(LED128_Controller_Inst_n33), .B2(
        LED128_Controller_Inst_n19), .ZN(LED128_Controller_Inst_n41) );
  NOR2_X1 LED128_Controller_Inst_U41 ( .A1(rst), .A2(
        LED128_Controller_Inst_n40), .ZN(LED128_Controller_Inst_n2) );
  NOR2_X1 LED128_Controller_Inst_U40 ( .A1(rst), .A2(
        LED128_Controller_Inst_n39), .ZN(LED128_Controller_Inst_n1) );
  NOR4_X1 LED128_Controller_Inst_U39 ( .A1(FSM[4]), .A2(
        LED128_Controller_Inst_n32), .A3(LED128_Controller_Inst_n31), .A4(
        LED128_Controller_Inst_n30), .ZN(done) );
  OAI221_X1 LED128_Controller_Inst_U38 ( .B1(FSM[2]), .B2(FSM[0]), .C1(
        LED128_Controller_Inst_n35), .C2(FSM[4]), .A(
        LED128_Controller_Inst_n29), .ZN(SelKey) );
  OAI22_X1 LED128_Controller_Inst_U37 ( .A1(LED128_Controller_Inst_n28), .A2(
        LED128_Controller_Inst_n27), .B1(LED128_Controller_Inst_n26), .B2(
        LED128_Controller_Inst_n31), .ZN(LED128_Controller_Inst_n29) );
  INV_X1 LED128_Controller_Inst_U36 ( .A(LED128_Controller_Inst_n25), .ZN(
        LED128_Controller_Inst_n31) );
  XOR2_X1 LED128_Controller_Inst_U35 ( .A(LED128_Controller_Inst_n26), .B(
        LED128_Controller_Inst_n36), .Z(LED128_Controller_Inst_n27) );
  NAND2_X1 LED128_Controller_Inst_U34 ( .A1(FSM[0]), .A2(FSM[2]), .ZN(
        LED128_Controller_Inst_n26) );
  NAND2_X1 LED128_Controller_Inst_U33 ( .A1(LED128_Controller_Inst_n34), .A2(
        LED128_Controller_Inst_n24), .ZN(LED128_Controller_Inst_n28) );
  INV_X1 LED128_Controller_Inst_U32 ( .A(FSM[2]), .ZN(
        LED128_Controller_Inst_n35) );
  AOI22_X1 LED128_Controller_Inst_U31 ( .A1(LED128_Controller_Inst_n18), .A2(
        LED128_Controller_Inst_n25), .B1(LED128_Controller_Inst_n17), .B2(
        LED128_Controller_Inst_n34), .ZN(LED128_Controller_Inst_n20) );
  AOI221_X1 LED128_Controller_Inst_U30 ( .B1(LED128_Controller_Inst_n16), .B2(
        FSM[1]), .C1(LED128_Controller_Inst_n14), .C2(
        LED128_Controller_Inst_n36), .A(LED128_Controller_Inst_n13), .ZN(
        LED128_Controller_Inst_n17) );
  NAND2_X1 LED128_Controller_Inst_U29 ( .A1(FSM[2]), .A2(FSM[4]), .ZN(
        LED128_Controller_Inst_n13) );
  INV_X1 LED128_Controller_Inst_U28 ( .A(FSM[1]), .ZN(
        LED128_Controller_Inst_n36) );
  INV_X1 LED128_Controller_Inst_U27 ( .A(LED128_Controller_Inst_n14), .ZN(
        LED128_Controller_Inst_n16) );
  NAND2_X1 LED128_Controller_Inst_U26 ( .A1(FSM[5]), .A2(
        LED128_Controller_Inst_n3), .ZN(LED128_Controller_Inst_n14) );
  NOR2_X1 LED128_Controller_Inst_U25 ( .A1(LED128_Controller_Inst_n34), .A2(
        FSM[5]), .ZN(LED128_Controller_Inst_n25) );
  OAI33_X1 LED128_Controller_Inst_U24 ( .A1(FSM[0]), .A2(FSM[4]), .A3(
        LED128_Controller_Inst_n30), .B1(LED128_Controller_Inst_n37), .B2(
        LED128_Controller_Inst_n33), .B3(LED128_Controller_Inst_n11), .ZN(
        LED128_Controller_Inst_n18) );
  OAI211_X1 LED128_Controller_Inst_U23 ( .C1(FSM[4]), .C2(
        LED128_Controller_Inst_n34), .A(FSM[0]), .B(LED128_Controller_Inst_n24), .ZN(LED128_Controller_Inst_n21) );
  INV_X1 LED128_Controller_Inst_U22 ( .A(LED128_Controller_Inst_n23), .ZN(
        LED128_Controller_Inst_n24) );
  INV_X1 LED128_Controller_Inst_U21 ( .A(LED128_Controller_Inst_n11), .ZN(
        LED128_Controller_Inst_n30) );
  NOR2_X1 LED128_Controller_Inst_U20 ( .A1(FSM[2]), .A2(FSM[1]), .ZN(
        LED128_Controller_Inst_n11) );
  NOR3_X1 LED128_Controller_Inst_U19 ( .A1(rst), .A2(LED128_Controller_Inst_n3), .A3(LED128_Controller_Inst_n8), .ZN(LED128_Controller_Inst_n32) );
  NOR2_X1 LED128_Controller_Inst_U18 ( .A1(rst), .A2(
        LED128_Controller_Inst_n15), .ZN(FSM[1]) );
  NOR2_X1 LED128_Controller_Inst_U17 ( .A1(rst), .A2(LED128_Controller_Inst_n7), .ZN(FSM[4]) );
  INV_X1 LED128_Controller_Inst_U16 ( .A(FSM[4]), .ZN(
        LED128_Controller_Inst_n33) );
  NOR2_X1 LED128_Controller_Inst_U15 ( .A1(rst), .A2(LED128_Controller_Inst_n6), .ZN(FSM[5]) );
  NOR2_X1 LED128_Controller_Inst_U14 ( .A1(LED128_Controller_Inst_n33), .A2(
        FSM[5]), .ZN(LED128_Controller_Inst_n23) );
  NOR2_X1 LED128_Controller_Inst_U13 ( .A1(rst), .A2(
        LED128_Controller_Inst_n12), .ZN(FSM[2]) );
  AOI21_X1 LED128_Controller_Inst_U12 ( .B1(LED128_Controller_Inst_n3), .B2(
        FSM[5]), .A(LED128_Controller_Inst_n32), .ZN(FSM[0]) );
  INV_X1 LED128_Controller_Inst_U11 ( .A(FSM[0]), .ZN(
        LED128_Controller_Inst_n37) );
  NOR2_X1 LED128_Controller_Inst_U10 ( .A1(FSM[2]), .A2(
        LED128_Controller_Inst_n37), .ZN(LED128_Controller_Inst_n22) );
  NOR2_X1 LED128_Controller_Inst_U9 ( .A1(rst), .A2(LED128_Controller_Inst_n9), 
        .ZN(FSM[3]) );
  INV_X1 LED128_Controller_Inst_U8 ( .A(FSM[3]), .ZN(
        LED128_Controller_Inst_n34) );
  NAND4_X1 LED128_Controller_Inst_U7 ( .A1(FSM[1]), .A2(
        LED128_Controller_Inst_n23), .A3(LED128_Controller_Inst_n22), .A4(
        LED128_Controller_Inst_n34), .ZN(RoundFunctionEN) );
  OAI21_X1 LED128_Controller_Inst_U6 ( .B1(LED128_Controller_Inst_n30), .B2(
        LED128_Controller_Inst_n21), .A(LED128_Controller_Inst_n20), .ZN(
        AddKey) );
  INV_X1 LED128_Controller_Inst_U5 ( .A(rst), .ZN(LED128_Controller_Inst_n10)
         );
  NAND2_X1 LED128_Controller_Inst_U4 ( .A1(LED128_Controller_Inst_n47), .A2(
        LED128_Controller_Inst_n10), .ZN(LED128_Controller_Inst_n19) );
  INV_X1 LED128_Controller_Inst_U3 ( .A(LED128_Controller_Inst_n19), .ZN(
        LED128_Controller_Inst_n48) );
  DFF_X1 LED128_Controller_Inst_FSM_EN_reg_reg_1_ ( .D(
        LED128_Controller_Inst_n1), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n40) );
  DFF_X1 LED128_Controller_Inst_FSM_EN_reg_reg_2_ ( .D(
        LED128_Controller_Inst_n2), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n47) );
  DFF_X1 LED128_Controller_Inst_FSM_reg_output_reg_4_ ( .D(
        LED128_Controller_Inst_n41), .CK(clk), .Q(LED128_Controller_Inst_n8), 
        .QN(LED128_Controller_Inst_n6) );
  DFF_X1 LED128_Controller_Inst_FSM_reg_output_reg_3_ ( .D(
        LED128_Controller_Inst_n42), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n7) );
  DFF_X1 LED128_Controller_Inst_FSM_reg_output_reg_2_ ( .D(
        LED128_Controller_Inst_n43), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n9) );
  DFF_X1 LED128_Controller_Inst_FSM_reg_output_reg_1_ ( .D(
        LED128_Controller_Inst_n44), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n12) );
  DFF_X1 LED128_Controller_Inst_FSM_reg_output_reg_0_ ( .D(
        LED128_Controller_Inst_n45), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n15) );
  DFF_X1 LED128_Controller_Inst_FSM_reg_output_reg_5_ ( .D(
        LED128_Controller_Inst_n46), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n3) );
  DFF_X1 LED128_Controller_Inst_FSM_EN_reg_reg_0_ ( .D(
        LED128_Controller_Inst_n19), .CK(clk), .Q(), .QN(
        LED128_Controller_Inst_n39) );
endmodule

