
module circuit ( ClkxCI, RstxBI, PTxDI, KxDI, PRNGQ, StartxSI, DonexSO, CxDO
 );
  input [23:0] PTxDI;
  input [23:0] KxDI;
  input [51:0] PRNGQ;
  output [23:0] CxDO;
  input ClkxCI, RstxBI, StartxSI;
  output DonexSO;
  wire   disableKeyRegsxS, ClkKeyRegxC, StateKEYSCHEDULExS, showRCONxS,
         StateKEYADDITION1o3xS, LastRoundxS, doMixColumnsxS, n170, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, aes_ctrl_lsfr_23_cycles_1_n24,
         aes_ctrl_lsfr_23_cycles_1_n23, aes_ctrl_lsfr_23_cycles_1_n22,
         aes_ctrl_lsfr_23_cycles_1_n21, aes_ctrl_lsfr_23_cycles_1_n20,
         aes_ctrl_lsfr_23_cycles_1_n19, aes_ctrl_lsfr_23_cycles_1_n18,
         aes_ctrl_lsfr_23_cycles_1_n17, aes_ctrl_lsfr_23_cycles_1_n16,
         aes_ctrl_lsfr_23_cycles_1_n15, aes_ctrl_lsfr_23_cycles_1_n14,
         aes_ctrl_lsfr_23_cycles_1_n13, aes_ctrl_lsfr_23_cycles_1_n11,
         aes_ctrl_lsfr_23_cycles_1_n10, aes_ctrl_lsfr_23_cycles_1_n8,
         aes_ctrl_lsfr_23_cycles_1_n7, aes_ctrl_lsfr_23_cycles_1_n5,
         aes_ctrl_lsfr_23_cycles_1_n3, aes_ctrl_lsfr_23_cycles_1_n1,
         aes_ctrl_lsfr_23_cycles_1_n39, aes_ctrl_lsfr_23_cycles_1_n38,
         aes_ctrl_lsfr_23_cycles_1_n37, aes_ctrl_lsfr_23_cycles_1_n36,
         aes_ctrl_lsfr_23_cycles_1_n35, aes_ctrl_lsfr_23_cycles_1_n12,
         aes_ctrl_lsfr_23_cycles_1_n9, aes_ctrl_lsfr_23_cycles_1_n6,
         aes_ctrl_lsfr_23_cycles_1_n4, aes_ctrl_lsfr_23_cycles_1_n2,
         aes_ctrl_lsfr_23_cycles_1_N83, aes_ctrl_lsfr_23_cycles_1_N66,
         aes_ctrl_lsfr_23_cycles_1_N16, rcon_1_n43, rcon_1_n42, rcon_1_n41,
         rcon_1_n40, rcon_1_n39, rcon_1_n38, rcon_1_n37, rcon_1_n36,
         rcon_1_n34, rcon_1_n33, rcon_1_n32, rcon_1_n31, rcon_1_n30,
         rcon_1_n29, rcon_1_n28, rcon_1_n16, rcon_1_n15, rcon_1_n14,
         rcon_1_n13, rcon_1_n12, rcon_1_n11, rcon_1_n35, rcon_1_n26,
         rcon_1_n25, rcon_1_n24, rcon_1_n23, rcon_1_n22, rcon_1_n21,
         rcon_1_n20, rcon_1_n19, rcon_1_n18, rcon_1_n17, rcon_1_n9, rcon_1_n4,
         SBOX_Zl_f1_0_, SBOX_Zl_f1_1_, SBOX_Zl_f1_3_, SBOX_Zl_f1_4_,
         SBOX_Zl_f1_5_, SBOX_Zl_f1_7_, SBOX_Zl_f1_8_, SBOX_Zl_f1_9_,
         SBOX_Zl_f1_11_, SBOX_Inst_f1_linearMapping_n32,
         SBOX_Inst_f1_linearMapping_n31, SBOX_Inst_f1_linearMapping_n30,
         SBOX_Inst_f1_linearMapping_n29, SBOX_Inst_f1_linearMapping_n28,
         SBOX_Inst_f1_linearMapping_n27, SBOX_Inst_f1_linearMapping_n26,
         SBOX_Inst_f1_linearMapping_n25, SBOX_Inst_f1_linearMapping_n24,
         SBOX_Inst_f1_linearMapping_n23, SBOX_Inst_f1_linearMapping_n22,
         SBOX_Inst_f1_linearMapping_n21, SBOX_Inst_f1_linearMapping_n20,
         SBOX_Inst_f1_linearMapping_n19, SBOX_Inst_f1_linearMapping_n18,
         SBOX_Inst_f1_linearMapping_n17, SBOX_Inst_f1_linearMapping_n16,
         SBOX_Inst_f1_linearMapping_n15, SBOX_Inst_f1_linearMapping_n14,
         SBOX_Inst_f1_linearMapping_n13, SBOX_Inst_f1_linearMapping_n12,
         SBOX_Inst_f1_phpplmul_himul_n172, SBOX_Inst_f1_phpplmul_himul_n171,
         SBOX_Inst_f1_phpplmul_himul_n170, SBOX_Inst_f1_phpplmul_himul_n169,
         SBOX_Inst_f1_phpplmul_himul_n168, SBOX_Inst_f1_phpplmul_himul_n167,
         SBOX_Inst_f1_phpplmul_himul_n166, SBOX_Inst_f1_phpplmul_himul_n165,
         SBOX_Inst_f1_phpplmul_himul_n164, SBOX_Inst_f1_phpplmul_himul_n163,
         SBOX_Inst_f1_phpplmul_himul_n162, SBOX_Inst_f1_phpplmul_himul_n161,
         SBOX_Inst_f1_phpplmul_himul_n160, SBOX_Inst_f1_phpplmul_himul_n159,
         SBOX_Inst_f1_phpplmul_himul_n158, SBOX_Inst_f1_phpplmul_himul_n157,
         SBOX_Inst_f1_phpplmul_himul_n156, SBOX_Inst_f1_phpplmul_himul_n155,
         SBOX_Inst_f1_phpplmul_himul_n154, SBOX_Inst_f1_phpplmul_himul_n153,
         SBOX_Inst_f1_phpplmul_himul_n152, SBOX_Inst_f1_phpplmul_himul_n151,
         SBOX_Inst_f1_phpplmul_himul_n150, SBOX_Inst_f1_phpplmul_himul_n149,
         SBOX_Inst_f1_phpplmul_himul_n148, SBOX_Inst_f1_phpplmul_himul_n147,
         SBOX_Inst_f1_phpplmul_himul_n146, SBOX_Inst_f1_phpplmul_himul_n145,
         SBOX_Inst_f1_phpplmul_himul_n144, SBOX_Inst_f1_phpplmul_himul_n143,
         SBOX_Inst_f1_phpplmul_himul_n142, SBOX_Inst_f1_phpplmul_himul_n141,
         SBOX_Inst_f1_phpplmul_himul_n140, SBOX_Inst_f1_phpplmul_himul_n139,
         SBOX_Inst_f1_phpplmul_himul_n138, SBOX_Inst_f1_phpplmul_himul_n137,
         SBOX_Inst_f1_phpplmul_himul_n136, SBOX_Inst_f1_phpplmul_himul_n135,
         SBOX_Inst_f1_phpplmul_himul_n134, SBOX_Inst_f1_phpplmul_himul_n133,
         SBOX_Inst_f1_phpplmul_himul_n132, SBOX_Inst_f1_phpplmul_himul_n131,
         SBOX_Inst_f1_phpplmul_himul_n130, SBOX_Inst_f1_phpplmul_himul_n129,
         SBOX_Inst_f1_phpplmul_himul_n128, SBOX_Inst_f1_phpplmul_himul_n127,
         SBOX_Inst_f1_phpplmul_himul_n126, SBOX_Inst_f1_phpplmul_himul_n125,
         SBOX_Inst_f1_phpplmul_himul_n124, SBOX_Inst_f1_phpplmul_himul_n123,
         SBOX_Inst_f1_phpplmul_himul_n122, SBOX_Inst_f1_phpplmul_himul_n121,
         SBOX_Inst_f1_phpplmul_himul_n120, SBOX_Inst_f1_phpplmul_himul_n119,
         SBOX_Inst_f1_phpplmul_himul_n118, SBOX_Inst_f1_phpplmul_himul_n117,
         SBOX_Inst_f1_phpplmul_himul_n116, SBOX_Inst_f1_phpplmul_himul_n115,
         SBOX_Inst_f1_phpplmul_himul_n114, SBOX_Inst_f1_phpplmul_himul_n113,
         SBOX_Inst_f1_phpplmul_himul_n112, SBOX_Inst_f1_phpplmul_himul_n111,
         SBOX_Inst_f1_phpplmul_himul_n110, SBOX_Inst_f1_phpplmul_himul_n109,
         SBOX_Inst_f1_phpplmul_himul_n108, SBOX_Inst_f1_phpplmul_himul_n107,
         SBOX_Inst_f1_phpplmul_himul_n106, SBOX_Inst_f1_phpplmul_himul_n105,
         SBOX_Inst_f1_phpplmul_himul_n104, SBOX_Inst_f1_phpplmul_himul_n103,
         SBOX_Inst_f1_phpplmul_himul_n102, SBOX_Inst_f1_phpplmul_himul_n101,
         SBOX_Inst_f1_phpplmul_himul_n100, SBOX_Inst_f1_phpplmul_himul_n99,
         SBOX_Inst_f1_phpplmul_himul_n98, SBOX_Inst_f1_phpplmul_himul_n97,
         SBOX_Inst_f1_phpplmul_himul_n96, SBOX_Inst_f1_phpplmul_himul_n95,
         SBOX_Inst_f1_phpplmul_himul_n94, SBOX_Inst_f1_phpplmul_himul_n93,
         SBOX_Inst_f1_phpplmul_himul_n92, SBOX_Inst_f1_phpplmul_himul_n91,
         SBOX_Inst_f1_phpplmul_himul_n90, SBOX_Inst_f1_phpplmul_himul_n89,
         SBOX_Inst_f1_phpplmul_himul_n88, SBOX_Inst_f1_phpplmul_himul_n87,
         SBOX_Inst_f1_phpplmul_himul_n86, SBOX_Inst_f1_phpplmul_himul_n85,
         SBOX_Inst_f1_phpplmul_himul_n84, SBOX_Inst_f1_phpplmul_himul_n83,
         SBOX_Inst_f1_phpplmul_himul_n82, SBOX_Inst_f1_phpplmul_himul_n81,
         SBOX_Inst_f1_phpplmul_himul_n80, SBOX_Inst_f1_phpplmul_himul_n79,
         SBOX_Inst_f1_phpplmul_himul_n78, SBOX_Inst_f1_phpplmul_himul_n77,
         SBOX_Inst_f1_phpplmul_himul_n76,
         SBOX_Inst_f1_phpplmul_AddNewMaskph_n6,
         SBOX_Inst_f1_phpplmul_AddNewMaskph_n5,
         SBOX_Inst_f1_phpplmul_summul_n300, SBOX_Inst_f1_phpplmul_summul_n299,
         SBOX_Inst_f1_phpplmul_summul_n298, SBOX_Inst_f1_phpplmul_summul_n297,
         SBOX_Inst_f1_phpplmul_summul_n296, SBOX_Inst_f1_phpplmul_summul_n295,
         SBOX_Inst_f1_phpplmul_summul_n294, SBOX_Inst_f1_phpplmul_summul_n293,
         SBOX_Inst_f1_phpplmul_summul_n292, SBOX_Inst_f1_phpplmul_summul_n291,
         SBOX_Inst_f1_phpplmul_summul_n290, SBOX_Inst_f1_phpplmul_summul_n289,
         SBOX_Inst_f1_phpplmul_summul_n288, SBOX_Inst_f1_phpplmul_summul_n287,
         SBOX_Inst_f1_phpplmul_summul_n286, SBOX_Inst_f1_phpplmul_summul_n285,
         SBOX_Inst_f1_phpplmul_summul_n284, SBOX_Inst_f1_phpplmul_summul_n283,
         SBOX_Inst_f1_phpplmul_summul_n282, SBOX_Inst_f1_phpplmul_summul_n281,
         SBOX_Inst_f1_phpplmul_summul_n280, SBOX_Inst_f1_phpplmul_summul_n279,
         SBOX_Inst_f1_phpplmul_summul_n278, SBOX_Inst_f1_phpplmul_summul_n277,
         SBOX_Inst_f1_phpplmul_summul_n276, SBOX_Inst_f1_phpplmul_summul_n275,
         SBOX_Inst_f1_phpplmul_summul_n274, SBOX_Inst_f1_phpplmul_summul_n273,
         SBOX_Inst_f1_phpplmul_summul_n272, SBOX_Inst_f1_phpplmul_summul_n271,
         SBOX_Inst_f1_phpplmul_summul_n270, SBOX_Inst_f1_phpplmul_summul_n269,
         SBOX_Inst_f1_phpplmul_summul_n268, SBOX_Inst_f1_phpplmul_summul_n267,
         SBOX_Inst_f1_phpplmul_summul_n266, SBOX_Inst_f1_phpplmul_summul_n265,
         SBOX_Inst_f1_phpplmul_summul_n264, SBOX_Inst_f1_phpplmul_summul_n263,
         SBOX_Inst_f1_phpplmul_summul_n262, SBOX_Inst_f1_phpplmul_summul_n261,
         SBOX_Inst_f1_phpplmul_summul_n260, SBOX_Inst_f1_phpplmul_summul_n259,
         SBOX_Inst_f1_phpplmul_summul_n258, SBOX_Inst_f1_phpplmul_summul_n257,
         SBOX_Inst_f1_phpplmul_summul_n256, SBOX_Inst_f1_phpplmul_summul_n255,
         SBOX_Inst_f1_phpplmul_summul_n254, SBOX_Inst_f1_phpplmul_summul_n253,
         SBOX_Inst_f1_phpplmul_summul_n252, SBOX_Inst_f1_phpplmul_summul_n251,
         SBOX_Inst_f1_phpplmul_summul_n250, SBOX_Inst_f1_phpplmul_summul_n249,
         SBOX_Inst_f1_phpplmul_summul_n248, SBOX_Inst_f1_phpplmul_summul_n247,
         SBOX_Inst_f1_phpplmul_summul_n246, SBOX_Inst_f1_phpplmul_summul_n245,
         SBOX_Inst_f1_phpplmul_summul_n244, SBOX_Inst_f1_phpplmul_summul_n243,
         SBOX_Inst_f1_phpplmul_summul_n242, SBOX_Inst_f1_phpplmul_summul_n241,
         SBOX_Inst_f1_phpplmul_summul_n240, SBOX_Inst_f1_phpplmul_summul_n239,
         SBOX_Inst_f1_phpplmul_summul_n238, SBOX_Inst_f1_phpplmul_summul_n237,
         SBOX_Inst_f1_phpplmul_summul_n236, SBOX_Inst_f1_phpplmul_summul_n235,
         SBOX_Inst_f1_phpplmul_summul_n234, SBOX_Inst_f1_phpplmul_summul_n233,
         SBOX_Inst_f1_phpplmul_summul_n232, SBOX_Inst_f1_phpplmul_summul_n231,
         SBOX_Inst_f1_phpplmul_summul_n230, SBOX_Inst_f1_phpplmul_summul_n229,
         SBOX_Inst_f1_phpplmul_summul_n228, SBOX_Inst_f1_phpplmul_summul_n227,
         SBOX_Inst_f1_phpplmul_summul_n226, SBOX_Inst_f1_phpplmul_summul_n225,
         SBOX_Inst_f1_phpplmul_summul_n224, SBOX_Inst_f1_phpplmul_summul_n223,
         SBOX_Inst_f1_phpplmul_summul_n222, SBOX_Inst_f1_phpplmul_summul_n221,
         SBOX_Inst_f1_phpplmul_summul_n220, SBOX_Inst_f1_phpplmul_summul_n219,
         SBOX_Inst_f1_phpplmul_summul_n218, SBOX_Inst_f1_phpplmul_summul_n217,
         SBOX_Inst_f1_phpplmul_summul_n216, SBOX_Inst_f1_phpplmul_summul_n215,
         SBOX_Inst_f1_phpplmul_AddNewMaskp_n6,
         SBOX_Inst_f1_phpplmul_AddNewMaskp_n5,
         SBOX_Inst_f1_phpplmul_lowmul_n302, SBOX_Inst_f1_phpplmul_lowmul_n301,
         SBOX_Inst_f1_phpplmul_lowmul_n300, SBOX_Inst_f1_phpplmul_lowmul_n299,
         SBOX_Inst_f1_phpplmul_lowmul_n298, SBOX_Inst_f1_phpplmul_lowmul_n297,
         SBOX_Inst_f1_phpplmul_lowmul_n296, SBOX_Inst_f1_phpplmul_lowmul_n295,
         SBOX_Inst_f1_phpplmul_lowmul_n294, SBOX_Inst_f1_phpplmul_lowmul_n293,
         SBOX_Inst_f1_phpplmul_lowmul_n292, SBOX_Inst_f1_phpplmul_lowmul_n291,
         SBOX_Inst_f1_phpplmul_lowmul_n290, SBOX_Inst_f1_phpplmul_lowmul_n289,
         SBOX_Inst_f1_phpplmul_lowmul_n288, SBOX_Inst_f1_phpplmul_lowmul_n287,
         SBOX_Inst_f1_phpplmul_lowmul_n286, SBOX_Inst_f1_phpplmul_lowmul_n285,
         SBOX_Inst_f1_phpplmul_lowmul_n284, SBOX_Inst_f1_phpplmul_lowmul_n283,
         SBOX_Inst_f1_phpplmul_lowmul_n282, SBOX_Inst_f1_phpplmul_lowmul_n281,
         SBOX_Inst_f1_phpplmul_lowmul_n280, SBOX_Inst_f1_phpplmul_lowmul_n279,
         SBOX_Inst_f1_phpplmul_lowmul_n278, SBOX_Inst_f1_phpplmul_lowmul_n277,
         SBOX_Inst_f1_phpplmul_lowmul_n276, SBOX_Inst_f1_phpplmul_lowmul_n275,
         SBOX_Inst_f1_phpplmul_lowmul_n274, SBOX_Inst_f1_phpplmul_lowmul_n273,
         SBOX_Inst_f1_phpplmul_lowmul_n272, SBOX_Inst_f1_phpplmul_lowmul_n271,
         SBOX_Inst_f1_phpplmul_lowmul_n270, SBOX_Inst_f1_phpplmul_lowmul_n269,
         SBOX_Inst_f1_phpplmul_lowmul_n268, SBOX_Inst_f1_phpplmul_lowmul_n267,
         SBOX_Inst_f1_phpplmul_lowmul_n266, SBOX_Inst_f1_phpplmul_lowmul_n265,
         SBOX_Inst_f1_phpplmul_lowmul_n264, SBOX_Inst_f1_phpplmul_lowmul_n263,
         SBOX_Inst_f1_phpplmul_lowmul_n262, SBOX_Inst_f1_phpplmul_lowmul_n261,
         SBOX_Inst_f1_phpplmul_lowmul_n260, SBOX_Inst_f1_phpplmul_lowmul_n259,
         SBOX_Inst_f1_phpplmul_lowmul_n258, SBOX_Inst_f1_phpplmul_lowmul_n257,
         SBOX_Inst_f1_phpplmul_lowmul_n256, SBOX_Inst_f1_phpplmul_lowmul_n255,
         SBOX_Inst_f1_phpplmul_lowmul_n254, SBOX_Inst_f1_phpplmul_lowmul_n253,
         SBOX_Inst_f1_phpplmul_lowmul_n252, SBOX_Inst_f1_phpplmul_lowmul_n251,
         SBOX_Inst_f1_phpplmul_lowmul_n250, SBOX_Inst_f1_phpplmul_lowmul_n249,
         SBOX_Inst_f1_phpplmul_lowmul_n248, SBOX_Inst_f1_phpplmul_lowmul_n247,
         SBOX_Inst_f1_phpplmul_lowmul_n246, SBOX_Inst_f1_phpplmul_lowmul_n245,
         SBOX_Inst_f1_phpplmul_lowmul_n244, SBOX_Inst_f1_phpplmul_lowmul_n243,
         SBOX_Inst_f1_phpplmul_lowmul_n242, SBOX_Inst_f1_phpplmul_lowmul_n241,
         SBOX_Inst_f1_phpplmul_lowmul_n240, SBOX_Inst_f1_phpplmul_lowmul_n239,
         SBOX_Inst_f1_phpplmul_lowmul_n238, SBOX_Inst_f1_phpplmul_lowmul_n237,
         SBOX_Inst_f1_phpplmul_lowmul_n236, SBOX_Inst_f1_phpplmul_lowmul_n235,
         SBOX_Inst_f1_phpplmul_lowmul_n234, SBOX_Inst_f1_phpplmul_lowmul_n233,
         SBOX_Inst_f1_phpplmul_lowmul_n232, SBOX_Inst_f1_phpplmul_lowmul_n231,
         SBOX_Inst_f1_phpplmul_lowmul_n230, SBOX_Inst_f1_phpplmul_lowmul_n229,
         SBOX_Inst_f1_phpplmul_lowmul_n228, SBOX_Inst_f1_phpplmul_lowmul_n227,
         SBOX_Inst_f1_phpplmul_lowmul_n226, SBOX_Inst_f1_phpplmul_lowmul_n225,
         SBOX_Inst_f1_phpplmul_lowmul_n224, SBOX_Inst_f1_phpplmul_lowmul_n223,
         SBOX_Inst_f1_phpplmul_lowmul_n222, SBOX_Inst_f1_phpplmul_lowmul_n221,
         SBOX_Inst_f1_phpplmul_lowmul_n220, SBOX_Inst_f1_phpplmul_lowmul_n219,
         SBOX_Inst_f1_phpplmul_lowmul_n218, SBOX_Inst_f1_phpplmul_lowmul_n217,
         SBOX_Inst_f1_phpplmul_lowmul_n216,
         SBOX_Inst_f1_phpplmul_AddNewMaskpl_n6,
         SBOX_Inst_f1_phpplmul_AddNewMaskpl_n5, SBOX_PL_1_n54, SBOX_PL_1_n53,
         SBOX_PL_1_n52, SBOX_PL_1_n51, SBOX_PL_1_n50, SBOX_PL_1_n49,
         SBOX_PL_1_n48, SBOX_PL_1_n47, SBOX_PL_1_n46, SBOX_PL_1_n45,
         SBOX_PL_1_n44, SBOX_PL_1_n43, SBOX_PL_1_n42, SBOX_PL_1_n41,
         SBOX_PL_1_n40, SBOX_PL_1_n39, SBOX_PL_1_n38, SBOX_PL_1_n37,
         SBOX_PL_1_n36, SBOX_PL_1_n35, SBOX_PL_1_n34, SBOX_PL_1_n33,
         SBOX_PL_1_n32, SBOX_PL_1_n31, SBOX_PL_1_n30, SBOX_PL_1_n29,
         SBOX_PL_1_n28, SBOX_PL_1_n27, SBOX_PL_1_n26, SBOX_PL_1_n25,
         SBOX_PL_1_n24, SBOX_PL_1_n23, SBOX_PL_1_n22, SBOX_PL_1_n21,
         SBOX_PL_1_n20, SBOX_PL_1_n19, SBOX_PL_1_n18, SBOX_PL_1_n17,
         SBOX_PL_1_n16, SBOX_PL_1_n15, SBOX_PL_1_n14, SBOX_PL_1_n13,
         SBOX_PL_1_n12, SBOX_PL_1_n11, SBOX_PL_1_n10, SBOX_PL_1_n9,
         SBOX_PL_1_n8, SBOX_PL_1_n7, SBOX_PL_1_n6, SBOX_PL_1_n5, SBOX_PL_1_n4,
         SBOX_PL_1_n3, SBOX_PL_1_n2, SBOX_PL_1_n1, SBOX_PL_1_n162,
         SBOX_PL_1_n161, SBOX_PL_1_n160, SBOX_PL_1_n159, SBOX_PL_1_n158,
         SBOX_PL_1_n157, SBOX_PL_1_n156, SBOX_PL_1_n155, SBOX_PL_1_n154,
         SBOX_PL_1_n153, SBOX_PL_1_n152, SBOX_PL_1_n151, SBOX_PL_1_n150,
         SBOX_PL_1_n149, SBOX_PL_1_n148, SBOX_PL_1_n147, SBOX_PL_1_n146,
         SBOX_PL_1_n145, SBOX_PL_1_n144, SBOX_PL_1_n143, SBOX_PL_1_n142,
         SBOX_PL_1_n141, SBOX_PL_1_n140, SBOX_PL_1_n139, SBOX_PL_1_n138,
         SBOX_PL_1_n137, SBOX_PL_1_n136, SBOX_PL_1_n135, SBOX_PL_1_n134,
         SBOX_PL_1_n133, SBOX_PL_1_n132, SBOX_PL_1_n131, SBOX_PL_1_n130,
         SBOX_PL_1_n129, SBOX_PL_1_n128, SBOX_PL_1_n127, SBOX_PL_1_n126,
         SBOX_PL_1_n125, SBOX_PL_1_n124, SBOX_PL_1_n123, SBOX_PL_1_n122,
         SBOX_PL_1_n121, SBOX_PL_1_n120, SBOX_PL_1_n119, SBOX_PL_1_n118,
         SBOX_PL_1_n117, SBOX_PL_1_n116, SBOX_PL_1_n115, SBOX_PL_1_n114,
         SBOX_PL_1_n113, SBOX_PL_1_n112, SBOX_PL_1_n111, SBOX_PL_1_n110,
         SBOX_PL_1_n109, SBOX_PL_1_n108, SBOX_PL_1_n107, SBOX_PL_1_n106,
         SBOX_PL_1_n105, SBOX_PL_1_n104, SBOX_PL_1_n103, SBOX_PL_1_n102,
         SBOX_PL_1_n101, SBOX_PL_1_n100, SBOX_PL_1_n99, SBOX_PL_1_n98,
         SBOX_PL_1_n97, SBOX_PL_1_n96, SBOX_PL_1_n95, SBOX_PL_1_n94,
         SBOX_PL_1_n93, SBOX_PL_1_n92, SBOX_PL_1_n91, SBOX_PL_1_n90,
         SBOX_PL_1_n89, SBOX_PL_1_n88, SBOX_PL_1_n87, SBOX_PL_1_n86,
         SBOX_PL_1_n85, SBOX_PL_1_n84, SBOX_PL_1_n83, SBOX_PL_1_n82,
         SBOX_PL_1_n81, SBOX_PL_1_n80, SBOX_PL_1_n79, SBOX_PL_1_n78,
         SBOX_PL_1_n77, SBOX_PL_1_n76, SBOX_PL_1_n75, SBOX_PL_1_n74,
         SBOX_PL_1_n73, SBOX_PL_1_n72, SBOX_PL_1_n71, SBOX_PL_1_n70,
         SBOX_PL_1_n69, SBOX_PL_1_n68, SBOX_PL_1_n67, SBOX_PL_1_n66,
         SBOX_PL_1_n65, SBOX_PL_1_n64, SBOX_PL_1_n63, SBOX_PL_1_n62,
         SBOX_PL_1_n61, SBOX_PL_1_n60, SBOX_PL_1_n59, SBOX_PL_1_n58,
         SBOX_PL_1_n57, SBOX_PL_1_n56, SBOX_PL_1_n55,
         SBOX_Inst_f2_abmul_pw2_0_, SBOX_Inst_f2_abmul_pw2_1_,
         SBOX_Inst_f2_abmul_pw2_2_, SBOX_Inst_f2_abmul_pw2_3_,
         SBOX_Inst_f2_abmul_pw2_4_, SBOX_Inst_f2_abmul_pw2_5_,
         SBOX_Inst_f2_dinv_1_mul_n303, SBOX_Inst_f2_dinv_1_mul_n302,
         SBOX_Inst_f2_dinv_1_mul_n301, SBOX_Inst_f2_dinv_1_mul_n300,
         SBOX_Inst_f2_dinv_1_mul_n299, SBOX_Inst_f2_dinv_1_mul_n298,
         SBOX_Inst_f2_dinv_1_mul_n297, SBOX_Inst_f2_dinv_1_mul_n296,
         SBOX_Inst_f2_dinv_1_mul_n295, SBOX_Inst_f2_dinv_1_mul_n294,
         SBOX_Inst_f2_dinv_1_mul_n293, SBOX_Inst_f2_dinv_1_mul_n292,
         SBOX_Inst_f2_dinv_1_mul_n291, SBOX_Inst_f2_dinv_1_mul_n290,
         SBOX_Inst_f2_dinv_1_mul_n289, SBOX_Inst_f2_dinv_1_mul_n288,
         SBOX_Inst_f2_dinv_1_mul_n287, SBOX_Inst_f2_dinv_1_mul_n286,
         SBOX_Inst_f2_dinv_1_mul_n285, SBOX_Inst_f2_dinv_1_mul_n284,
         SBOX_Inst_f2_dinv_1_mul_n283, SBOX_Inst_f2_dinv_1_mul_n282,
         SBOX_Inst_f2_dinv_1_mul_n281, SBOX_Inst_f2_dinv_1_mul_n280,
         SBOX_Inst_f2_dinv_1_mul_n279, SBOX_Inst_f2_dinv_1_mul_n278,
         SBOX_Inst_f2_dinv_1_mul_n277, SBOX_Inst_f2_dinv_1_mul_n276,
         SBOX_Inst_f2_dinv_1_mul_n275, SBOX_Inst_f2_dinv_1_mul_n274,
         SBOX_Inst_f2_dinv_1_mul_n273, SBOX_Inst_f2_dinv_1_mul_n272,
         SBOX_Inst_f2_dinv_1_mul_n271, SBOX_Inst_f2_dinv_1_mul_n270,
         SBOX_Inst_f2_dinv_1_mul_n269, SBOX_Inst_f2_dinv_1_mul_n268,
         SBOX_Inst_f2_dinv_1_mul_n267, SBOX_Inst_f2_dinv_1_mul_n266,
         SBOX_Inst_f2_dinv_1_mul_n265, SBOX_Inst_f2_dinv_1_mul_n264,
         SBOX_Inst_f2_dinv_1_mul_n263, SBOX_Inst_f2_dinv_1_mul_n262,
         SBOX_Inst_f2_dinv_1_mul_n261, SBOX_Inst_f2_dinv_1_mul_n260,
         SBOX_Inst_f2_dinv_1_mul_n259, SBOX_Inst_f2_dinv_1_mul_n258,
         SBOX_Inst_f2_dinv_1_mul_n257, SBOX_Inst_f2_dinv_1_mul_n256,
         SBOX_Inst_f2_dinv_1_mul_n255, SBOX_Inst_f2_dinv_1_mul_n254,
         SBOX_Inst_f2_dinv_1_mul_n253, SBOX_Inst_f2_dinv_1_mul_n252,
         SBOX_Inst_f2_dinv_1_mul_n251, SBOX_Inst_f2_dinv_1_mul_n250,
         SBOX_Inst_f2_dinv_1_mul_n249, SBOX_Inst_f2_dinv_1_mul_n248,
         SBOX_Inst_f2_dinv_1_mul_n247, SBOX_Inst_f2_dinv_1_mul_n246,
         SBOX_Inst_f2_dinv_1_mul_n245, SBOX_Inst_f2_dinv_1_mul_n244,
         SBOX_Inst_f2_dinv_1_mul_n243, SBOX_Inst_f2_dinv_1_mul_n242,
         SBOX_Inst_f2_dinv_1_mul_n241, SBOX_Inst_f2_dinv_1_mul_n240,
         SBOX_Inst_f2_dinv_1_mul_n239, SBOX_Inst_f2_dinv_1_mul_n238,
         SBOX_Inst_f2_dinv_1_mul_n237, SBOX_Inst_f2_dinv_1_mul_n236,
         SBOX_Inst_f2_dinv_1_mul_n235, SBOX_Inst_f2_dinv_1_mul_n234,
         SBOX_Inst_f2_dinv_1_mul_n233, SBOX_Inst_f2_dinv_1_mul_n232,
         SBOX_Inst_f2_dinv_1_mul_n231, SBOX_Inst_f2_dinv_1_mul_n230,
         SBOX_Inst_f2_dinv_1_mul_n229, SBOX_Inst_f2_dinv_1_mul_n228,
         SBOX_Inst_f2_dinv_1_mul_n227, SBOX_Inst_f2_dinv_1_mul_n226,
         SBOX_Inst_f2_dinv_1_mul_n225, SBOX_Inst_f2_dinv_1_mul_n224,
         SBOX_Inst_f2_dinv_1_mul_n223, SBOX_Inst_f2_dinv_1_mul_n222,
         SBOX_Inst_f2_dinv_1_mul_n221, SBOX_Inst_f2_dinv_1_mul_n220,
         SBOX_Inst_f2_dinv_1_mul_n219, SBOX_Inst_f2_dinv_1_mul_n218,
         SBOX_Inst_f2_dinv_1_mul_n217, SBOX_Inst_f2_dinv_1_mul_n216,
         SBOX_Inst_f2_dinv_1_mul_n215, SBOX_Inst_f2_dinv_1_AddNewMaskab_n6,
         SBOX_Inst_f2_dinv_1_AddNewMaskab_n5,
         SBOX_Inst_f2_dinv_1_AddNewMasksA2N_n6,
         SBOX_Inst_f2_dinv_1_AddNewMasksA2N_n5, SBOX_PL_2_n48, SBOX_PL_2_n47,
         SBOX_PL_2_n46, SBOX_PL_2_n45, SBOX_PL_2_n44, SBOX_PL_2_n43,
         SBOX_PL_2_n42, SBOX_PL_2_n41, SBOX_PL_2_n40, SBOX_PL_2_n39,
         SBOX_PL_2_n38, SBOX_PL_2_n37, SBOX_PL_2_n36, SBOX_PL_2_n35,
         SBOX_PL_2_n34, SBOX_PL_2_n33, SBOX_PL_2_n32, SBOX_PL_2_n31,
         SBOX_PL_2_n30, SBOX_PL_2_n29, SBOX_PL_2_n28, SBOX_PL_2_n27,
         SBOX_PL_2_n26, SBOX_PL_2_n25, SBOX_PL_2_n24, SBOX_PL_2_n23,
         SBOX_PL_2_n22, SBOX_PL_2_n21, SBOX_PL_2_n20, SBOX_PL_2_n19,
         SBOX_PL_2_n18, SBOX_PL_2_n17, SBOX_PL_2_n16, SBOX_PL_2_n15,
         SBOX_PL_2_n14, SBOX_PL_2_n13, SBOX_PL_2_n12, SBOX_PL_2_n11,
         SBOX_PL_2_n10, SBOX_PL_2_n9, SBOX_PL_2_n8, SBOX_PL_2_n7, SBOX_PL_2_n6,
         SBOX_PL_2_n5, SBOX_PL_2_n4, SBOX_PL_2_n3, SBOX_PL_2_n2, SBOX_PL_2_n1,
         SBOX_PL_2_n144, SBOX_PL_2_n143, SBOX_PL_2_n142, SBOX_PL_2_n141,
         SBOX_PL_2_n140, SBOX_PL_2_n139, SBOX_PL_2_n138, SBOX_PL_2_n137,
         SBOX_PL_2_n136, SBOX_PL_2_n135, SBOX_PL_2_n134, SBOX_PL_2_n133,
         SBOX_PL_2_n132, SBOX_PL_2_n131, SBOX_PL_2_n130, SBOX_PL_2_n129,
         SBOX_PL_2_n128, SBOX_PL_2_n127, SBOX_PL_2_n126, SBOX_PL_2_n125,
         SBOX_PL_2_n124, SBOX_PL_2_n123, SBOX_PL_2_n122, SBOX_PL_2_n121,
         SBOX_PL_2_n120, SBOX_PL_2_n119, SBOX_PL_2_n118, SBOX_PL_2_n117,
         SBOX_PL_2_n116, SBOX_PL_2_n115, SBOX_PL_2_n114, SBOX_PL_2_n113,
         SBOX_PL_2_n112, SBOX_PL_2_n111, SBOX_PL_2_n110, SBOX_PL_2_n109,
         SBOX_PL_2_n108, SBOX_PL_2_n107, SBOX_PL_2_n106, SBOX_PL_2_n105,
         SBOX_PL_2_n104, SBOX_PL_2_n103, SBOX_PL_2_n102, SBOX_PL_2_n101,
         SBOX_PL_2_n100, SBOX_PL_2_n99, SBOX_PL_2_n98, SBOX_PL_2_n97,
         SBOX_PL_2_n96, SBOX_PL_2_n95, SBOX_PL_2_n94, SBOX_PL_2_n93,
         SBOX_PL_2_n92, SBOX_PL_2_n91, SBOX_PL_2_n90, SBOX_PL_2_n89,
         SBOX_PL_2_n88, SBOX_PL_2_n87, SBOX_PL_2_n86, SBOX_PL_2_n85,
         SBOX_PL_2_n84, SBOX_PL_2_n83, SBOX_PL_2_n82, SBOX_PL_2_n81,
         SBOX_PL_2_n80, SBOX_PL_2_n79, SBOX_PL_2_n78, SBOX_PL_2_n77,
         SBOX_PL_2_n76, SBOX_PL_2_n75, SBOX_PL_2_n74, SBOX_PL_2_n73,
         SBOX_PL_2_n72, SBOX_PL_2_n71, SBOX_PL_2_n70, SBOX_PL_2_n69,
         SBOX_PL_2_n68, SBOX_PL_2_n67, SBOX_PL_2_n66, SBOX_PL_2_n65,
         SBOX_PL_2_n64, SBOX_PL_2_n63, SBOX_PL_2_n62, SBOX_PL_2_n61,
         SBOX_PL_2_n60, SBOX_PL_2_n59, SBOX_PL_2_n58, SBOX_PL_2_n57,
         SBOX_PL_2_n56, SBOX_PL_2_n55, SBOX_PL_2_n54, SBOX_PL_2_n53,
         SBOX_PL_2_n52, SBOX_PL_2_n51, SBOX_PL_2_n50, SBOX_PL_2_n49,
         SBOX_Inst_f3_dinv_2_d_0_, SBOX_Inst_f3_dinv_2_d_1_,
         SBOX_Inst_f3_dinv_2_d_2_, SBOX_Inst_f3_dinv_2_d_3_,
         SBOX_Inst_f3_dinv_2_d_4_, SBOX_Inst_f3_dinv_2_d_5_,
         SBOX_Inst_f3_dinv_2_himul_n308, SBOX_Inst_f3_dinv_2_himul_n307,
         SBOX_Inst_f3_dinv_2_himul_n306, SBOX_Inst_f3_dinv_2_himul_n305,
         SBOX_Inst_f3_dinv_2_himul_n304, SBOX_Inst_f3_dinv_2_himul_n303,
         SBOX_Inst_f3_dinv_2_himul_n302, SBOX_Inst_f3_dinv_2_himul_n301,
         SBOX_Inst_f3_dinv_2_himul_n300, SBOX_Inst_f3_dinv_2_himul_n299,
         SBOX_Inst_f3_dinv_2_himul_n298, SBOX_Inst_f3_dinv_2_himul_n297,
         SBOX_Inst_f3_dinv_2_himul_n296, SBOX_Inst_f3_dinv_2_himul_n295,
         SBOX_Inst_f3_dinv_2_himul_n294, SBOX_Inst_f3_dinv_2_himul_n293,
         SBOX_Inst_f3_dinv_2_himul_n292, SBOX_Inst_f3_dinv_2_himul_n291,
         SBOX_Inst_f3_dinv_2_himul_n290, SBOX_Inst_f3_dinv_2_himul_n289,
         SBOX_Inst_f3_dinv_2_himul_n288, SBOX_Inst_f3_dinv_2_himul_n287,
         SBOX_Inst_f3_dinv_2_himul_n286, SBOX_Inst_f3_dinv_2_himul_n285,
         SBOX_Inst_f3_dinv_2_himul_n284, SBOX_Inst_f3_dinv_2_himul_n283,
         SBOX_Inst_f3_dinv_2_himul_n282, SBOX_Inst_f3_dinv_2_himul_n281,
         SBOX_Inst_f3_dinv_2_himul_n280, SBOX_Inst_f3_dinv_2_himul_n279,
         SBOX_Inst_f3_dinv_2_himul_n278, SBOX_Inst_f3_dinv_2_himul_n277,
         SBOX_Inst_f3_dinv_2_himul_n276, SBOX_Inst_f3_dinv_2_himul_n275,
         SBOX_Inst_f3_dinv_2_himul_n274, SBOX_Inst_f3_dinv_2_himul_n273,
         SBOX_Inst_f3_dinv_2_himul_n272, SBOX_Inst_f3_dinv_2_himul_n271,
         SBOX_Inst_f3_dinv_2_himul_n270, SBOX_Inst_f3_dinv_2_himul_n269,
         SBOX_Inst_f3_dinv_2_himul_n268, SBOX_Inst_f3_dinv_2_himul_n267,
         SBOX_Inst_f3_dinv_2_himul_n266, SBOX_Inst_f3_dinv_2_himul_n265,
         SBOX_Inst_f3_dinv_2_himul_n264, SBOX_Inst_f3_dinv_2_himul_n263,
         SBOX_Inst_f3_dinv_2_himul_n262, SBOX_Inst_f3_dinv_2_himul_n261,
         SBOX_Inst_f3_dinv_2_himul_n260, SBOX_Inst_f3_dinv_2_himul_n259,
         SBOX_Inst_f3_dinv_2_himul_n258, SBOX_Inst_f3_dinv_2_himul_n257,
         SBOX_Inst_f3_dinv_2_himul_n256, SBOX_Inst_f3_dinv_2_himul_n255,
         SBOX_Inst_f3_dinv_2_himul_n254, SBOX_Inst_f3_dinv_2_himul_n253,
         SBOX_Inst_f3_dinv_2_himul_n252, SBOX_Inst_f3_dinv_2_himul_n251,
         SBOX_Inst_f3_dinv_2_himul_n250, SBOX_Inst_f3_dinv_2_himul_n249,
         SBOX_Inst_f3_dinv_2_himul_n248, SBOX_Inst_f3_dinv_2_himul_n247,
         SBOX_Inst_f3_dinv_2_himul_n246, SBOX_Inst_f3_dinv_2_himul_n245,
         SBOX_Inst_f3_dinv_2_himul_n244, SBOX_Inst_f3_dinv_2_himul_n243,
         SBOX_Inst_f3_dinv_2_himul_n242, SBOX_Inst_f3_dinv_2_himul_n241,
         SBOX_Inst_f3_dinv_2_himul_n240, SBOX_Inst_f3_dinv_2_himul_n239,
         SBOX_Inst_f3_dinv_2_himul_n238, SBOX_Inst_f3_dinv_2_himul_n237,
         SBOX_Inst_f3_dinv_2_himul_n236, SBOX_Inst_f3_dinv_2_himul_n235,
         SBOX_Inst_f3_dinv_2_himul_n234, SBOX_Inst_f3_dinv_2_himul_n233,
         SBOX_Inst_f3_dinv_2_himul_n232, SBOX_Inst_f3_dinv_2_himul_n231,
         SBOX_Inst_f3_dinv_2_himul_n230, SBOX_Inst_f3_dinv_2_himul_n229,
         SBOX_Inst_f3_dinv_2_himul_n228, SBOX_Inst_f3_dinv_2_himul_n227,
         SBOX_Inst_f3_dinv_2_himul_n226, SBOX_Inst_f3_dinv_2_himul_n225,
         SBOX_Inst_f3_dinv_2_himul_n224, SBOX_Inst_f3_dinv_2_himul_n223,
         SBOX_Inst_f3_dinv_2_himul_n222, SBOX_Inst_f3_dinv_2_himul_n221,
         SBOX_Inst_f3_dinv_2_himul_n220, SBOX_Inst_f3_dinv_2_himul_n219,
         SBOX_Inst_f3_dinv_2_himul_n218, SBOX_Inst_f3_dinv_2_himul_n217,
         SBOX_Inst_f3_dinv_2_himul_n216, SBOX_Inst_f3_dinv_2_himul_n215,
         SBOX_Inst_f3_dinv_2_lowmul_n308, SBOX_Inst_f3_dinv_2_lowmul_n307,
         SBOX_Inst_f3_dinv_2_lowmul_n306, SBOX_Inst_f3_dinv_2_lowmul_n305,
         SBOX_Inst_f3_dinv_2_lowmul_n304, SBOX_Inst_f3_dinv_2_lowmul_n303,
         SBOX_Inst_f3_dinv_2_lowmul_n302, SBOX_Inst_f3_dinv_2_lowmul_n301,
         SBOX_Inst_f3_dinv_2_lowmul_n300, SBOX_Inst_f3_dinv_2_lowmul_n299,
         SBOX_Inst_f3_dinv_2_lowmul_n298, SBOX_Inst_f3_dinv_2_lowmul_n297,
         SBOX_Inst_f3_dinv_2_lowmul_n296, SBOX_Inst_f3_dinv_2_lowmul_n295,
         SBOX_Inst_f3_dinv_2_lowmul_n294, SBOX_Inst_f3_dinv_2_lowmul_n293,
         SBOX_Inst_f3_dinv_2_lowmul_n292, SBOX_Inst_f3_dinv_2_lowmul_n291,
         SBOX_Inst_f3_dinv_2_lowmul_n290, SBOX_Inst_f3_dinv_2_lowmul_n289,
         SBOX_Inst_f3_dinv_2_lowmul_n288, SBOX_Inst_f3_dinv_2_lowmul_n287,
         SBOX_Inst_f3_dinv_2_lowmul_n286, SBOX_Inst_f3_dinv_2_lowmul_n285,
         SBOX_Inst_f3_dinv_2_lowmul_n284, SBOX_Inst_f3_dinv_2_lowmul_n283,
         SBOX_Inst_f3_dinv_2_lowmul_n282, SBOX_Inst_f3_dinv_2_lowmul_n281,
         SBOX_Inst_f3_dinv_2_lowmul_n280, SBOX_Inst_f3_dinv_2_lowmul_n279,
         SBOX_Inst_f3_dinv_2_lowmul_n278, SBOX_Inst_f3_dinv_2_lowmul_n277,
         SBOX_Inst_f3_dinv_2_lowmul_n276, SBOX_Inst_f3_dinv_2_lowmul_n275,
         SBOX_Inst_f3_dinv_2_lowmul_n274, SBOX_Inst_f3_dinv_2_lowmul_n273,
         SBOX_Inst_f3_dinv_2_lowmul_n272, SBOX_Inst_f3_dinv_2_lowmul_n271,
         SBOX_Inst_f3_dinv_2_lowmul_n270, SBOX_Inst_f3_dinv_2_lowmul_n269,
         SBOX_Inst_f3_dinv_2_lowmul_n268, SBOX_Inst_f3_dinv_2_lowmul_n267,
         SBOX_Inst_f3_dinv_2_lowmul_n266, SBOX_Inst_f3_dinv_2_lowmul_n265,
         SBOX_Inst_f3_dinv_2_lowmul_n264, SBOX_Inst_f3_dinv_2_lowmul_n263,
         SBOX_Inst_f3_dinv_2_lowmul_n262, SBOX_Inst_f3_dinv_2_lowmul_n261,
         SBOX_Inst_f3_dinv_2_lowmul_n260, SBOX_Inst_f3_dinv_2_lowmul_n259,
         SBOX_Inst_f3_dinv_2_lowmul_n258, SBOX_Inst_f3_dinv_2_lowmul_n257,
         SBOX_Inst_f3_dinv_2_lowmul_n256, SBOX_Inst_f3_dinv_2_lowmul_n255,
         SBOX_Inst_f3_dinv_2_lowmul_n254, SBOX_Inst_f3_dinv_2_lowmul_n253,
         SBOX_Inst_f3_dinv_2_lowmul_n252, SBOX_Inst_f3_dinv_2_lowmul_n251,
         SBOX_Inst_f3_dinv_2_lowmul_n250, SBOX_Inst_f3_dinv_2_lowmul_n249,
         SBOX_Inst_f3_dinv_2_lowmul_n248, SBOX_Inst_f3_dinv_2_lowmul_n247,
         SBOX_Inst_f3_dinv_2_lowmul_n246, SBOX_Inst_f3_dinv_2_lowmul_n245,
         SBOX_Inst_f3_dinv_2_lowmul_n244, SBOX_Inst_f3_dinv_2_lowmul_n243,
         SBOX_Inst_f3_dinv_2_lowmul_n242, SBOX_Inst_f3_dinv_2_lowmul_n241,
         SBOX_Inst_f3_dinv_2_lowmul_n240, SBOX_Inst_f3_dinv_2_lowmul_n239,
         SBOX_Inst_f3_dinv_2_lowmul_n238, SBOX_Inst_f3_dinv_2_lowmul_n237,
         SBOX_Inst_f3_dinv_2_lowmul_n236, SBOX_Inst_f3_dinv_2_lowmul_n235,
         SBOX_Inst_f3_dinv_2_lowmul_n234, SBOX_Inst_f3_dinv_2_lowmul_n233,
         SBOX_Inst_f3_dinv_2_lowmul_n232, SBOX_Inst_f3_dinv_2_lowmul_n231,
         SBOX_Inst_f3_dinv_2_lowmul_n230, SBOX_Inst_f3_dinv_2_lowmul_n229,
         SBOX_Inst_f3_dinv_2_lowmul_n228, SBOX_Inst_f3_dinv_2_lowmul_n227,
         SBOX_Inst_f3_dinv_2_lowmul_n226, SBOX_Inst_f3_dinv_2_lowmul_n225,
         SBOX_Inst_f3_dinv_2_lowmul_n224, SBOX_Inst_f3_dinv_2_lowmul_n223,
         SBOX_Inst_f3_dinv_2_lowmul_n222, SBOX_Inst_f3_dinv_2_lowmul_n221,
         SBOX_Inst_f3_dinv_2_lowmul_n220, SBOX_Inst_f3_dinv_2_lowmul_n219,
         SBOX_Inst_f3_dinv_2_lowmul_n218, SBOX_Inst_f3_dinv_2_lowmul_n217,
         SBOX_Inst_f3_dinv_2_lowmul_n216, SBOX_Inst_f3_dinv_2_lowmul_n215,
         SBOX_Inst_f3_dinv_2_AddNewMaskQ_n4,
         SBOX_Inst_f3_dinv_2_AddNewMaskQ_n3,
         SBOX_Inst_f3_dinv_2_AddNewMaskQ_n2,
         SBOX_Inst_f3_dinv_2_AddNewMaskQ_n1, SBOX_PL_3_n252, SBOX_PL_3_n251,
         SBOX_PL_3_n250, SBOX_PL_3_n249, SBOX_PL_3_n248, SBOX_PL_3_n247,
         SBOX_PL_3_n246, SBOX_PL_3_n245, SBOX_PL_3_n244, SBOX_PL_3_n243,
         SBOX_PL_3_n242, SBOX_PL_3_n241, SBOX_PL_3_n240, SBOX_PL_3_n239,
         SBOX_PL_3_n238, SBOX_PL_3_n237, SBOX_PL_3_n236, SBOX_PL_3_n235,
         SBOX_PL_3_n234, SBOX_PL_3_n233, SBOX_PL_3_n232, SBOX_PL_3_n231,
         SBOX_PL_3_n230, SBOX_PL_3_n229, SBOX_PL_3_n228, SBOX_PL_3_n227,
         SBOX_PL_3_n226, SBOX_PL_3_n225, SBOX_PL_3_n224, SBOX_PL_3_n223,
         SBOX_PL_3_n222, SBOX_PL_3_n221, SBOX_PL_3_n220, SBOX_PL_3_n219,
         SBOX_PL_3_n218, SBOX_PL_3_n217, SBOX_PL_3_n180, SBOX_PL_3_n179,
         SBOX_PL_3_n178, SBOX_PL_3_n177, SBOX_PL_3_n176, SBOX_PL_3_n175,
         SBOX_PL_3_n174, SBOX_PL_3_n173, SBOX_PL_3_n172, SBOX_PL_3_n171,
         SBOX_PL_3_n170, SBOX_PL_3_n169, SBOX_PL_3_n168, SBOX_PL_3_n167,
         SBOX_PL_3_n166, SBOX_PL_3_n165, SBOX_PL_3_n164, SBOX_PL_3_n163,
         SBOX_PL_3_n162, SBOX_PL_3_n161, SBOX_PL_3_n160, SBOX_PL_3_n159,
         SBOX_PL_3_n158, SBOX_PL_3_n157, SBOX_PL_3_n156, SBOX_PL_3_n155,
         SBOX_PL_3_n154, SBOX_PL_3_n153, SBOX_PL_3_n152, SBOX_PL_3_n151,
         SBOX_PL_3_n150, SBOX_PL_3_n149, SBOX_PL_3_n148, SBOX_PL_3_n147,
         SBOX_PL_3_n146, SBOX_PL_3_n145, SBOX_PL_3_n144, SBOX_PL_3_n143,
         SBOX_PL_3_n142, SBOX_PL_3_n141, SBOX_PL_3_n140, SBOX_PL_3_n139,
         SBOX_PL_3_n138, SBOX_PL_3_n137, SBOX_PL_3_n136, SBOX_PL_3_n135,
         SBOX_PL_3_n134, SBOX_PL_3_n133, SBOX_PL_3_n132, SBOX_PL_3_n131,
         SBOX_PL_3_n130, SBOX_PL_3_n129, SBOX_PL_3_n128, SBOX_PL_3_n127,
         SBOX_PL_3_n126, SBOX_PL_3_n125, SBOX_PL_3_n124, SBOX_PL_3_n123,
         SBOX_PL_3_n122, SBOX_PL_3_n121, SBOX_PL_3_n120, SBOX_PL_3_n119,
         SBOX_PL_3_n118, SBOX_PL_3_n117, SBOX_PL_3_n116, SBOX_PL_3_n115,
         SBOX_PL_3_n114, SBOX_PL_3_n113, SBOX_PL_3_n112, SBOX_PL_3_n111,
         SBOX_PL_3_n110, SBOX_PL_3_n109, SBOX_Inst_f4_multd_L_himul_n302,
         SBOX_Inst_f4_multd_L_himul_n301, SBOX_Inst_f4_multd_L_himul_n300,
         SBOX_Inst_f4_multd_L_himul_n299, SBOX_Inst_f4_multd_L_himul_n298,
         SBOX_Inst_f4_multd_L_himul_n297, SBOX_Inst_f4_multd_L_himul_n296,
         SBOX_Inst_f4_multd_L_himul_n295, SBOX_Inst_f4_multd_L_himul_n294,
         SBOX_Inst_f4_multd_L_himul_n293, SBOX_Inst_f4_multd_L_himul_n292,
         SBOX_Inst_f4_multd_L_himul_n291, SBOX_Inst_f4_multd_L_himul_n290,
         SBOX_Inst_f4_multd_L_himul_n289, SBOX_Inst_f4_multd_L_himul_n288,
         SBOX_Inst_f4_multd_L_himul_n287, SBOX_Inst_f4_multd_L_himul_n286,
         SBOX_Inst_f4_multd_L_himul_n285, SBOX_Inst_f4_multd_L_himul_n284,
         SBOX_Inst_f4_multd_L_himul_n283, SBOX_Inst_f4_multd_L_himul_n282,
         SBOX_Inst_f4_multd_L_himul_n281, SBOX_Inst_f4_multd_L_himul_n280,
         SBOX_Inst_f4_multd_L_himul_n279, SBOX_Inst_f4_multd_L_himul_n278,
         SBOX_Inst_f4_multd_L_himul_n277, SBOX_Inst_f4_multd_L_himul_n276,
         SBOX_Inst_f4_multd_L_himul_n275, SBOX_Inst_f4_multd_L_himul_n274,
         SBOX_Inst_f4_multd_L_himul_n273, SBOX_Inst_f4_multd_L_himul_n272,
         SBOX_Inst_f4_multd_L_himul_n271, SBOX_Inst_f4_multd_L_himul_n270,
         SBOX_Inst_f4_multd_L_himul_n269, SBOX_Inst_f4_multd_L_himul_n268,
         SBOX_Inst_f4_multd_L_himul_n267, SBOX_Inst_f4_multd_L_himul_n266,
         SBOX_Inst_f4_multd_L_himul_n265, SBOX_Inst_f4_multd_L_himul_n264,
         SBOX_Inst_f4_multd_L_himul_n263, SBOX_Inst_f4_multd_L_himul_n262,
         SBOX_Inst_f4_multd_L_himul_n261, SBOX_Inst_f4_multd_L_himul_n260,
         SBOX_Inst_f4_multd_L_himul_n259, SBOX_Inst_f4_multd_L_himul_n258,
         SBOX_Inst_f4_multd_L_himul_n257, SBOX_Inst_f4_multd_L_himul_n256,
         SBOX_Inst_f4_multd_L_himul_n255, SBOX_Inst_f4_multd_L_himul_n254,
         SBOX_Inst_f4_multd_L_himul_n253, SBOX_Inst_f4_multd_L_himul_n252,
         SBOX_Inst_f4_multd_L_himul_n251, SBOX_Inst_f4_multd_L_himul_n250,
         SBOX_Inst_f4_multd_L_himul_n249, SBOX_Inst_f4_multd_L_himul_n248,
         SBOX_Inst_f4_multd_L_himul_n247, SBOX_Inst_f4_multd_L_himul_n246,
         SBOX_Inst_f4_multd_L_himul_n245, SBOX_Inst_f4_multd_L_himul_n244,
         SBOX_Inst_f4_multd_L_himul_n243, SBOX_Inst_f4_multd_L_himul_n242,
         SBOX_Inst_f4_multd_L_himul_n241, SBOX_Inst_f4_multd_L_himul_n240,
         SBOX_Inst_f4_multd_L_himul_n239, SBOX_Inst_f4_multd_L_himul_n238,
         SBOX_Inst_f4_multd_L_himul_n237, SBOX_Inst_f4_multd_L_himul_n236,
         SBOX_Inst_f4_multd_L_himul_n235, SBOX_Inst_f4_multd_L_himul_n234,
         SBOX_Inst_f4_multd_L_himul_n233, SBOX_Inst_f4_multd_L_himul_n232,
         SBOX_Inst_f4_multd_L_himul_n231, SBOX_Inst_f4_multd_L_himul_n230,
         SBOX_Inst_f4_multd_L_himul_n229, SBOX_Inst_f4_multd_L_himul_n228,
         SBOX_Inst_f4_multd_L_himul_n227, SBOX_Inst_f4_multd_L_himul_n226,
         SBOX_Inst_f4_multd_L_himul_n225, SBOX_Inst_f4_multd_L_himul_n224,
         SBOX_Inst_f4_multd_L_himul_n223, SBOX_Inst_f4_multd_L_himul_n222,
         SBOX_Inst_f4_multd_L_himul_n221, SBOX_Inst_f4_multd_L_himul_n220,
         SBOX_Inst_f4_multd_L_himul_n219, SBOX_Inst_f4_multd_L_himul_n218,
         SBOX_Inst_f4_multd_L_himul_n217, SBOX_Inst_f4_multd_L_himul_n216,
         SBOX_Inst_f4_multd_L_AddNewMaskph_n6,
         SBOX_Inst_f4_multd_L_AddNewMaskph_n5,
         SBOX_Inst_f4_multd_L_summul_n298, SBOX_Inst_f4_multd_L_summul_n297,
         SBOX_Inst_f4_multd_L_summul_n296, SBOX_Inst_f4_multd_L_summul_n295,
         SBOX_Inst_f4_multd_L_summul_n294, SBOX_Inst_f4_multd_L_summul_n293,
         SBOX_Inst_f4_multd_L_summul_n292, SBOX_Inst_f4_multd_L_summul_n291,
         SBOX_Inst_f4_multd_L_summul_n290, SBOX_Inst_f4_multd_L_summul_n289,
         SBOX_Inst_f4_multd_L_summul_n288, SBOX_Inst_f4_multd_L_summul_n287,
         SBOX_Inst_f4_multd_L_summul_n286, SBOX_Inst_f4_multd_L_summul_n285,
         SBOX_Inst_f4_multd_L_summul_n284, SBOX_Inst_f4_multd_L_summul_n283,
         SBOX_Inst_f4_multd_L_summul_n282, SBOX_Inst_f4_multd_L_summul_n281,
         SBOX_Inst_f4_multd_L_summul_n280, SBOX_Inst_f4_multd_L_summul_n279,
         SBOX_Inst_f4_multd_L_summul_n278, SBOX_Inst_f4_multd_L_summul_n277,
         SBOX_Inst_f4_multd_L_summul_n276, SBOX_Inst_f4_multd_L_summul_n275,
         SBOX_Inst_f4_multd_L_summul_n274, SBOX_Inst_f4_multd_L_summul_n273,
         SBOX_Inst_f4_multd_L_summul_n272, SBOX_Inst_f4_multd_L_summul_n271,
         SBOX_Inst_f4_multd_L_summul_n270, SBOX_Inst_f4_multd_L_summul_n269,
         SBOX_Inst_f4_multd_L_summul_n268, SBOX_Inst_f4_multd_L_summul_n267,
         SBOX_Inst_f4_multd_L_summul_n266, SBOX_Inst_f4_multd_L_summul_n265,
         SBOX_Inst_f4_multd_L_summul_n264, SBOX_Inst_f4_multd_L_summul_n263,
         SBOX_Inst_f4_multd_L_summul_n262, SBOX_Inst_f4_multd_L_summul_n261,
         SBOX_Inst_f4_multd_L_summul_n260, SBOX_Inst_f4_multd_L_summul_n259,
         SBOX_Inst_f4_multd_L_summul_n258, SBOX_Inst_f4_multd_L_summul_n257,
         SBOX_Inst_f4_multd_L_summul_n256, SBOX_Inst_f4_multd_L_summul_n255,
         SBOX_Inst_f4_multd_L_summul_n254, SBOX_Inst_f4_multd_L_summul_n253,
         SBOX_Inst_f4_multd_L_summul_n252, SBOX_Inst_f4_multd_L_summul_n251,
         SBOX_Inst_f4_multd_L_summul_n250, SBOX_Inst_f4_multd_L_summul_n249,
         SBOX_Inst_f4_multd_L_summul_n248, SBOX_Inst_f4_multd_L_summul_n247,
         SBOX_Inst_f4_multd_L_summul_n246, SBOX_Inst_f4_multd_L_summul_n245,
         SBOX_Inst_f4_multd_L_summul_n244, SBOX_Inst_f4_multd_L_summul_n243,
         SBOX_Inst_f4_multd_L_summul_n242, SBOX_Inst_f4_multd_L_summul_n241,
         SBOX_Inst_f4_multd_L_summul_n240, SBOX_Inst_f4_multd_L_summul_n239,
         SBOX_Inst_f4_multd_L_summul_n238, SBOX_Inst_f4_multd_L_summul_n237,
         SBOX_Inst_f4_multd_L_summul_n236, SBOX_Inst_f4_multd_L_summul_n235,
         SBOX_Inst_f4_multd_L_summul_n234, SBOX_Inst_f4_multd_L_summul_n233,
         SBOX_Inst_f4_multd_L_summul_n232, SBOX_Inst_f4_multd_L_summul_n231,
         SBOX_Inst_f4_multd_L_summul_n230, SBOX_Inst_f4_multd_L_summul_n229,
         SBOX_Inst_f4_multd_L_summul_n228, SBOX_Inst_f4_multd_L_summul_n227,
         SBOX_Inst_f4_multd_L_summul_n226, SBOX_Inst_f4_multd_L_summul_n225,
         SBOX_Inst_f4_multd_L_summul_n224, SBOX_Inst_f4_multd_L_summul_n223,
         SBOX_Inst_f4_multd_L_summul_n222, SBOX_Inst_f4_multd_L_summul_n221,
         SBOX_Inst_f4_multd_L_summul_n220, SBOX_Inst_f4_multd_L_summul_n219,
         SBOX_Inst_f4_multd_L_summul_n218, SBOX_Inst_f4_multd_L_summul_n217,
         SBOX_Inst_f4_multd_L_summul_n216, SBOX_Inst_f4_multd_L_summul_n215,
         SBOX_Inst_f4_multd_L_AddNewMaskp_n6,
         SBOX_Inst_f4_multd_L_AddNewMaskp_n5, SBOX_Inst_f4_multd_L_lowmul_n302,
         SBOX_Inst_f4_multd_L_lowmul_n301, SBOX_Inst_f4_multd_L_lowmul_n300,
         SBOX_Inst_f4_multd_L_lowmul_n299, SBOX_Inst_f4_multd_L_lowmul_n298,
         SBOX_Inst_f4_multd_L_lowmul_n297, SBOX_Inst_f4_multd_L_lowmul_n296,
         SBOX_Inst_f4_multd_L_lowmul_n295, SBOX_Inst_f4_multd_L_lowmul_n294,
         SBOX_Inst_f4_multd_L_lowmul_n293, SBOX_Inst_f4_multd_L_lowmul_n292,
         SBOX_Inst_f4_multd_L_lowmul_n291, SBOX_Inst_f4_multd_L_lowmul_n290,
         SBOX_Inst_f4_multd_L_lowmul_n289, SBOX_Inst_f4_multd_L_lowmul_n288,
         SBOX_Inst_f4_multd_L_lowmul_n287, SBOX_Inst_f4_multd_L_lowmul_n286,
         SBOX_Inst_f4_multd_L_lowmul_n285, SBOX_Inst_f4_multd_L_lowmul_n284,
         SBOX_Inst_f4_multd_L_lowmul_n283, SBOX_Inst_f4_multd_L_lowmul_n282,
         SBOX_Inst_f4_multd_L_lowmul_n281, SBOX_Inst_f4_multd_L_lowmul_n280,
         SBOX_Inst_f4_multd_L_lowmul_n279, SBOX_Inst_f4_multd_L_lowmul_n278,
         SBOX_Inst_f4_multd_L_lowmul_n277, SBOX_Inst_f4_multd_L_lowmul_n276,
         SBOX_Inst_f4_multd_L_lowmul_n275, SBOX_Inst_f4_multd_L_lowmul_n274,
         SBOX_Inst_f4_multd_L_lowmul_n273, SBOX_Inst_f4_multd_L_lowmul_n272,
         SBOX_Inst_f4_multd_L_lowmul_n271, SBOX_Inst_f4_multd_L_lowmul_n270,
         SBOX_Inst_f4_multd_L_lowmul_n269, SBOX_Inst_f4_multd_L_lowmul_n268,
         SBOX_Inst_f4_multd_L_lowmul_n267, SBOX_Inst_f4_multd_L_lowmul_n266,
         SBOX_Inst_f4_multd_L_lowmul_n265, SBOX_Inst_f4_multd_L_lowmul_n264,
         SBOX_Inst_f4_multd_L_lowmul_n263, SBOX_Inst_f4_multd_L_lowmul_n262,
         SBOX_Inst_f4_multd_L_lowmul_n261, SBOX_Inst_f4_multd_L_lowmul_n260,
         SBOX_Inst_f4_multd_L_lowmul_n259, SBOX_Inst_f4_multd_L_lowmul_n258,
         SBOX_Inst_f4_multd_L_lowmul_n257, SBOX_Inst_f4_multd_L_lowmul_n256,
         SBOX_Inst_f4_multd_L_lowmul_n255, SBOX_Inst_f4_multd_L_lowmul_n254,
         SBOX_Inst_f4_multd_L_lowmul_n253, SBOX_Inst_f4_multd_L_lowmul_n252,
         SBOX_Inst_f4_multd_L_lowmul_n251, SBOX_Inst_f4_multd_L_lowmul_n250,
         SBOX_Inst_f4_multd_L_lowmul_n249, SBOX_Inst_f4_multd_L_lowmul_n248,
         SBOX_Inst_f4_multd_L_lowmul_n247, SBOX_Inst_f4_multd_L_lowmul_n246,
         SBOX_Inst_f4_multd_L_lowmul_n245, SBOX_Inst_f4_multd_L_lowmul_n244,
         SBOX_Inst_f4_multd_L_lowmul_n243, SBOX_Inst_f4_multd_L_lowmul_n242,
         SBOX_Inst_f4_multd_L_lowmul_n241, SBOX_Inst_f4_multd_L_lowmul_n240,
         SBOX_Inst_f4_multd_L_lowmul_n239, SBOX_Inst_f4_multd_L_lowmul_n238,
         SBOX_Inst_f4_multd_L_lowmul_n237, SBOX_Inst_f4_multd_L_lowmul_n236,
         SBOX_Inst_f4_multd_L_lowmul_n235, SBOX_Inst_f4_multd_L_lowmul_n234,
         SBOX_Inst_f4_multd_L_lowmul_n233, SBOX_Inst_f4_multd_L_lowmul_n232,
         SBOX_Inst_f4_multd_L_lowmul_n231, SBOX_Inst_f4_multd_L_lowmul_n230,
         SBOX_Inst_f4_multd_L_lowmul_n229, SBOX_Inst_f4_multd_L_lowmul_n228,
         SBOX_Inst_f4_multd_L_lowmul_n227, SBOX_Inst_f4_multd_L_lowmul_n226,
         SBOX_Inst_f4_multd_L_lowmul_n225, SBOX_Inst_f4_multd_L_lowmul_n224,
         SBOX_Inst_f4_multd_L_lowmul_n223, SBOX_Inst_f4_multd_L_lowmul_n222,
         SBOX_Inst_f4_multd_L_lowmul_n221, SBOX_Inst_f4_multd_L_lowmul_n220,
         SBOX_Inst_f4_multd_L_lowmul_n219, SBOX_Inst_f4_multd_L_lowmul_n218,
         SBOX_Inst_f4_multd_L_lowmul_n217, SBOX_Inst_f4_multd_L_lowmul_n216,
         SBOX_Inst_f4_multd_L_AddNewMaskpl_n6,
         SBOX_Inst_f4_multd_L_AddNewMaskpl_n5, SBOX_Inst_f4_multd_H_himul_n308,
         SBOX_Inst_f4_multd_H_himul_n307, SBOX_Inst_f4_multd_H_himul_n306,
         SBOX_Inst_f4_multd_H_himul_n305, SBOX_Inst_f4_multd_H_himul_n304,
         SBOX_Inst_f4_multd_H_himul_n303, SBOX_Inst_f4_multd_H_himul_n302,
         SBOX_Inst_f4_multd_H_himul_n301, SBOX_Inst_f4_multd_H_himul_n300,
         SBOX_Inst_f4_multd_H_himul_n299, SBOX_Inst_f4_multd_H_himul_n298,
         SBOX_Inst_f4_multd_H_himul_n297, SBOX_Inst_f4_multd_H_himul_n296,
         SBOX_Inst_f4_multd_H_himul_n295, SBOX_Inst_f4_multd_H_himul_n294,
         SBOX_Inst_f4_multd_H_himul_n293, SBOX_Inst_f4_multd_H_himul_n292,
         SBOX_Inst_f4_multd_H_himul_n291, SBOX_Inst_f4_multd_H_himul_n290,
         SBOX_Inst_f4_multd_H_himul_n289, SBOX_Inst_f4_multd_H_himul_n288,
         SBOX_Inst_f4_multd_H_himul_n287, SBOX_Inst_f4_multd_H_himul_n286,
         SBOX_Inst_f4_multd_H_himul_n285, SBOX_Inst_f4_multd_H_himul_n284,
         SBOX_Inst_f4_multd_H_himul_n283, SBOX_Inst_f4_multd_H_himul_n282,
         SBOX_Inst_f4_multd_H_himul_n281, SBOX_Inst_f4_multd_H_himul_n280,
         SBOX_Inst_f4_multd_H_himul_n279, SBOX_Inst_f4_multd_H_himul_n278,
         SBOX_Inst_f4_multd_H_himul_n277, SBOX_Inst_f4_multd_H_himul_n276,
         SBOX_Inst_f4_multd_H_himul_n275, SBOX_Inst_f4_multd_H_himul_n274,
         SBOX_Inst_f4_multd_H_himul_n273, SBOX_Inst_f4_multd_H_himul_n272,
         SBOX_Inst_f4_multd_H_himul_n271, SBOX_Inst_f4_multd_H_himul_n270,
         SBOX_Inst_f4_multd_H_himul_n269, SBOX_Inst_f4_multd_H_himul_n268,
         SBOX_Inst_f4_multd_H_himul_n267, SBOX_Inst_f4_multd_H_himul_n266,
         SBOX_Inst_f4_multd_H_himul_n265, SBOX_Inst_f4_multd_H_himul_n264,
         SBOX_Inst_f4_multd_H_himul_n263, SBOX_Inst_f4_multd_H_himul_n262,
         SBOX_Inst_f4_multd_H_himul_n261, SBOX_Inst_f4_multd_H_himul_n260,
         SBOX_Inst_f4_multd_H_himul_n259, SBOX_Inst_f4_multd_H_himul_n258,
         SBOX_Inst_f4_multd_H_himul_n257, SBOX_Inst_f4_multd_H_himul_n256,
         SBOX_Inst_f4_multd_H_himul_n255, SBOX_Inst_f4_multd_H_himul_n254,
         SBOX_Inst_f4_multd_H_himul_n253, SBOX_Inst_f4_multd_H_himul_n252,
         SBOX_Inst_f4_multd_H_himul_n251, SBOX_Inst_f4_multd_H_himul_n250,
         SBOX_Inst_f4_multd_H_himul_n249, SBOX_Inst_f4_multd_H_himul_n248,
         SBOX_Inst_f4_multd_H_himul_n247, SBOX_Inst_f4_multd_H_himul_n246,
         SBOX_Inst_f4_multd_H_himul_n245, SBOX_Inst_f4_multd_H_himul_n244,
         SBOX_Inst_f4_multd_H_himul_n243, SBOX_Inst_f4_multd_H_himul_n242,
         SBOX_Inst_f4_multd_H_himul_n241, SBOX_Inst_f4_multd_H_himul_n240,
         SBOX_Inst_f4_multd_H_himul_n239, SBOX_Inst_f4_multd_H_himul_n238,
         SBOX_Inst_f4_multd_H_himul_n237, SBOX_Inst_f4_multd_H_himul_n236,
         SBOX_Inst_f4_multd_H_himul_n235, SBOX_Inst_f4_multd_H_himul_n234,
         SBOX_Inst_f4_multd_H_himul_n233, SBOX_Inst_f4_multd_H_himul_n232,
         SBOX_Inst_f4_multd_H_himul_n231, SBOX_Inst_f4_multd_H_himul_n230,
         SBOX_Inst_f4_multd_H_himul_n229, SBOX_Inst_f4_multd_H_himul_n228,
         SBOX_Inst_f4_multd_H_himul_n227, SBOX_Inst_f4_multd_H_himul_n226,
         SBOX_Inst_f4_multd_H_himul_n225, SBOX_Inst_f4_multd_H_himul_n224,
         SBOX_Inst_f4_multd_H_himul_n223, SBOX_Inst_f4_multd_H_himul_n222,
         SBOX_Inst_f4_multd_H_himul_n221, SBOX_Inst_f4_multd_H_himul_n220,
         SBOX_Inst_f4_multd_H_himul_n219, SBOX_Inst_f4_multd_H_himul_n218,
         SBOX_Inst_f4_multd_H_himul_n217, SBOX_Inst_f4_multd_H_himul_n216,
         SBOX_Inst_f4_multd_H_himul_n215, SBOX_Inst_f4_multd_H_AddNewMaskph_n6,
         SBOX_Inst_f4_multd_H_AddNewMaskph_n5,
         SBOX_Inst_f4_multd_H_summul_n308, SBOX_Inst_f4_multd_H_summul_n307,
         SBOX_Inst_f4_multd_H_summul_n306, SBOX_Inst_f4_multd_H_summul_n305,
         SBOX_Inst_f4_multd_H_summul_n304, SBOX_Inst_f4_multd_H_summul_n303,
         SBOX_Inst_f4_multd_H_summul_n302, SBOX_Inst_f4_multd_H_summul_n301,
         SBOX_Inst_f4_multd_H_summul_n300, SBOX_Inst_f4_multd_H_summul_n299,
         SBOX_Inst_f4_multd_H_summul_n298, SBOX_Inst_f4_multd_H_summul_n297,
         SBOX_Inst_f4_multd_H_summul_n296, SBOX_Inst_f4_multd_H_summul_n295,
         SBOX_Inst_f4_multd_H_summul_n294, SBOX_Inst_f4_multd_H_summul_n293,
         SBOX_Inst_f4_multd_H_summul_n292, SBOX_Inst_f4_multd_H_summul_n291,
         SBOX_Inst_f4_multd_H_summul_n290, SBOX_Inst_f4_multd_H_summul_n289,
         SBOX_Inst_f4_multd_H_summul_n288, SBOX_Inst_f4_multd_H_summul_n287,
         SBOX_Inst_f4_multd_H_summul_n286, SBOX_Inst_f4_multd_H_summul_n285,
         SBOX_Inst_f4_multd_H_summul_n284, SBOX_Inst_f4_multd_H_summul_n283,
         SBOX_Inst_f4_multd_H_summul_n282, SBOX_Inst_f4_multd_H_summul_n281,
         SBOX_Inst_f4_multd_H_summul_n280, SBOX_Inst_f4_multd_H_summul_n279,
         SBOX_Inst_f4_multd_H_summul_n278, SBOX_Inst_f4_multd_H_summul_n277,
         SBOX_Inst_f4_multd_H_summul_n276, SBOX_Inst_f4_multd_H_summul_n275,
         SBOX_Inst_f4_multd_H_summul_n274, SBOX_Inst_f4_multd_H_summul_n273,
         SBOX_Inst_f4_multd_H_summul_n272, SBOX_Inst_f4_multd_H_summul_n271,
         SBOX_Inst_f4_multd_H_summul_n270, SBOX_Inst_f4_multd_H_summul_n269,
         SBOX_Inst_f4_multd_H_summul_n268, SBOX_Inst_f4_multd_H_summul_n267,
         SBOX_Inst_f4_multd_H_summul_n266, SBOX_Inst_f4_multd_H_summul_n265,
         SBOX_Inst_f4_multd_H_summul_n264, SBOX_Inst_f4_multd_H_summul_n263,
         SBOX_Inst_f4_multd_H_summul_n262, SBOX_Inst_f4_multd_H_summul_n261,
         SBOX_Inst_f4_multd_H_summul_n260, SBOX_Inst_f4_multd_H_summul_n259,
         SBOX_Inst_f4_multd_H_summul_n258, SBOX_Inst_f4_multd_H_summul_n257,
         SBOX_Inst_f4_multd_H_summul_n256, SBOX_Inst_f4_multd_H_summul_n255,
         SBOX_Inst_f4_multd_H_summul_n254, SBOX_Inst_f4_multd_H_summul_n253,
         SBOX_Inst_f4_multd_H_summul_n252, SBOX_Inst_f4_multd_H_summul_n251,
         SBOX_Inst_f4_multd_H_summul_n250, SBOX_Inst_f4_multd_H_summul_n249,
         SBOX_Inst_f4_multd_H_summul_n248, SBOX_Inst_f4_multd_H_summul_n247,
         SBOX_Inst_f4_multd_H_summul_n246, SBOX_Inst_f4_multd_H_summul_n245,
         SBOX_Inst_f4_multd_H_summul_n244, SBOX_Inst_f4_multd_H_summul_n243,
         SBOX_Inst_f4_multd_H_summul_n242, SBOX_Inst_f4_multd_H_summul_n241,
         SBOX_Inst_f4_multd_H_summul_n240, SBOX_Inst_f4_multd_H_summul_n239,
         SBOX_Inst_f4_multd_H_summul_n238, SBOX_Inst_f4_multd_H_summul_n237,
         SBOX_Inst_f4_multd_H_summul_n236, SBOX_Inst_f4_multd_H_summul_n235,
         SBOX_Inst_f4_multd_H_summul_n234, SBOX_Inst_f4_multd_H_summul_n233,
         SBOX_Inst_f4_multd_H_summul_n232, SBOX_Inst_f4_multd_H_summul_n231,
         SBOX_Inst_f4_multd_H_summul_n230, SBOX_Inst_f4_multd_H_summul_n229,
         SBOX_Inst_f4_multd_H_summul_n228, SBOX_Inst_f4_multd_H_summul_n227,
         SBOX_Inst_f4_multd_H_summul_n226, SBOX_Inst_f4_multd_H_summul_n225,
         SBOX_Inst_f4_multd_H_summul_n224, SBOX_Inst_f4_multd_H_summul_n223,
         SBOX_Inst_f4_multd_H_summul_n222, SBOX_Inst_f4_multd_H_summul_n221,
         SBOX_Inst_f4_multd_H_summul_n220, SBOX_Inst_f4_multd_H_summul_n219,
         SBOX_Inst_f4_multd_H_summul_n218, SBOX_Inst_f4_multd_H_summul_n217,
         SBOX_Inst_f4_multd_H_summul_n216, SBOX_Inst_f4_multd_H_summul_n215,
         SBOX_Inst_f4_multd_H_AddNewMaskp_n6,
         SBOX_Inst_f4_multd_H_AddNewMaskp_n5, SBOX_Inst_f4_multd_H_lowmul_n308,
         SBOX_Inst_f4_multd_H_lowmul_n307, SBOX_Inst_f4_multd_H_lowmul_n306,
         SBOX_Inst_f4_multd_H_lowmul_n305, SBOX_Inst_f4_multd_H_lowmul_n304,
         SBOX_Inst_f4_multd_H_lowmul_n303, SBOX_Inst_f4_multd_H_lowmul_n302,
         SBOX_Inst_f4_multd_H_lowmul_n301, SBOX_Inst_f4_multd_H_lowmul_n300,
         SBOX_Inst_f4_multd_H_lowmul_n299, SBOX_Inst_f4_multd_H_lowmul_n298,
         SBOX_Inst_f4_multd_H_lowmul_n297, SBOX_Inst_f4_multd_H_lowmul_n296,
         SBOX_Inst_f4_multd_H_lowmul_n295, SBOX_Inst_f4_multd_H_lowmul_n294,
         SBOX_Inst_f4_multd_H_lowmul_n293, SBOX_Inst_f4_multd_H_lowmul_n292,
         SBOX_Inst_f4_multd_H_lowmul_n291, SBOX_Inst_f4_multd_H_lowmul_n290,
         SBOX_Inst_f4_multd_H_lowmul_n289, SBOX_Inst_f4_multd_H_lowmul_n288,
         SBOX_Inst_f4_multd_H_lowmul_n287, SBOX_Inst_f4_multd_H_lowmul_n286,
         SBOX_Inst_f4_multd_H_lowmul_n285, SBOX_Inst_f4_multd_H_lowmul_n284,
         SBOX_Inst_f4_multd_H_lowmul_n283, SBOX_Inst_f4_multd_H_lowmul_n282,
         SBOX_Inst_f4_multd_H_lowmul_n281, SBOX_Inst_f4_multd_H_lowmul_n280,
         SBOX_Inst_f4_multd_H_lowmul_n279, SBOX_Inst_f4_multd_H_lowmul_n278,
         SBOX_Inst_f4_multd_H_lowmul_n277, SBOX_Inst_f4_multd_H_lowmul_n276,
         SBOX_Inst_f4_multd_H_lowmul_n275, SBOX_Inst_f4_multd_H_lowmul_n274,
         SBOX_Inst_f4_multd_H_lowmul_n273, SBOX_Inst_f4_multd_H_lowmul_n272,
         SBOX_Inst_f4_multd_H_lowmul_n271, SBOX_Inst_f4_multd_H_lowmul_n270,
         SBOX_Inst_f4_multd_H_lowmul_n269, SBOX_Inst_f4_multd_H_lowmul_n268,
         SBOX_Inst_f4_multd_H_lowmul_n267, SBOX_Inst_f4_multd_H_lowmul_n266,
         SBOX_Inst_f4_multd_H_lowmul_n265, SBOX_Inst_f4_multd_H_lowmul_n264,
         SBOX_Inst_f4_multd_H_lowmul_n263, SBOX_Inst_f4_multd_H_lowmul_n262,
         SBOX_Inst_f4_multd_H_lowmul_n261, SBOX_Inst_f4_multd_H_lowmul_n260,
         SBOX_Inst_f4_multd_H_lowmul_n259, SBOX_Inst_f4_multd_H_lowmul_n258,
         SBOX_Inst_f4_multd_H_lowmul_n257, SBOX_Inst_f4_multd_H_lowmul_n256,
         SBOX_Inst_f4_multd_H_lowmul_n255, SBOX_Inst_f4_multd_H_lowmul_n254,
         SBOX_Inst_f4_multd_H_lowmul_n253, SBOX_Inst_f4_multd_H_lowmul_n252,
         SBOX_Inst_f4_multd_H_lowmul_n251, SBOX_Inst_f4_multd_H_lowmul_n250,
         SBOX_Inst_f4_multd_H_lowmul_n249, SBOX_Inst_f4_multd_H_lowmul_n248,
         SBOX_Inst_f4_multd_H_lowmul_n247, SBOX_Inst_f4_multd_H_lowmul_n246,
         SBOX_Inst_f4_multd_H_lowmul_n245, SBOX_Inst_f4_multd_H_lowmul_n244,
         SBOX_Inst_f4_multd_H_lowmul_n243, SBOX_Inst_f4_multd_H_lowmul_n242,
         SBOX_Inst_f4_multd_H_lowmul_n241, SBOX_Inst_f4_multd_H_lowmul_n240,
         SBOX_Inst_f4_multd_H_lowmul_n239, SBOX_Inst_f4_multd_H_lowmul_n238,
         SBOX_Inst_f4_multd_H_lowmul_n237, SBOX_Inst_f4_multd_H_lowmul_n236,
         SBOX_Inst_f4_multd_H_lowmul_n235, SBOX_Inst_f4_multd_H_lowmul_n234,
         SBOX_Inst_f4_multd_H_lowmul_n233, SBOX_Inst_f4_multd_H_lowmul_n232,
         SBOX_Inst_f4_multd_H_lowmul_n231, SBOX_Inst_f4_multd_H_lowmul_n230,
         SBOX_Inst_f4_multd_H_lowmul_n229, SBOX_Inst_f4_multd_H_lowmul_n228,
         SBOX_Inst_f4_multd_H_lowmul_n227, SBOX_Inst_f4_multd_H_lowmul_n226,
         SBOX_Inst_f4_multd_H_lowmul_n225, SBOX_Inst_f4_multd_H_lowmul_n224,
         SBOX_Inst_f4_multd_H_lowmul_n223, SBOX_Inst_f4_multd_H_lowmul_n222,
         SBOX_Inst_f4_multd_H_lowmul_n221, SBOX_Inst_f4_multd_H_lowmul_n220,
         SBOX_Inst_f4_multd_H_lowmul_n219, SBOX_Inst_f4_multd_H_lowmul_n218,
         SBOX_Inst_f4_multd_H_lowmul_n217, SBOX_Inst_f4_multd_H_lowmul_n216,
         SBOX_Inst_f4_multd_H_lowmul_n215,
         SBOX_Inst_f4_multd_H_AddNewMaskpl_n6,
         SBOX_Inst_f4_multd_H_AddNewMaskpl_n5, SBOX_PL_4_n252, SBOX_PL_4_n251,
         SBOX_PL_4_n250, SBOX_PL_4_n249, SBOX_PL_4_n248, SBOX_PL_4_n247,
         SBOX_PL_4_n246, SBOX_PL_4_n245, SBOX_PL_4_n244, SBOX_PL_4_n243,
         SBOX_PL_4_n242, SBOX_PL_4_n241, SBOX_PL_4_n240, SBOX_PL_4_n239,
         SBOX_PL_4_n238, SBOX_PL_4_n237, SBOX_PL_4_n236, SBOX_PL_4_n235,
         SBOX_PL_4_n234, SBOX_PL_4_n233, SBOX_PL_4_n232, SBOX_PL_4_n231,
         SBOX_PL_4_n230, SBOX_PL_4_n229, SBOX_PL_4_n228, SBOX_PL_4_n227,
         SBOX_PL_4_n226, SBOX_PL_4_n225, SBOX_PL_4_n224, SBOX_PL_4_n223,
         SBOX_PL_4_n222, SBOX_PL_4_n221, SBOX_PL_4_n220, SBOX_PL_4_n219,
         SBOX_PL_4_n218, SBOX_PL_4_n217, SBOX_PL_4_n180, SBOX_PL_4_n179,
         SBOX_PL_4_n178, SBOX_PL_4_n177, SBOX_PL_4_n176, SBOX_PL_4_n175,
         SBOX_PL_4_n174, SBOX_PL_4_n173, SBOX_PL_4_n172, SBOX_PL_4_n171,
         SBOX_PL_4_n170, SBOX_PL_4_n169, SBOX_PL_4_n168, SBOX_PL_4_n167,
         SBOX_PL_4_n166, SBOX_PL_4_n165, SBOX_PL_4_n164, SBOX_PL_4_n163,
         SBOX_PL_4_n162, SBOX_PL_4_n161, SBOX_PL_4_n160, SBOX_PL_4_n159,
         SBOX_PL_4_n158, SBOX_PL_4_n157, SBOX_PL_4_n156, SBOX_PL_4_n155,
         SBOX_PL_4_n154, SBOX_PL_4_n153, SBOX_PL_4_n152, SBOX_PL_4_n151,
         SBOX_PL_4_n150, SBOX_PL_4_n149, SBOX_PL_4_n148, SBOX_PL_4_n147,
         SBOX_PL_4_n146, SBOX_PL_4_n145, SBOX_PL_4_n144, SBOX_PL_4_n143,
         SBOX_PL_4_n142, SBOX_PL_4_n141, SBOX_PL_4_n140, SBOX_PL_4_n139,
         SBOX_PL_4_n138, SBOX_PL_4_n137, SBOX_PL_4_n136, SBOX_PL_4_n135,
         SBOX_PL_4_n134, SBOX_PL_4_n133, SBOX_PL_4_n132, SBOX_PL_4_n131,
         SBOX_PL_4_n130, SBOX_PL_4_n129, SBOX_PL_4_n128, SBOX_PL_4_n127,
         SBOX_PL_4_n126, SBOX_PL_4_n125, SBOX_PL_4_n124, SBOX_PL_4_n123,
         SBOX_PL_4_n122, SBOX_PL_4_n121, SBOX_PL_4_n120, SBOX_PL_4_n119,
         SBOX_PL_4_n118, SBOX_PL_4_n117, SBOX_PL_4_n116, SBOX_PL_4_n115,
         SBOX_PL_4_n114, SBOX_PL_4_n113, SBOX_PL_4_n112, SBOX_PL_4_n111,
         SBOX_PL_4_n110, SBOX_PL_4_n109, SBOX_Inst_f5_phwillwin_pw2_0_,
         SBOX_Inst_f5_phwillwin_pw2_1_, SBOX_Inst_f5_phwillwin_pw2_2_,
         SBOX_Inst_f5_phwillwin_pw2_3_, SBOX_Inst_f5_phwillwin_pw2_4_,
         SBOX_Inst_f5_phwillwin_pw2_5_, SBOX_Inst_f5_plwillwin_pw2_0_,
         SBOX_Inst_f5_plwillwin_pw2_1_, SBOX_Inst_f5_plwillwin_pw2_2_,
         SBOX_Inst_f5_plwillwin_pw2_3_, SBOX_Inst_f5_plwillwin_pw2_4_,
         SBOX_Inst_f5_plwillwin_pw2_5_, SBOX_Inst_f5_invlinearMapping_n9,
         SBOX_Inst_f5_invlinearMapping_n8, SBOX_Inst_f5_invlinearMapping_n7,
         SBOX_Inst_f5_invlinearMapping_n6, SBOX_Inst_f5_invlinearMapping_n5,
         SBOX_Inst_f5_invlinearMapping_n4, SBOX_Inst_f5_invlinearMapping_n3,
         SBOX_Inst_f5_invlinearMapping_n2, SBOX_Inst_f5_invlinearMapping_n1,
         SBOX_PL_5_n168, SBOX_PL_5_n167, SBOX_PL_5_n166, SBOX_PL_5_n165,
         SBOX_PL_5_n164, SBOX_PL_5_n163, SBOX_PL_5_n162, SBOX_PL_5_n161,
         SBOX_PL_5_n160, SBOX_PL_5_n159, SBOX_PL_5_n158, SBOX_PL_5_n157,
         SBOX_PL_5_n156, SBOX_PL_5_n155, SBOX_PL_5_n154, SBOX_PL_5_n153,
         SBOX_PL_5_n152, SBOX_PL_5_n151, SBOX_PL_5_n150, SBOX_PL_5_n149,
         SBOX_PL_5_n148, SBOX_PL_5_n147, SBOX_PL_5_n146, SBOX_PL_5_n145,
         SBOX_PL_5_n120, SBOX_PL_5_n119, SBOX_PL_5_n118, SBOX_PL_5_n117,
         SBOX_PL_5_n116, SBOX_PL_5_n115, SBOX_PL_5_n114, SBOX_PL_5_n113,
         SBOX_PL_5_n112, SBOX_PL_5_n111, SBOX_PL_5_n110, SBOX_PL_5_n109,
         SBOX_PL_5_n108, SBOX_PL_5_n107, SBOX_PL_5_n106, SBOX_PL_5_n105,
         SBOX_PL_5_n104, SBOX_PL_5_n103, SBOX_PL_5_n102, SBOX_PL_5_n101,
         SBOX_PL_5_n100, SBOX_PL_5_n99, SBOX_PL_5_n98, SBOX_PL_5_n97,
         SBOX_PL_5_n96, SBOX_PL_5_n95, SBOX_PL_5_n94, SBOX_PL_5_n93,
         SBOX_PL_5_n92, SBOX_PL_5_n91, SBOX_PL_5_n90, SBOX_PL_5_n89,
         SBOX_PL_5_n88, SBOX_PL_5_n87, SBOX_PL_5_n86, SBOX_PL_5_n85,
         SBOX_PL_5_n84, SBOX_PL_5_n83, SBOX_PL_5_n82, SBOX_PL_5_n81,
         SBOX_PL_5_n80, SBOX_PL_5_n79, SBOX_PL_5_n78, SBOX_PL_5_n77,
         SBOX_PL_5_n76, SBOX_PL_5_n75, SBOX_PL_5_n74, SBOX_PL_5_n73,
         SBOX_PL_6_n168, SBOX_PL_6_n167, SBOX_PL_6_n166, SBOX_PL_6_n165,
         SBOX_PL_6_n164, SBOX_PL_6_n163, SBOX_PL_6_n162, SBOX_PL_6_n161,
         SBOX_PL_6_n160, SBOX_PL_6_n159, SBOX_PL_6_n158, SBOX_PL_6_n157,
         SBOX_PL_6_n156, SBOX_PL_6_n155, SBOX_PL_6_n154, SBOX_PL_6_n153,
         SBOX_PL_6_n152, SBOX_PL_6_n151, SBOX_PL_6_n150, SBOX_PL_6_n149,
         SBOX_PL_6_n148, SBOX_PL_6_n147, SBOX_PL_6_n146, SBOX_PL_6_n145,
         SBOX_PL_6_n120, SBOX_PL_6_n119, SBOX_PL_6_n118, SBOX_PL_6_n117,
         SBOX_PL_6_n116, SBOX_PL_6_n115, SBOX_PL_6_n114, SBOX_PL_6_n113,
         SBOX_PL_6_n112, SBOX_PL_6_n111, SBOX_PL_6_n110, SBOX_PL_6_n109,
         SBOX_PL_6_n108, SBOX_PL_6_n107, SBOX_PL_6_n106, SBOX_PL_6_n105,
         SBOX_PL_6_n104, SBOX_PL_6_n103, SBOX_PL_6_n102, SBOX_PL_6_n101,
         SBOX_PL_6_n100, SBOX_PL_6_n99, SBOX_PL_6_n98, SBOX_PL_6_n97,
         SBOX_PL_6_n96, SBOX_PL_6_n95, SBOX_PL_6_n94, SBOX_PL_6_n93,
         SBOX_PL_6_n92, SBOX_PL_6_n91, SBOX_PL_6_n90, SBOX_PL_6_n89,
         SBOX_PL_6_n88, SBOX_PL_6_n87, SBOX_PL_6_n86, SBOX_PL_6_n85,
         SBOX_PL_6_n84, SBOX_PL_6_n83, SBOX_PL_6_n82, SBOX_PL_6_n81,
         SBOX_PL_6_n80, SBOX_PL_6_n79, SBOX_PL_6_n78, SBOX_PL_6_n77,
         SBOX_PL_6_n76, SBOX_PL_6_n75, SBOX_PL_6_n74, SBOX_PL_6_n73,
         SBOX_PL_7_n168, SBOX_PL_7_n167, SBOX_PL_7_n166, SBOX_PL_7_n165,
         SBOX_PL_7_n164, SBOX_PL_7_n163, SBOX_PL_7_n162, SBOX_PL_7_n161,
         SBOX_PL_7_n160, SBOX_PL_7_n159, SBOX_PL_7_n158, SBOX_PL_7_n157,
         SBOX_PL_7_n156, SBOX_PL_7_n155, SBOX_PL_7_n154, SBOX_PL_7_n153,
         SBOX_PL_7_n152, SBOX_PL_7_n151, SBOX_PL_7_n150, SBOX_PL_7_n149,
         SBOX_PL_7_n148, SBOX_PL_7_n147, SBOX_PL_7_n146, SBOX_PL_7_n145,
         SBOX_PL_7_n120, SBOX_PL_7_n119, SBOX_PL_7_n118, SBOX_PL_7_n117,
         SBOX_PL_7_n116, SBOX_PL_7_n115, SBOX_PL_7_n114, SBOX_PL_7_n113,
         SBOX_PL_7_n112, SBOX_PL_7_n111, SBOX_PL_7_n110, SBOX_PL_7_n109,
         SBOX_PL_7_n108, SBOX_PL_7_n107, SBOX_PL_7_n106, SBOX_PL_7_n105,
         SBOX_PL_7_n104, SBOX_PL_7_n103, SBOX_PL_7_n102, SBOX_PL_7_n101,
         SBOX_PL_7_n100, SBOX_PL_7_n99, SBOX_PL_7_n98, SBOX_PL_7_n97,
         SBOX_PL_7_n96, SBOX_PL_7_n95, SBOX_PL_7_n94, SBOX_PL_7_n93,
         SBOX_PL_7_n92, SBOX_PL_7_n91, SBOX_PL_7_n90, SBOX_PL_7_n89,
         SBOX_PL_7_n88, SBOX_PL_7_n87, SBOX_PL_7_n86, SBOX_PL_7_n85,
         SBOX_PL_7_n84, SBOX_PL_7_n83, SBOX_PL_7_n82, SBOX_PL_7_n81,
         SBOX_PL_7_n80, SBOX_PL_7_n79, SBOX_PL_7_n78, SBOX_PL_7_n77,
         SBOX_PL_7_n76, SBOX_PL_7_n75, SBOX_PL_7_n74, SBOX_PL_7_n73,
         aes_key_regs_2_n3, aes_key_regs_2_K02xDP_0_, aes_key_regs_2_K02xDP_1_,
         aes_key_regs_2_K02xDP_2_, aes_key_regs_2_K02xDP_3_,
         aes_key_regs_2_K02xDP_4_, aes_key_regs_2_K02xDP_5_,
         aes_key_regs_2_K02xDP_6_, aes_key_regs_2_K02xDP_7_,
         aes_key_regs_2_K01xDP_0_, aes_key_regs_2_K01xDP_1_,
         aes_key_regs_2_K01xDP_2_, aes_key_regs_2_K01xDP_3_,
         aes_key_regs_2_K01xDP_4_, aes_key_regs_2_K01xDP_5_,
         aes_key_regs_2_K01xDP_6_, aes_key_regs_2_K01xDP_7_,
         aes_state_regs_2_n118, aes_state_regs_2_n117, aes_state_regs_2_n116,
         aes_state_regs_2_n115, aes_state_regs_2_n114, aes_state_regs_2_n113,
         aes_state_regs_2_n112, aes_state_regs_2_n111, aes_state_regs_2_n110,
         aes_state_regs_2_n109, aes_state_regs_2_n108, aes_state_regs_2_n107,
         aes_state_regs_2_n81, aes_state_regs_2_n80, aes_state_regs_2_n79,
         aes_state_regs_2_n78, aes_state_regs_2_n77, aes_state_regs_2_n76,
         aes_state_regs_2_n75, aes_state_regs_2_n74, aes_state_regs_2_n73,
         aes_state_regs_2_n72, aes_state_regs_2_n71, aes_state_regs_2_n70,
         aes_state_regs_2_n69, aes_state_regs_2_n68, aes_state_regs_2_n67,
         aes_state_regs_2_n65, aes_state_regs_2_n64, aes_state_regs_2_n63,
         aes_state_regs_2_n56, aes_state_regs_2_n46, aes_state_regs_2_n45,
         aes_state_regs_2_n105, aes_state_regs_2_n104, aes_state_regs_2_n103,
         aes_state_regs_2_n102, aes_state_regs_2_n101, aes_state_regs_2_n100,
         aes_state_regs_2_n99, aes_state_regs_2_n98, aes_state_regs_2_n97,
         aes_state_regs_2_n96, aes_state_regs_2_n95, aes_state_regs_2_n94,
         aes_state_regs_2_n93, aes_state_regs_2_n92, aes_state_regs_2_n91,
         aes_state_regs_2_n90, aes_state_regs_2_n89, aes_state_regs_2_n88,
         aes_state_regs_2_n87, aes_state_regs_2_n86, aes_state_regs_2_n85,
         aes_state_regs_2_n84, aes_state_regs_2_n83, aes_state_regs_2_n82,
         aes_state_regs_2_n66, aes_state_regs_2_n62, aes_state_regs_2_n61,
         aes_state_regs_2_n60, aes_state_regs_2_n59, aes_state_regs_2_n58,
         aes_state_regs_2_n57, aes_state_regs_2_n55, aes_state_regs_2_n54,
         aes_state_regs_2_n53, aes_state_regs_2_n52, aes_state_regs_2_n51,
         aes_state_regs_2_n50, aes_state_regs_2_n49, aes_state_regs_2_n48,
         aes_state_regs_2_n47, aes_state_regs_2_n38, aes_state_regs_2_n37,
         aes_state_regs_2_n36, aes_state_regs_2_n35, aes_state_regs_2_n34,
         aes_state_regs_2_n33, aes_state_regs_2_n32, aes_state_regs_2_n31,
         aes_state_regs_2_n30, aes_state_regs_2_n29, aes_state_regs_2_n28,
         aes_state_regs_2_n27, aes_state_regs_2_n26, aes_state_regs_2_n25,
         aes_state_regs_2_n24, aes_state_regs_2_n23, aes_state_regs_2_n22,
         aes_state_regs_2_n21, aes_state_regs_2_n20, aes_state_regs_2_n19,
         aes_state_regs_2_n18, aes_state_regs_2_n17, aes_state_regs_2_n16,
         aes_state_regs_2_n15, aes_state_regs_2_n14, aes_state_regs_2_n13,
         aes_state_regs_2_n12, aes_state_regs_2_n11, aes_state_regs_2_n10,
         aes_state_regs_2_n9, aes_state_regs_2_n8, aes_state_regs_2_n7,
         aes_state_regs_2_n6, aes_state_regs_2_n5, aes_state_regs_2_n4,
         aes_state_regs_2_n3, aes_state_regs_2_n2, aes_state_regs_2_n1,
         aes_state_regs_2_S03xDP_0_, aes_state_regs_2_S02xDP_0_,
         aes_state_regs_2_S02xDP_1_, aes_state_regs_2_S02xDP_2_,
         aes_state_regs_2_S02xDP_3_, aes_state_regs_2_S02xDP_4_,
         aes_state_regs_2_S02xDP_5_, aes_state_regs_2_S02xDP_6_,
         aes_state_regs_2_S02xDP_7_, aes_state_regs_2_S31xDP_0_,
         aes_state_regs_2_S30xDP_0_, aes_state_regs_2_S30xDP_1_,
         aes_state_regs_2_S30xDP_2_, aes_state_regs_2_S30xDP_3_,
         aes_state_regs_2_S30xDP_4_, aes_state_regs_2_S30xDP_5_,
         aes_state_regs_2_S30xDP_6_, aes_state_regs_2_S30xDP_7_,
         aes_state_regs_2_S20xDP_0_, aes_state_regs_2_S20xDP_1_,
         aes_state_regs_2_S20xDP_2_, aes_state_regs_2_S20xDP_3_,
         aes_state_regs_2_S20xDP_4_, aes_state_regs_2_S20xDP_5_,
         aes_state_regs_2_S20xDP_6_, aes_state_regs_2_S20xDP_7_,
         aes_state_regs_2_S23xDP_0_, aes_state_regs_2_S23xDP_1_,
         aes_state_regs_2_S23xDP_2_, aes_state_regs_2_S23xDP_3_,
         aes_state_regs_2_S23xDP_4_, aes_state_regs_2_S23xDP_5_,
         aes_state_regs_2_S23xDP_6_, aes_state_regs_2_S23xDP_7_,
         aes_state_regs_2_S22xDP_0_, aes_state_regs_2_S10xDP_0_,
         aes_state_regs_2_S10xDP_1_, aes_state_regs_2_S10xDP_2_,
         aes_state_regs_2_S10xDP_3_, aes_state_regs_2_S10xDP_4_,
         aes_state_regs_2_S10xDP_5_, aes_state_regs_2_S10xDP_6_,
         aes_state_regs_2_S10xDP_7_, aes_state_regs_2_S01xDO_0_,
         aes_state_regs_2_S01xDO_1_, aes_state_regs_2_S01xDO_2_,
         aes_state_regs_2_S01xDO_3_, aes_state_regs_2_S01xDO_4_,
         aes_state_regs_2_S01xDO_5_, aes_state_regs_2_S01xDO_6_,
         aes_state_regs_2_S01xDO_7_, aes_state_regs_2_mix_columns_1_n245,
         aes_state_regs_2_mix_columns_1_n244,
         aes_state_regs_2_mix_columns_1_n243,
         aes_state_regs_2_mix_columns_1_n242,
         aes_state_regs_2_mix_columns_1_n241,
         aes_state_regs_2_mix_columns_1_n240,
         aes_state_regs_2_mix_columns_1_n239,
         aes_state_regs_2_mix_columns_1_n238,
         aes_state_regs_2_mix_columns_1_n237,
         aes_state_regs_2_mix_columns_1_n236,
         aes_state_regs_2_mix_columns_1_n235,
         aes_state_regs_2_mix_columns_1_n234,
         aes_state_regs_2_mix_columns_1_n233,
         aes_state_regs_2_mix_columns_1_n232,
         aes_state_regs_2_mix_columns_1_n231,
         aes_state_regs_2_mix_columns_1_n230,
         aes_state_regs_2_mix_columns_1_n229,
         aes_state_regs_2_mix_columns_1_n228,
         aes_state_regs_2_mix_columns_1_n227,
         aes_state_regs_2_mix_columns_1_n226,
         aes_state_regs_2_mix_columns_1_n225,
         aes_state_regs_2_mix_columns_1_n224,
         aes_state_regs_2_mix_columns_1_n223,
         aes_state_regs_2_mix_columns_1_n222,
         aes_state_regs_2_mix_columns_1_n221,
         aes_state_regs_2_mix_columns_1_n220,
         aes_state_regs_2_mix_columns_1_n219,
         aes_state_regs_2_mix_columns_1_n218,
         aes_state_regs_2_mix_columns_1_n217,
         aes_state_regs_2_mix_columns_1_n216,
         aes_state_regs_2_mix_columns_1_n215,
         aes_state_regs_2_mix_columns_1_n214,
         aes_state_regs_2_mix_columns_1_n213,
         aes_state_regs_2_mix_columns_1_n212,
         aes_state_regs_2_mix_columns_1_n211,
         aes_state_regs_2_mix_columns_1_n210,
         aes_state_regs_2_mix_columns_1_n209,
         aes_state_regs_2_mix_columns_1_n208,
         aes_state_regs_2_mix_columns_1_n207,
         aes_state_regs_2_mix_columns_1_n206,
         aes_state_regs_2_mix_columns_1_n205,
         aes_state_regs_2_mix_columns_1_n204,
         aes_state_regs_2_mix_columns_1_n203,
         aes_state_regs_2_mix_columns_1_n202,
         aes_state_regs_2_mix_columns_1_n201,
         aes_state_regs_2_mix_columns_1_n200,
         aes_state_regs_2_mix_columns_1_n199,
         aes_state_regs_2_mix_columns_1_n198,
         aes_state_regs_2_mix_columns_1_n197,
         aes_state_regs_2_mix_columns_1_n196,
         aes_state_regs_2_mix_columns_1_n195,
         aes_state_regs_2_mix_columns_1_n194,
         aes_state_regs_2_mix_columns_1_n193,
         aes_state_regs_2_mix_columns_1_n192,
         aes_state_regs_2_mix_columns_1_n191,
         aes_state_regs_2_mix_columns_1_n190,
         aes_state_regs_2_mix_columns_1_n189,
         aes_state_regs_2_mix_columns_1_n188,
         aes_state_regs_2_mix_columns_1_n187,
         aes_state_regs_2_mix_columns_1_n186,
         aes_state_regs_2_mix_columns_1_n185,
         aes_state_regs_2_mix_columns_1_n184,
         aes_state_regs_2_mix_columns_1_n183,
         aes_state_regs_2_mix_columns_1_n182,
         aes_state_regs_2_mix_columns_1_n181,
         aes_state_regs_2_mix_columns_1_n180,
         aes_state_regs_2_mix_columns_1_n179,
         aes_state_regs_2_mix_columns_1_n178,
         aes_state_regs_2_mix_columns_1_n177,
         aes_state_regs_2_mix_columns_1_n176,
         aes_state_regs_2_mix_columns_1_n175,
         aes_state_regs_2_mix_columns_1_n174,
         aes_state_regs_2_mix_columns_1_n173,
         aes_state_regs_2_mix_columns_1_n172,
         aes_state_regs_2_mix_columns_1_n171,
         aes_state_regs_2_mix_columns_1_n170,
         aes_state_regs_2_mix_columns_1_n169,
         aes_state_regs_2_mix_columns_1_n168,
         aes_state_regs_2_mix_columns_1_n167,
         aes_state_regs_2_mix_columns_1_n166,
         aes_state_regs_2_mix_columns_1_n165,
         aes_state_regs_2_mix_columns_1_n164,
         aes_state_regs_2_mix_columns_1_n163,
         aes_state_regs_2_mix_columns_1_n162,
         aes_state_regs_2_mix_columns_1_n161,
         aes_state_regs_2_mix_columns_1_n160,
         aes_state_regs_2_mix_columns_1_n159, aes_key_regs_1_n4,
         aes_key_regs_1_K02xDP_0_, aes_key_regs_1_K02xDP_1_,
         aes_key_regs_1_K02xDP_2_, aes_key_regs_1_K02xDP_3_,
         aes_key_regs_1_K02xDP_4_, aes_key_regs_1_K02xDP_5_,
         aes_key_regs_1_K02xDP_6_, aes_key_regs_1_K02xDP_7_,
         aes_key_regs_1_K01xDP_0_, aes_key_regs_1_K01xDP_1_,
         aes_key_regs_1_K01xDP_2_, aes_key_regs_1_K01xDP_3_,
         aes_key_regs_1_K01xDP_4_, aes_key_regs_1_K01xDP_5_,
         aes_key_regs_1_K01xDP_6_, aes_key_regs_1_K01xDP_7_,
         aes_state_regs_1_n202, aes_state_regs_1_n201, aes_state_regs_1_n200,
         aes_state_regs_1_n199, aes_state_regs_1_n198, aes_state_regs_1_n197,
         aes_state_regs_1_n196, aes_state_regs_1_n195, aes_state_regs_1_n194,
         aes_state_regs_1_n193, aes_state_regs_1_n192, aes_state_regs_1_n191,
         aes_state_regs_1_n190, aes_state_regs_1_n189, aes_state_regs_1_n188,
         aes_state_regs_1_n187, aes_state_regs_1_n186, aes_state_regs_1_n185,
         aes_state_regs_1_n184, aes_state_regs_1_n183, aes_state_regs_1_n182,
         aes_state_regs_1_n180, aes_state_regs_1_n179, aes_state_regs_1_n178,
         aes_state_regs_1_n177, aes_state_regs_1_n176, aes_state_regs_1_n175,
         aes_state_regs_1_n174, aes_state_regs_1_n51, aes_state_regs_1_n50,
         aes_state_regs_1_n49, aes_state_regs_1_n48, aes_state_regs_1_n47,
         aes_state_regs_1_n46, aes_state_regs_1_n45, aes_state_regs_1_n44,
         aes_state_regs_1_n43, aes_state_regs_1_n42, aes_state_regs_1_n41,
         aes_state_regs_1_n40, aes_state_regs_1_n39, aes_state_regs_1_n38,
         aes_state_regs_1_n37, aes_state_regs_1_n36, aes_state_regs_1_n35,
         aes_state_regs_1_n34, aes_state_regs_1_n33, aes_state_regs_1_n32,
         aes_state_regs_1_n31, aes_state_regs_1_n30, aes_state_regs_1_n29,
         aes_state_regs_1_n28, aes_state_regs_1_n173, aes_state_regs_1_n172,
         aes_state_regs_1_n171, aes_state_regs_1_n170, aes_state_regs_1_n169,
         aes_state_regs_1_n168, aes_state_regs_1_n167, aes_state_regs_1_n166,
         aes_state_regs_1_n165, aes_state_regs_1_n164, aes_state_regs_1_n163,
         aes_state_regs_1_n162, aes_state_regs_1_n161, aes_state_regs_1_n160,
         aes_state_regs_1_n159, aes_state_regs_1_n158, aes_state_regs_1_n157,
         aes_state_regs_1_n156, aes_state_regs_1_n155, aes_state_regs_1_n154,
         aes_state_regs_1_n153, aes_state_regs_1_n152, aes_state_regs_1_n151,
         aes_state_regs_1_n150, aes_state_regs_1_n149, aes_state_regs_1_n148,
         aes_state_regs_1_n147, aes_state_regs_1_n146, aes_state_regs_1_n145,
         aes_state_regs_1_n144, aes_state_regs_1_n143, aes_state_regs_1_n142,
         aes_state_regs_1_n141, aes_state_regs_1_n140, aes_state_regs_1_n139,
         aes_state_regs_1_n138, aes_state_regs_1_n137, aes_state_regs_1_n136,
         aes_state_regs_1_n127, aes_state_regs_1_n126, aes_state_regs_1_n125,
         aes_state_regs_1_n124, aes_state_regs_1_n123, aes_state_regs_1_n122,
         aes_state_regs_1_n121, aes_state_regs_1_n109,
         aes_state_regs_1_S03xDP_0_, aes_state_regs_1_S02xDP_0_,
         aes_state_regs_1_S02xDP_1_, aes_state_regs_1_S02xDP_2_,
         aes_state_regs_1_S02xDP_3_, aes_state_regs_1_S02xDP_4_,
         aes_state_regs_1_S02xDP_5_, aes_state_regs_1_S02xDP_6_,
         aes_state_regs_1_S02xDP_7_, aes_state_regs_1_S31xDP_0_,
         aes_state_regs_1_S30xDP_0_, aes_state_regs_1_S30xDP_1_,
         aes_state_regs_1_S30xDP_2_, aes_state_regs_1_S30xDP_3_,
         aes_state_regs_1_S30xDP_4_, aes_state_regs_1_S30xDP_5_,
         aes_state_regs_1_S30xDP_6_, aes_state_regs_1_S30xDP_7_,
         aes_state_regs_1_S20xDP_0_, aes_state_regs_1_S20xDP_1_,
         aes_state_regs_1_S20xDP_2_, aes_state_regs_1_S20xDP_3_,
         aes_state_regs_1_S20xDP_4_, aes_state_regs_1_S20xDP_5_,
         aes_state_regs_1_S20xDP_6_, aes_state_regs_1_S20xDP_7_,
         aes_state_regs_1_S23xDP_0_, aes_state_regs_1_S23xDP_1_,
         aes_state_regs_1_S23xDP_2_, aes_state_regs_1_S23xDP_3_,
         aes_state_regs_1_S23xDP_4_, aes_state_regs_1_S23xDP_5_,
         aes_state_regs_1_S23xDP_6_, aes_state_regs_1_S23xDP_7_,
         aes_state_regs_1_S22xDP_0_, aes_state_regs_1_S10xDP_0_,
         aes_state_regs_1_S10xDP_1_, aes_state_regs_1_S10xDP_2_,
         aes_state_regs_1_S10xDP_3_, aes_state_regs_1_S10xDP_4_,
         aes_state_regs_1_S10xDP_5_, aes_state_regs_1_S10xDP_6_,
         aes_state_regs_1_S10xDP_7_, aes_state_regs_1_S01xDO_0_,
         aes_state_regs_1_S01xDO_1_, aes_state_regs_1_S01xDO_2_,
         aes_state_regs_1_S01xDO_3_, aes_state_regs_1_S01xDO_4_,
         aes_state_regs_1_S01xDO_5_, aes_state_regs_1_S01xDO_6_,
         aes_state_regs_1_S01xDO_7_, aes_state_regs_1_mix_columns_1_n245,
         aes_state_regs_1_mix_columns_1_n244,
         aes_state_regs_1_mix_columns_1_n243,
         aes_state_regs_1_mix_columns_1_n242,
         aes_state_regs_1_mix_columns_1_n241,
         aes_state_regs_1_mix_columns_1_n240,
         aes_state_regs_1_mix_columns_1_n239,
         aes_state_regs_1_mix_columns_1_n238,
         aes_state_regs_1_mix_columns_1_n237,
         aes_state_regs_1_mix_columns_1_n236,
         aes_state_regs_1_mix_columns_1_n235,
         aes_state_regs_1_mix_columns_1_n234,
         aes_state_regs_1_mix_columns_1_n233,
         aes_state_regs_1_mix_columns_1_n232,
         aes_state_regs_1_mix_columns_1_n231,
         aes_state_regs_1_mix_columns_1_n230,
         aes_state_regs_1_mix_columns_1_n229,
         aes_state_regs_1_mix_columns_1_n228,
         aes_state_regs_1_mix_columns_1_n227,
         aes_state_regs_1_mix_columns_1_n226,
         aes_state_regs_1_mix_columns_1_n225,
         aes_state_regs_1_mix_columns_1_n224,
         aes_state_regs_1_mix_columns_1_n223,
         aes_state_regs_1_mix_columns_1_n222,
         aes_state_regs_1_mix_columns_1_n221,
         aes_state_regs_1_mix_columns_1_n220,
         aes_state_regs_1_mix_columns_1_n219,
         aes_state_regs_1_mix_columns_1_n218,
         aes_state_regs_1_mix_columns_1_n217,
         aes_state_regs_1_mix_columns_1_n216,
         aes_state_regs_1_mix_columns_1_n215,
         aes_state_regs_1_mix_columns_1_n214,
         aes_state_regs_1_mix_columns_1_n213,
         aes_state_regs_1_mix_columns_1_n212,
         aes_state_regs_1_mix_columns_1_n211,
         aes_state_regs_1_mix_columns_1_n210,
         aes_state_regs_1_mix_columns_1_n209,
         aes_state_regs_1_mix_columns_1_n208,
         aes_state_regs_1_mix_columns_1_n207,
         aes_state_regs_1_mix_columns_1_n206,
         aes_state_regs_1_mix_columns_1_n205,
         aes_state_regs_1_mix_columns_1_n204,
         aes_state_regs_1_mix_columns_1_n203,
         aes_state_regs_1_mix_columns_1_n202,
         aes_state_regs_1_mix_columns_1_n201,
         aes_state_regs_1_mix_columns_1_n200,
         aes_state_regs_1_mix_columns_1_n199,
         aes_state_regs_1_mix_columns_1_n198,
         aes_state_regs_1_mix_columns_1_n197,
         aes_state_regs_1_mix_columns_1_n196,
         aes_state_regs_1_mix_columns_1_n195,
         aes_state_regs_1_mix_columns_1_n194,
         aes_state_regs_1_mix_columns_1_n193,
         aes_state_regs_1_mix_columns_1_n192,
         aes_state_regs_1_mix_columns_1_n191,
         aes_state_regs_1_mix_columns_1_n190,
         aes_state_regs_1_mix_columns_1_n189,
         aes_state_regs_1_mix_columns_1_n188,
         aes_state_regs_1_mix_columns_1_n187,
         aes_state_regs_1_mix_columns_1_n186,
         aes_state_regs_1_mix_columns_1_n185,
         aes_state_regs_1_mix_columns_1_n184,
         aes_state_regs_1_mix_columns_1_n183,
         aes_state_regs_1_mix_columns_1_n182,
         aes_state_regs_1_mix_columns_1_n181,
         aes_state_regs_1_mix_columns_1_n180,
         aes_state_regs_1_mix_columns_1_n179,
         aes_state_regs_1_mix_columns_1_n178,
         aes_state_regs_1_mix_columns_1_n177,
         aes_state_regs_1_mix_columns_1_n176,
         aes_state_regs_1_mix_columns_1_n175,
         aes_state_regs_1_mix_columns_1_n174,
         aes_state_regs_1_mix_columns_1_n173,
         aes_state_regs_1_mix_columns_1_n172,
         aes_state_regs_1_mix_columns_1_n171,
         aes_state_regs_1_mix_columns_1_n170,
         aes_state_regs_1_mix_columns_1_n169,
         aes_state_regs_1_mix_columns_1_n168,
         aes_state_regs_1_mix_columns_1_n167,
         aes_state_regs_1_mix_columns_1_n166,
         aes_state_regs_1_mix_columns_1_n165,
         aes_state_regs_1_mix_columns_1_n164,
         aes_state_regs_1_mix_columns_1_n163,
         aes_state_regs_1_mix_columns_1_n162,
         aes_state_regs_1_mix_columns_1_n161,
         aes_state_regs_1_mix_columns_1_n160,
         aes_state_regs_1_mix_columns_1_n159, aes_key_regs_0_n4,
         aes_key_regs_0_K02xDP_0_, aes_key_regs_0_K02xDP_1_,
         aes_key_regs_0_K02xDP_2_, aes_key_regs_0_K02xDP_3_,
         aes_key_regs_0_K02xDP_4_, aes_key_regs_0_K02xDP_5_,
         aes_key_regs_0_K02xDP_6_, aes_key_regs_0_K02xDP_7_,
         aes_key_regs_0_K01xDP_0_, aes_key_regs_0_K01xDP_1_,
         aes_key_regs_0_K01xDP_2_, aes_key_regs_0_K01xDP_3_,
         aes_key_regs_0_K01xDP_4_, aes_key_regs_0_K01xDP_5_,
         aes_key_regs_0_K01xDP_6_, aes_key_regs_0_K01xDP_7_,
         aes_state_regs_0_n203, aes_state_regs_0_n202, aes_state_regs_0_n201,
         aes_state_regs_0_n200, aes_state_regs_0_n199, aes_state_regs_0_n198,
         aes_state_regs_0_n197, aes_state_regs_0_n196, aes_state_regs_0_n195,
         aes_state_regs_0_n194, aes_state_regs_0_n193, aes_state_regs_0_n192,
         aes_state_regs_0_n191, aes_state_regs_0_n190, aes_state_regs_0_n189,
         aes_state_regs_0_n188, aes_state_regs_0_n187, aes_state_regs_0_n186,
         aes_state_regs_0_n185, aes_state_regs_0_n184, aes_state_regs_0_n183,
         aes_state_regs_0_n182, aes_state_regs_0_n181, aes_state_regs_0_n180,
         aes_state_regs_0_n179, aes_state_regs_0_n178, aes_state_regs_0_n176,
         aes_state_regs_0_n175, aes_state_regs_0_n174, aes_state_regs_0_n51,
         aes_state_regs_0_n50, aes_state_regs_0_n49, aes_state_regs_0_n48,
         aes_state_regs_0_n47, aes_state_regs_0_n46, aes_state_regs_0_n45,
         aes_state_regs_0_n44, aes_state_regs_0_n43, aes_state_regs_0_n42,
         aes_state_regs_0_n41, aes_state_regs_0_n40, aes_state_regs_0_n39,
         aes_state_regs_0_n38, aes_state_regs_0_n37, aes_state_regs_0_n36,
         aes_state_regs_0_n35, aes_state_regs_0_n34, aes_state_regs_0_n33,
         aes_state_regs_0_n32, aes_state_regs_0_n31, aes_state_regs_0_n30,
         aes_state_regs_0_n29, aes_state_regs_0_n28, aes_state_regs_0_n173,
         aes_state_regs_0_n172, aes_state_regs_0_n171, aes_state_regs_0_n170,
         aes_state_regs_0_n169, aes_state_regs_0_n168, aes_state_regs_0_n167,
         aes_state_regs_0_n166, aes_state_regs_0_n165, aes_state_regs_0_n164,
         aes_state_regs_0_n163, aes_state_regs_0_n162, aes_state_regs_0_n161,
         aes_state_regs_0_n160, aes_state_regs_0_n159, aes_state_regs_0_n158,
         aes_state_regs_0_n157, aes_state_regs_0_n156, aes_state_regs_0_n155,
         aes_state_regs_0_n154, aes_state_regs_0_n153, aes_state_regs_0_n152,
         aes_state_regs_0_n151, aes_state_regs_0_n150, aes_state_regs_0_n149,
         aes_state_regs_0_n148, aes_state_regs_0_n147, aes_state_regs_0_n146,
         aes_state_regs_0_n145, aes_state_regs_0_n144, aes_state_regs_0_n143,
         aes_state_regs_0_n142, aes_state_regs_0_n141, aes_state_regs_0_n140,
         aes_state_regs_0_n139, aes_state_regs_0_n138, aes_state_regs_0_n137,
         aes_state_regs_0_n136, aes_state_regs_0_n127, aes_state_regs_0_n126,
         aes_state_regs_0_n125, aes_state_regs_0_n124, aes_state_regs_0_n123,
         aes_state_regs_0_n122, aes_state_regs_0_n121, aes_state_regs_0_n109,
         aes_state_regs_0_S03xDP_0_, aes_state_regs_0_S02xDP_0_,
         aes_state_regs_0_S02xDP_1_, aes_state_regs_0_S02xDP_2_,
         aes_state_regs_0_S02xDP_3_, aes_state_regs_0_S02xDP_4_,
         aes_state_regs_0_S02xDP_5_, aes_state_regs_0_S02xDP_6_,
         aes_state_regs_0_S02xDP_7_, aes_state_regs_0_S31xDP_0_,
         aes_state_regs_0_S30xDP_0_, aes_state_regs_0_S30xDP_1_,
         aes_state_regs_0_S30xDP_2_, aes_state_regs_0_S30xDP_3_,
         aes_state_regs_0_S30xDP_4_, aes_state_regs_0_S30xDP_5_,
         aes_state_regs_0_S30xDP_6_, aes_state_regs_0_S30xDP_7_,
         aes_state_regs_0_S20xDP_0_, aes_state_regs_0_S20xDP_1_,
         aes_state_regs_0_S20xDP_2_, aes_state_regs_0_S20xDP_3_,
         aes_state_regs_0_S20xDP_4_, aes_state_regs_0_S20xDP_5_,
         aes_state_regs_0_S20xDP_6_, aes_state_regs_0_S20xDP_7_,
         aes_state_regs_0_S23xDP_0_, aes_state_regs_0_S23xDP_1_,
         aes_state_regs_0_S23xDP_2_, aes_state_regs_0_S23xDP_3_,
         aes_state_regs_0_S23xDP_4_, aes_state_regs_0_S23xDP_5_,
         aes_state_regs_0_S23xDP_6_, aes_state_regs_0_S23xDP_7_,
         aes_state_regs_0_S22xDP_0_, aes_state_regs_0_S10xDP_0_,
         aes_state_regs_0_S10xDP_1_, aes_state_regs_0_S10xDP_2_,
         aes_state_regs_0_S10xDP_3_, aes_state_regs_0_S10xDP_4_,
         aes_state_regs_0_S10xDP_5_, aes_state_regs_0_S10xDP_6_,
         aes_state_regs_0_S10xDP_7_, aes_state_regs_0_S01xDO_0_,
         aes_state_regs_0_S01xDO_1_, aes_state_regs_0_S01xDO_2_,
         aes_state_regs_0_S01xDO_3_, aes_state_regs_0_S01xDO_4_,
         aes_state_regs_0_S01xDO_5_, aes_state_regs_0_S01xDO_6_,
         aes_state_regs_0_S01xDO_7_, aes_state_regs_0_mix_columns_1_n245,
         aes_state_regs_0_mix_columns_1_n244,
         aes_state_regs_0_mix_columns_1_n243,
         aes_state_regs_0_mix_columns_1_n242,
         aes_state_regs_0_mix_columns_1_n241,
         aes_state_regs_0_mix_columns_1_n240,
         aes_state_regs_0_mix_columns_1_n239,
         aes_state_regs_0_mix_columns_1_n238,
         aes_state_regs_0_mix_columns_1_n237,
         aes_state_regs_0_mix_columns_1_n236,
         aes_state_regs_0_mix_columns_1_n235,
         aes_state_regs_0_mix_columns_1_n234,
         aes_state_regs_0_mix_columns_1_n233,
         aes_state_regs_0_mix_columns_1_n232,
         aes_state_regs_0_mix_columns_1_n231,
         aes_state_regs_0_mix_columns_1_n230,
         aes_state_regs_0_mix_columns_1_n229,
         aes_state_regs_0_mix_columns_1_n228,
         aes_state_regs_0_mix_columns_1_n227,
         aes_state_regs_0_mix_columns_1_n226,
         aes_state_regs_0_mix_columns_1_n225,
         aes_state_regs_0_mix_columns_1_n224,
         aes_state_regs_0_mix_columns_1_n223,
         aes_state_regs_0_mix_columns_1_n222,
         aes_state_regs_0_mix_columns_1_n221,
         aes_state_regs_0_mix_columns_1_n220,
         aes_state_regs_0_mix_columns_1_n219,
         aes_state_regs_0_mix_columns_1_n218,
         aes_state_regs_0_mix_columns_1_n217,
         aes_state_regs_0_mix_columns_1_n216,
         aes_state_regs_0_mix_columns_1_n215,
         aes_state_regs_0_mix_columns_1_n214,
         aes_state_regs_0_mix_columns_1_n213,
         aes_state_regs_0_mix_columns_1_n212,
         aes_state_regs_0_mix_columns_1_n211,
         aes_state_regs_0_mix_columns_1_n210,
         aes_state_regs_0_mix_columns_1_n209,
         aes_state_regs_0_mix_columns_1_n208,
         aes_state_regs_0_mix_columns_1_n207,
         aes_state_regs_0_mix_columns_1_n206,
         aes_state_regs_0_mix_columns_1_n205,
         aes_state_regs_0_mix_columns_1_n204,
         aes_state_regs_0_mix_columns_1_n203,
         aes_state_regs_0_mix_columns_1_n202,
         aes_state_regs_0_mix_columns_1_n201,
         aes_state_regs_0_mix_columns_1_n200,
         aes_state_regs_0_mix_columns_1_n199,
         aes_state_regs_0_mix_columns_1_n198,
         aes_state_regs_0_mix_columns_1_n197,
         aes_state_regs_0_mix_columns_1_n196,
         aes_state_regs_0_mix_columns_1_n195,
         aes_state_regs_0_mix_columns_1_n194,
         aes_state_regs_0_mix_columns_1_n193,
         aes_state_regs_0_mix_columns_1_n192,
         aes_state_regs_0_mix_columns_1_n191,
         aes_state_regs_0_mix_columns_1_n190,
         aes_state_regs_0_mix_columns_1_n189,
         aes_state_regs_0_mix_columns_1_n188,
         aes_state_regs_0_mix_columns_1_n187,
         aes_state_regs_0_mix_columns_1_n186,
         aes_state_regs_0_mix_columns_1_n185,
         aes_state_regs_0_mix_columns_1_n184,
         aes_state_regs_0_mix_columns_1_n183,
         aes_state_regs_0_mix_columns_1_n182,
         aes_state_regs_0_mix_columns_1_n181,
         aes_state_regs_0_mix_columns_1_n180,
         aes_state_regs_0_mix_columns_1_n179,
         aes_state_regs_0_mix_columns_1_n178,
         aes_state_regs_0_mix_columns_1_n177,
         aes_state_regs_0_mix_columns_1_n176,
         aes_state_regs_0_mix_columns_1_n175,
         aes_state_regs_0_mix_columns_1_n174,
         aes_state_regs_0_mix_columns_1_n173,
         aes_state_regs_0_mix_columns_1_n172,
         aes_state_regs_0_mix_columns_1_n171,
         aes_state_regs_0_mix_columns_1_n170,
         aes_state_regs_0_mix_columns_1_n169,
         aes_state_regs_0_mix_columns_1_n168,
         aes_state_regs_0_mix_columns_1_n167,
         aes_state_regs_0_mix_columns_1_n166,
         aes_state_regs_0_mix_columns_1_n165,
         aes_state_regs_0_mix_columns_1_n164,
         aes_state_regs_0_mix_columns_1_n163,
         aes_state_regs_0_mix_columns_1_n162,
         aes_state_regs_0_mix_columns_1_n161,
         aes_state_regs_0_mix_columns_1_n160,
         aes_state_regs_0_mix_columns_1_n159;
  wire   [23:0] KeyToSboxOutxD;
  wire   [23:0] KeyInxD;
  wire   [23:0] StateOutxD;
  wire   [23:0] StateInxD;
  wire   [23:0] KeyOutxD;
  wire   [23:0] K03xD;
  wire   [7:0] RCONxD;
  wire   [23:0] SBOX_Qreg6;
  wire   [23:0] SBOX_Qreg5;
  wire   [23:0] SBOX_Qoutput;
  wire   [35:0] SBOX_FF4_out;
  wire   [5:0] SBOX_pl_L;
  wire   [5:0] SBOX_p_L;
  wire   [5:0] SBOX_ph_L;
  wire   [5:0] SBOX_pl_H;
  wire   [5:0] SBOX_p_H;
  wire   [5:0] SBOX_ph_H;
  wire   [35:0] SBOX_FF3_out;
  wire   [11:0] SBOX_muld;
  wire   [11:0] SBOX_Zl_f3;
  wire   [11:0] SBOX_Zh_f3;
  wire   [23:0] SBOX_FF2_out;
  wire   [5:0] SBOX_gamma0;
  wire   [5:0] SBOX_ab;
  wire   [5:0] SBOX_sA2N;
  wire   [5:0] SBOX_gamma1;
  wire   [11:0] SBOX_Zl_f2;
  wire   [11:0] SBOX_Zh_f2;
  wire   [29:0] SBOX_FF1_out;
  wire   [5:0] SBOX_pl;
  wire   [5:0] SBOX_p;
  wire   [5:0] SBOX_ph;
  wire   [11:0] SBOX_ab2;
  wire   [11:0] SBOX_Zh_f1;
  wire   [11:1] SBOX_Inst_f1_sZ;
  wire   [5:0] SBOX_Inst_f1_phpplmul_Orig_pl;
  wire   [5:0] SBOX_Inst_f1_phpplmul_Orig_p;
  wire   [5:0] SBOX_Inst_f1_phpplmul_Orig_ph;
  wire   [5:0] SBOX_Inst_f1_phpplmul_sB;
  wire   [5:0] SBOX_Inst_f1_phpplmul_sA;
  wire   [11:0] SBOX_Inst_f2_abin;
  wire   [5:0] SBOX_Inst_f2_dinv_1_Orig_sA2N;
  wire   [5:1] SBOX_Inst_f2_dinv_1_sA2;
  wire   [5:0] SBOX_Inst_f2_dinv_1_Orig_ab;
  wire   [5:0] SBOX_Inst_f3_dinv_2_ph;
  wire   [5:0] SBOX_Inst_f3_dinv_2_pl;
  wire   [5:0] SBOX_Inst_f4_multd_L_Orig_pl;
  wire   [5:0] SBOX_Inst_f4_multd_L_Orig_p;
  wire   [5:0] SBOX_Inst_f4_multd_L_Orig_ph;
  wire   [5:0] SBOX_Inst_f4_multd_L_sB;
  wire   [5:0] SBOX_Inst_f4_multd_L_sA;
  wire   [5:0] SBOX_Inst_f4_multd_H_Orig_pl;
  wire   [5:0] SBOX_Inst_f4_multd_H_Orig_p;
  wire   [5:0] SBOX_Inst_f4_multd_H_Orig_ph;
  wire   [5:0] SBOX_Inst_f4_multd_H_sB;
  wire   [5:0] SBOX_Inst_f4_multd_H_sA;
  wire   [11:0] SBOX_Inst_f5_pl;
  wire   [11:0] SBOX_Inst_f5_ph;
  wire   [7:0] aes_key_regs_2_K23xDN;
  wire   [7:0] aes_key_regs_2_K22xDN;
  wire   [7:0] aes_key_regs_2_K21xDN;
  wire   [7:0] aes_key_regs_2_K20xDN;
  wire   [7:0] aes_key_regs_2_K13xDN;
  wire   [7:0] aes_key_regs_2_K12xDN;
  wire   [7:0] aes_key_regs_2_K11xDN;
  wire   [7:0] aes_key_regs_2_K10xDN;
  wire   [7:0] aes_key_regs_2_K02xDN;
  wire   [7:0] aes_key_regs_2_K01xDN;
  wire   [7:0] aes_key_regs_2_K00xDN;
  wire   [7:0] aes_state_regs_2_MixColumnsS3xD;
  wire   [7:0] aes_state_regs_2_MixColumnsS2xD;
  wire   [7:0] aes_state_regs_2_MixColumnsS1xD;
  wire   [7:0] aes_state_regs_2_MixColumnsS0xD;
  wire   [7:0] aes_state_regs_2_S20xDN;
  wire   [7:1] aes_state_regs_2_S21xDP;
  wire   [7:0] aes_state_regs_2_S10xDN;
  wire   [7:0] aes_state_regs_2_S03xDN;
  wire   [7:0] aes_state_regs_2_S02xDN;
  wire   [7:0] aes_state_regs_2_S01xDN;
  wire   [7:0] aes_state_regs_2_S00xDP;
  wire   [7:0] aes_key_regs_1_K23xDN;
  wire   [7:0] aes_key_regs_1_K22xDN;
  wire   [7:0] aes_key_regs_1_K21xDN;
  wire   [7:0] aes_key_regs_1_K20xDN;
  wire   [7:0] aes_key_regs_1_K13xDN;
  wire   [7:0] aes_key_regs_1_K12xDN;
  wire   [7:0] aes_key_regs_1_K11xDN;
  wire   [7:0] aes_key_regs_1_K10xDN;
  wire   [7:0] aes_key_regs_1_K02xDN;
  wire   [7:0] aes_key_regs_1_K01xDN;
  wire   [7:0] aes_key_regs_1_K00xDN;
  wire   [7:0] aes_state_regs_1_MixColumnsS3xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS2xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS1xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS0xD;
  wire   [7:0] aes_state_regs_1_S20xDN;
  wire   [7:1] aes_state_regs_1_S21xDP;
  wire   [7:0] aes_state_regs_1_S10xDN;
  wire   [7:0] aes_state_regs_1_S03xDN;
  wire   [7:0] aes_state_regs_1_S02xDN;
  wire   [7:0] aes_state_regs_1_S01xDN;
  wire   [7:0] aes_state_regs_1_S00xDP;
  wire   [7:0] aes_key_regs_0_K23xDN;
  wire   [7:0] aes_key_regs_0_K22xDN;
  wire   [7:0] aes_key_regs_0_K21xDN;
  wire   [7:0] aes_key_regs_0_K20xDN;
  wire   [7:0] aes_key_regs_0_K13xDN;
  wire   [7:0] aes_key_regs_0_K12xDN;
  wire   [7:0] aes_key_regs_0_K11xDN;
  wire   [7:0] aes_key_regs_0_K10xDN;
  wire   [7:0] aes_key_regs_0_K02xDN;
  wire   [7:0] aes_key_regs_0_K01xDN;
  wire   [7:0] aes_key_regs_0_K00xDN;
  wire   [7:0] aes_state_regs_0_MixColumnsS3xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS2xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS1xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS0xD;
  wire   [7:0] aes_state_regs_0_S20xDN;
  wire   [7:1] aes_state_regs_0_S21xDP;
  wire   [7:0] aes_state_regs_0_S10xDN;
  wire   [7:0] aes_state_regs_0_S03xDN;
  wire   [7:0] aes_state_regs_0_S02xDN;
  wire   [7:0] aes_state_regs_0_S01xDN;
  wire   [7:0] aes_state_regs_0_S00xDP;

  DFFS_X1 disableKeyRegsxSP_reg ( .D(disableKeyRegsxS), .CK(ClkxCI), .SN(
        RstxBI), .Q(n330), .QN() );
  NAND2_X1 U424 ( .A1(n454), .A2(n464), .ZN(n498) );
  INV_X1 U425 ( .A(n497), .ZN(n458) );
  OAI22_X1 U426 ( .A1(StateOutxD[16]), .A2(n458), .B1(PTxDI[16]), .B2(n460), 
        .ZN(n492) );
  INV_X1 U427 ( .A(n497), .ZN(n459) );
  INV_X1 U428 ( .A(n461), .ZN(n460) );
  INV_X1 U429 ( .A(n459), .ZN(n457) );
  INV_X2 U430 ( .A(n498), .ZN(n461) );
  NOR2_X1 U431 ( .A1(StateKEYSCHEDULExS), .A2(n453), .ZN(n464) );
  OR2_X1 U432 ( .A1(n454), .A2(StateKEYADDITION1o3xS), .ZN(n455) );
  NOR2_X2 U433 ( .A1(n454), .A2(n463), .ZN(n495) );
  INV_X1 U434 ( .A(StateKEYADDITION1o3xS), .ZN(n463) );
  INV_X2 U435 ( .A(n455), .ZN(n456) );
  INV_X2 U436 ( .A(n495), .ZN(n496) );
  AOI22_X1 U437 ( .A1(KeyToSboxOutxD[0]), .A2(n170), .B1(n465), .B2(KeyInxD[0]), .ZN(n466) );
  AOI22_X1 U438 ( .A1(n457), .A2(StateOutxD[0]), .B1(n461), .B2(PTxDI[0]), 
        .ZN(n467) );
  OAI21_X1 U439 ( .B1(n470), .B2(KeyInxD[1]), .A(n469), .ZN(CxDO[1]) );
  AOI22_X1 U440 ( .A1(KeyToSboxOutxD[1]), .A2(n170), .B1(n468), .B2(KeyInxD[1]), .ZN(n469) );
  OAI21_X1 U441 ( .B1(n473), .B2(KeyInxD[3]), .A(n472), .ZN(CxDO[3]) );
  AOI22_X1 U442 ( .A1(KeyToSboxOutxD[3]), .A2(n170), .B1(n471), .B2(KeyInxD[3]), .ZN(n472) );
  AOI22_X1 U443 ( .A1(n457), .A2(StateOutxD[3]), .B1(n461), .B2(PTxDI[3]), 
        .ZN(n473) );
  OAI22_X1 U444 ( .A1(StateOutxD[3]), .A2(n458), .B1(PTxDI[3]), .B2(n498), 
        .ZN(n471) );
  OAI21_X1 U445 ( .B1(n476), .B2(KeyInxD[4]), .A(n475), .ZN(CxDO[4]) );
  AOI22_X1 U446 ( .A1(KeyToSboxOutxD[4]), .A2(n170), .B1(n474), .B2(KeyInxD[4]), .ZN(n475) );
  AOI22_X1 U447 ( .A1(n457), .A2(StateOutxD[4]), .B1(n461), .B2(PTxDI[4]), 
        .ZN(n476) );
  OAI22_X1 U448 ( .A1(StateOutxD[4]), .A2(n458), .B1(PTxDI[4]), .B2(n498), 
        .ZN(n474) );
  OAI21_X1 U449 ( .B1(n479), .B2(KeyInxD[5]), .A(n478), .ZN(CxDO[5]) );
  AOI22_X1 U450 ( .A1(KeyToSboxOutxD[5]), .A2(n170), .B1(n477), .B2(KeyInxD[5]), .ZN(n478) );
  OAI22_X1 U451 ( .A1(StateOutxD[5]), .A2(n458), .B1(PTxDI[5]), .B2(n498), 
        .ZN(n477) );
  AOI22_X1 U452 ( .A1(KeyToSboxOutxD[8]), .A2(n170), .B1(n480), .B2(KeyInxD[8]), .ZN(n481) );
  AOI22_X1 U453 ( .A1(n457), .A2(StateOutxD[8]), .B1(n461), .B2(PTxDI[8]), 
        .ZN(n482) );
  OAI21_X1 U454 ( .B1(n485), .B2(KeyInxD[9]), .A(n484), .ZN(CxDO[9]) );
  AOI22_X1 U455 ( .A1(KeyToSboxOutxD[9]), .A2(n170), .B1(n483), .B2(KeyInxD[9]), .ZN(n484) );
  OAI22_X1 U456 ( .A1(StateOutxD[9]), .A2(n458), .B1(PTxDI[9]), .B2(n498), 
        .ZN(n483) );
  OAI21_X1 U457 ( .B1(n488), .B2(KeyInxD[11]), .A(n487), .ZN(CxDO[11]) );
  AOI22_X1 U458 ( .A1(KeyToSboxOutxD[11]), .A2(n170), .B1(n486), .B2(
        KeyInxD[11]), .ZN(n487) );
  OAI22_X1 U459 ( .A1(StateOutxD[11]), .A2(n458), .B1(PTxDI[11]), .B2(n498), 
        .ZN(n486) );
  OAI21_X1 U460 ( .B1(n491), .B2(KeyInxD[13]), .A(n490), .ZN(CxDO[13]) );
  AOI22_X1 U461 ( .A1(KeyToSboxOutxD[13]), .A2(n170), .B1(n489), .B2(
        KeyInxD[13]), .ZN(n490) );
  AOI22_X1 U462 ( .A1(n457), .A2(StateOutxD[13]), .B1(n461), .B2(PTxDI[13]), 
        .ZN(n491) );
  OAI22_X1 U463 ( .A1(StateOutxD[13]), .A2(n458), .B1(PTxDI[13]), .B2(n460), 
        .ZN(n489) );
  AOI22_X1 U464 ( .A1(KeyToSboxOutxD[16]), .A2(n170), .B1(n492), .B2(
        KeyInxD[16]), .ZN(n493) );
  AOI22_X1 U465 ( .A1(n457), .A2(StateOutxD[16]), .B1(n461), .B2(PTxDI[16]), 
        .ZN(n494) );
  AND2_X1 U466 ( .A1(LastRoundxS), .A2(showRCONxS), .ZN(DonexSO) );
  AOI22_X1 U467 ( .A1(n497), .A2(StateOutxD[2]), .B1(n461), .B2(PTxDI[2]), 
        .ZN(n331) );
  OAI22_X1 U468 ( .A1(n498), .A2(PTxDI[2]), .B1(n458), .B2(StateOutxD[2]), 
        .ZN(n332) );
  AOI22_X1 U469 ( .A1(n170), .A2(KeyToSboxOutxD[2]), .B1(KeyInxD[2]), .B2(n332), .ZN(n333) );
  OAI21_X1 U470 ( .B1(KeyInxD[2]), .B2(n331), .A(n333), .ZN(CxDO[2]) );
  AOI22_X1 U471 ( .A1(n495), .A2(StateInxD[8]), .B1(n456), .B2(K03xD[8]), .ZN(
        n334) );
  OAI22_X1 U472 ( .A1(n455), .A2(K03xD[8]), .B1(n496), .B2(StateInxD[8]), .ZN(
        n335) );
  AOI22_X1 U473 ( .A1(n454), .A2(KxDI[8]), .B1(KeyOutxD[8]), .B2(n335), .ZN(
        n336) );
  OAI21_X1 U474 ( .B1(KeyOutxD[8]), .B2(n334), .A(n336), .ZN(KeyInxD[8]) );
  AOI22_X1 U475 ( .A1(n461), .A2(PTxDI[17]), .B1(n457), .B2(StateOutxD[17]), 
        .ZN(n337) );
  OAI22_X1 U476 ( .A1(n459), .A2(StateOutxD[17]), .B1(n460), .B2(PTxDI[17]), 
        .ZN(n338) );
  AOI22_X1 U477 ( .A1(n170), .A2(KeyToSboxOutxD[17]), .B1(KeyInxD[17]), .B2(
        n338), .ZN(n339) );
  OAI21_X1 U478 ( .B1(KeyInxD[17]), .B2(n337), .A(n339), .ZN(CxDO[17]) );
  AOI22_X1 U479 ( .A1(n495), .A2(StateInxD[9]), .B1(n456), .B2(K03xD[9]), .ZN(
        n340) );
  OAI22_X1 U480 ( .A1(n455), .A2(K03xD[9]), .B1(n496), .B2(StateInxD[9]), .ZN(
        n341) );
  AOI22_X1 U481 ( .A1(n454), .A2(KxDI[9]), .B1(KeyOutxD[9]), .B2(n341), .ZN(
        n342) );
  OAI21_X1 U482 ( .B1(KeyOutxD[9]), .B2(n340), .A(n342), .ZN(KeyInxD[9]) );
  AOI22_X1 U483 ( .A1(n497), .A2(StateOutxD[6]), .B1(n461), .B2(PTxDI[6]), 
        .ZN(n343) );
  OAI22_X1 U484 ( .A1(n498), .A2(PTxDI[6]), .B1(StateOutxD[6]), .B2(n458), 
        .ZN(n344) );
  AOI22_X1 U485 ( .A1(n170), .A2(KeyToSboxOutxD[6]), .B1(KeyInxD[6]), .B2(n344), .ZN(n345) );
  OAI21_X1 U486 ( .B1(KeyInxD[6]), .B2(n343), .A(n345), .ZN(CxDO[6]) );
  AOI22_X1 U487 ( .A1(n495), .A2(StateInxD[10]), .B1(n456), .B2(K03xD[10]), 
        .ZN(n346) );
  OAI22_X1 U488 ( .A1(n455), .A2(K03xD[10]), .B1(n496), .B2(StateInxD[10]), 
        .ZN(n347) );
  AOI22_X1 U489 ( .A1(n454), .A2(KxDI[10]), .B1(KeyOutxD[10]), .B2(n347), .ZN(
        n348) );
  OAI21_X1 U490 ( .B1(KeyOutxD[10]), .B2(n346), .A(n348), .ZN(KeyInxD[10]) );
  AOI22_X1 U491 ( .A1(n457), .A2(StateOutxD[7]), .B1(n461), .B2(PTxDI[7]), 
        .ZN(n349) );
  OAI22_X1 U492 ( .A1(n498), .A2(PTxDI[7]), .B1(n458), .B2(StateOutxD[7]), 
        .ZN(n350) );
  AOI22_X1 U493 ( .A1(n170), .A2(KeyToSboxOutxD[7]), .B1(KeyInxD[7]), .B2(n350), .ZN(n351) );
  OAI21_X1 U494 ( .B1(KeyInxD[7]), .B2(n349), .A(n351), .ZN(CxDO[7]) );
  AOI22_X1 U495 ( .A1(n495), .A2(StateInxD[11]), .B1(n456), .B2(K03xD[11]), 
        .ZN(n352) );
  OAI22_X1 U496 ( .A1(n455), .A2(K03xD[11]), .B1(n496), .B2(StateInxD[11]), 
        .ZN(n353) );
  AOI22_X1 U497 ( .A1(n454), .A2(KxDI[11]), .B1(KeyOutxD[11]), .B2(n353), .ZN(
        n354) );
  OAI21_X1 U498 ( .B1(KeyOutxD[11]), .B2(n352), .A(n354), .ZN(KeyInxD[11]) );
  AOI22_X1 U499 ( .A1(n497), .A2(StateOutxD[10]), .B1(n461), .B2(PTxDI[10]), 
        .ZN(n355) );
  OAI22_X1 U500 ( .A1(n498), .A2(PTxDI[10]), .B1(n458), .B2(StateOutxD[10]), 
        .ZN(n356) );
  AOI22_X1 U501 ( .A1(n170), .A2(KeyToSboxOutxD[10]), .B1(KeyInxD[10]), .B2(
        n356), .ZN(n357) );
  OAI21_X1 U502 ( .B1(KeyInxD[10]), .B2(n355), .A(n357), .ZN(CxDO[10]) );
  AOI22_X1 U503 ( .A1(n495), .A2(StateInxD[12]), .B1(n456), .B2(K03xD[12]), 
        .ZN(n358) );
  OAI22_X1 U504 ( .A1(n455), .A2(K03xD[12]), .B1(n496), .B2(StateInxD[12]), 
        .ZN(n359) );
  AOI22_X1 U505 ( .A1(n454), .A2(KxDI[12]), .B1(KeyOutxD[12]), .B2(n359), .ZN(
        n360) );
  OAI21_X1 U506 ( .B1(KeyOutxD[12]), .B2(n358), .A(n360), .ZN(KeyInxD[12]) );
  AOI22_X1 U507 ( .A1(n461), .A2(PTxDI[14]), .B1(n457), .B2(StateOutxD[14]), 
        .ZN(n361) );
  OAI22_X1 U508 ( .A1(n460), .A2(PTxDI[14]), .B1(n458), .B2(StateOutxD[14]), 
        .ZN(n362) );
  AOI22_X1 U509 ( .A1(n170), .A2(KeyToSboxOutxD[14]), .B1(KeyInxD[14]), .B2(
        n362), .ZN(n363) );
  OAI21_X1 U510 ( .B1(KeyInxD[14]), .B2(n361), .A(n363), .ZN(CxDO[14]) );
  AOI22_X1 U511 ( .A1(n495), .A2(StateInxD[13]), .B1(n456), .B2(K03xD[13]), 
        .ZN(n364) );
  OAI22_X1 U512 ( .A1(n455), .A2(K03xD[13]), .B1(n496), .B2(StateInxD[13]), 
        .ZN(n365) );
  AOI22_X1 U513 ( .A1(n454), .A2(KxDI[13]), .B1(KeyOutxD[13]), .B2(n365), .ZN(
        n366) );
  OAI21_X1 U514 ( .B1(KeyOutxD[13]), .B2(n364), .A(n366), .ZN(KeyInxD[13]) );
  AOI22_X1 U515 ( .A1(n461), .A2(PTxDI[15]), .B1(n457), .B2(StateOutxD[15]), 
        .ZN(n367) );
  OAI22_X1 U516 ( .A1(n460), .A2(PTxDI[15]), .B1(n458), .B2(StateOutxD[15]), 
        .ZN(n368) );
  AOI22_X1 U517 ( .A1(n170), .A2(KeyToSboxOutxD[15]), .B1(KeyInxD[15]), .B2(
        n368), .ZN(n369) );
  OAI21_X1 U518 ( .B1(KeyInxD[15]), .B2(n367), .A(n369), .ZN(CxDO[15]) );
  AOI22_X1 U519 ( .A1(n495), .A2(StateInxD[14]), .B1(n456), .B2(K03xD[14]), 
        .ZN(n370) );
  OAI22_X1 U520 ( .A1(n455), .A2(K03xD[14]), .B1(n496), .B2(StateInxD[14]), 
        .ZN(n371) );
  AOI22_X1 U521 ( .A1(n454), .A2(KxDI[14]), .B1(KeyOutxD[14]), .B2(n371), .ZN(
        n372) );
  OAI21_X1 U522 ( .B1(KeyOutxD[14]), .B2(n370), .A(n372), .ZN(KeyInxD[14]) );
  AOI22_X1 U523 ( .A1(n461), .A2(PTxDI[23]), .B1(n457), .B2(StateOutxD[23]), 
        .ZN(n373) );
  OAI22_X1 U524 ( .A1(n459), .A2(StateOutxD[23]), .B1(n460), .B2(PTxDI[23]), 
        .ZN(n374) );
  AOI22_X1 U525 ( .A1(n170), .A2(KeyToSboxOutxD[23]), .B1(KeyInxD[23]), .B2(
        n374), .ZN(n375) );
  OAI21_X1 U526 ( .B1(KeyInxD[23]), .B2(n373), .A(n375), .ZN(CxDO[23]) );
  AOI22_X1 U527 ( .A1(n495), .A2(StateInxD[15]), .B1(n456), .B2(K03xD[15]), 
        .ZN(n376) );
  OAI22_X1 U528 ( .A1(n455), .A2(K03xD[15]), .B1(n496), .B2(StateInxD[15]), 
        .ZN(n377) );
  AOI22_X1 U529 ( .A1(n454), .A2(KxDI[15]), .B1(KeyOutxD[15]), .B2(n377), .ZN(
        n378) );
  OAI21_X1 U530 ( .B1(KeyOutxD[15]), .B2(n376), .A(n378), .ZN(KeyInxD[15]) );
  AOI22_X1 U531 ( .A1(n461), .A2(PTxDI[12]), .B1(n457), .B2(StateOutxD[12]), 
        .ZN(n379) );
  OAI22_X1 U532 ( .A1(n460), .A2(PTxDI[12]), .B1(n458), .B2(StateOutxD[12]), 
        .ZN(n380) );
  AOI22_X1 U533 ( .A1(n170), .A2(KeyToSboxOutxD[12]), .B1(KeyInxD[12]), .B2(
        n380), .ZN(n381) );
  OAI21_X1 U534 ( .B1(KeyInxD[12]), .B2(n379), .A(n381), .ZN(CxDO[12]) );
  XOR2_X1 U535 ( .A(StateInxD[0]), .B(KeyOutxD[0]), .Z(n382) );
  XNOR2_X1 U536 ( .A(RCONxD[0]), .B(n382), .ZN(n383) );
  XOR2_X1 U537 ( .A(KeyOutxD[0]), .B(K03xD[0]), .Z(n384) );
  AOI22_X1 U538 ( .A1(n456), .A2(n384), .B1(KxDI[0]), .B2(n454), .ZN(n385) );
  OAI21_X1 U539 ( .B1(n496), .B2(n383), .A(n385), .ZN(KeyInxD[0]) );
  AOI22_X1 U540 ( .A1(n495), .A2(StateInxD[16]), .B1(n456), .B2(K03xD[16]), 
        .ZN(n386) );
  OAI22_X1 U541 ( .A1(n455), .A2(K03xD[16]), .B1(n496), .B2(StateInxD[16]), 
        .ZN(n387) );
  AOI22_X1 U542 ( .A1(n454), .A2(KxDI[16]), .B1(KeyOutxD[16]), .B2(n387), .ZN(
        n388) );
  OAI21_X1 U543 ( .B1(KeyOutxD[16]), .B2(n386), .A(n388), .ZN(KeyInxD[16]) );
  AOI22_X1 U544 ( .A1(n461), .A2(PTxDI[21]), .B1(n457), .B2(StateOutxD[21]), 
        .ZN(n389) );
  OAI22_X1 U545 ( .A1(n459), .A2(StateOutxD[21]), .B1(n460), .B2(PTxDI[21]), 
        .ZN(n390) );
  AOI22_X1 U546 ( .A1(n170), .A2(KeyToSboxOutxD[21]), .B1(KeyInxD[21]), .B2(
        n390), .ZN(n391) );
  OAI21_X1 U547 ( .B1(KeyInxD[21]), .B2(n389), .A(n391), .ZN(CxDO[21]) );
  XOR2_X1 U548 ( .A(StateInxD[1]), .B(KeyOutxD[1]), .Z(n392) );
  XNOR2_X1 U549 ( .A(RCONxD[1]), .B(n392), .ZN(n393) );
  XOR2_X1 U550 ( .A(KeyOutxD[1]), .B(K03xD[1]), .Z(n394) );
  AOI22_X1 U551 ( .A1(n454), .A2(KxDI[1]), .B1(n456), .B2(n394), .ZN(n395) );
  OAI21_X1 U552 ( .B1(n496), .B2(n393), .A(n395), .ZN(KeyInxD[1]) );
  AOI22_X1 U553 ( .A1(n495), .A2(StateInxD[17]), .B1(n456), .B2(K03xD[17]), 
        .ZN(n396) );
  OAI22_X1 U554 ( .A1(n455), .A2(K03xD[17]), .B1(n496), .B2(StateInxD[17]), 
        .ZN(n397) );
  AOI22_X1 U555 ( .A1(n454), .A2(KxDI[17]), .B1(KeyOutxD[17]), .B2(n397), .ZN(
        n398) );
  OAI21_X1 U556 ( .B1(KeyOutxD[17]), .B2(n396), .A(n398), .ZN(KeyInxD[17]) );
  AOI22_X1 U557 ( .A1(n461), .A2(PTxDI[20]), .B1(n457), .B2(StateOutxD[20]), 
        .ZN(n399) );
  OAI22_X1 U558 ( .A1(n459), .A2(StateOutxD[20]), .B1(n460), .B2(PTxDI[20]), 
        .ZN(n400) );
  AOI22_X1 U559 ( .A1(n170), .A2(KeyToSboxOutxD[20]), .B1(KeyInxD[20]), .B2(
        n400), .ZN(n401) );
  OAI21_X1 U560 ( .B1(KeyInxD[20]), .B2(n399), .A(n401), .ZN(CxDO[20]) );
  XOR2_X1 U561 ( .A(StateInxD[3]), .B(KeyOutxD[3]), .Z(n402) );
  XNOR2_X1 U562 ( .A(RCONxD[3]), .B(n402), .ZN(n403) );
  XOR2_X1 U563 ( .A(KeyOutxD[3]), .B(K03xD[3]), .Z(n404) );
  AOI22_X1 U564 ( .A1(n454), .A2(KxDI[3]), .B1(n456), .B2(n404), .ZN(n405) );
  OAI21_X1 U565 ( .B1(n496), .B2(n403), .A(n405), .ZN(KeyInxD[3]) );
  AOI22_X1 U566 ( .A1(n495), .A2(StateInxD[18]), .B1(n456), .B2(K03xD[18]), 
        .ZN(n406) );
  OAI22_X1 U567 ( .A1(n455), .A2(K03xD[18]), .B1(n496), .B2(StateInxD[18]), 
        .ZN(n407) );
  AOI22_X1 U568 ( .A1(n454), .A2(KxDI[18]), .B1(KeyOutxD[18]), .B2(n407), .ZN(
        n408) );
  OAI21_X1 U569 ( .B1(KeyOutxD[18]), .B2(n406), .A(n408), .ZN(KeyInxD[18]) );
  AOI22_X1 U570 ( .A1(n461), .A2(PTxDI[22]), .B1(n457), .B2(StateOutxD[22]), 
        .ZN(n409) );
  OAI22_X1 U571 ( .A1(n459), .A2(StateOutxD[22]), .B1(n460), .B2(PTxDI[22]), 
        .ZN(n410) );
  AOI22_X1 U572 ( .A1(n170), .A2(KeyToSboxOutxD[22]), .B1(KeyInxD[22]), .B2(
        n410), .ZN(n411) );
  OAI21_X1 U573 ( .B1(KeyInxD[22]), .B2(n409), .A(n411), .ZN(CxDO[22]) );
  XOR2_X1 U574 ( .A(StateInxD[7]), .B(KeyOutxD[7]), .Z(n412) );
  XNOR2_X1 U575 ( .A(RCONxD[7]), .B(n412), .ZN(n413) );
  XOR2_X1 U576 ( .A(KeyOutxD[7]), .B(K03xD[7]), .Z(n414) );
  AOI22_X1 U577 ( .A1(n454), .A2(KxDI[7]), .B1(n456), .B2(n414), .ZN(n415) );
  OAI21_X1 U578 ( .B1(n496), .B2(n413), .A(n415), .ZN(KeyInxD[7]) );
  AOI22_X1 U579 ( .A1(n495), .A2(StateInxD[19]), .B1(n456), .B2(K03xD[19]), 
        .ZN(n416) );
  OAI22_X1 U580 ( .A1(n455), .A2(K03xD[19]), .B1(n496), .B2(StateInxD[19]), 
        .ZN(n417) );
  AOI22_X1 U581 ( .A1(n454), .A2(KxDI[19]), .B1(KeyOutxD[19]), .B2(n417), .ZN(
        n418) );
  OAI21_X1 U582 ( .B1(KeyOutxD[19]), .B2(n416), .A(n418), .ZN(KeyInxD[19]) );
  AOI22_X1 U583 ( .A1(n461), .A2(PTxDI[19]), .B1(n457), .B2(StateOutxD[19]), 
        .ZN(n419) );
  OAI22_X1 U584 ( .A1(n459), .A2(StateOutxD[19]), .B1(n460), .B2(PTxDI[19]), 
        .ZN(n420) );
  AOI22_X1 U585 ( .A1(n170), .A2(KeyToSboxOutxD[19]), .B1(KeyInxD[19]), .B2(
        n420), .ZN(n421) );
  OAI21_X1 U586 ( .B1(KeyInxD[19]), .B2(n419), .A(n421), .ZN(CxDO[19]) );
  XOR2_X1 U587 ( .A(StateInxD[2]), .B(KeyOutxD[2]), .Z(n422) );
  XNOR2_X1 U588 ( .A(RCONxD[2]), .B(n422), .ZN(n423) );
  XOR2_X1 U589 ( .A(KeyOutxD[2]), .B(K03xD[2]), .Z(n424) );
  AOI22_X1 U590 ( .A1(n454), .A2(KxDI[2]), .B1(n456), .B2(n424), .ZN(n425) );
  OAI21_X1 U591 ( .B1(n496), .B2(n423), .A(n425), .ZN(KeyInxD[2]) );
  AOI22_X1 U592 ( .A1(n495), .A2(StateInxD[20]), .B1(n456), .B2(K03xD[20]), 
        .ZN(n426) );
  OAI22_X1 U593 ( .A1(n455), .A2(K03xD[20]), .B1(n496), .B2(StateInxD[20]), 
        .ZN(n427) );
  AOI22_X1 U594 ( .A1(n454), .A2(KxDI[20]), .B1(KeyOutxD[20]), .B2(n427), .ZN(
        n428) );
  OAI21_X1 U595 ( .B1(KeyOutxD[20]), .B2(n426), .A(n428), .ZN(KeyInxD[20]) );
  AOI22_X1 U596 ( .A1(n461), .A2(PTxDI[18]), .B1(n457), .B2(StateOutxD[18]), 
        .ZN(n429) );
  OAI22_X1 U597 ( .A1(n459), .A2(StateOutxD[18]), .B1(n460), .B2(PTxDI[18]), 
        .ZN(n430) );
  AOI22_X1 U598 ( .A1(n170), .A2(KeyToSboxOutxD[18]), .B1(KeyInxD[18]), .B2(
        n430), .ZN(n431) );
  OAI21_X1 U599 ( .B1(KeyInxD[18]), .B2(n429), .A(n431), .ZN(CxDO[18]) );
  XOR2_X1 U600 ( .A(StateInxD[4]), .B(KeyOutxD[4]), .Z(n432) );
  XNOR2_X1 U601 ( .A(RCONxD[4]), .B(n432), .ZN(n433) );
  XOR2_X1 U602 ( .A(KeyOutxD[4]), .B(K03xD[4]), .Z(n434) );
  AOI22_X1 U603 ( .A1(n454), .A2(KxDI[4]), .B1(n456), .B2(n434), .ZN(n435) );
  OAI21_X1 U604 ( .B1(n496), .B2(n433), .A(n435), .ZN(KeyInxD[4]) );
  AOI22_X1 U605 ( .A1(n495), .A2(StateInxD[21]), .B1(n456), .B2(K03xD[21]), 
        .ZN(n436) );
  OAI22_X1 U606 ( .A1(n455), .A2(K03xD[21]), .B1(n496), .B2(StateInxD[21]), 
        .ZN(n437) );
  AOI22_X1 U607 ( .A1(n454), .A2(KxDI[21]), .B1(KeyOutxD[21]), .B2(n437), .ZN(
        n438) );
  OAI21_X1 U608 ( .B1(KeyOutxD[21]), .B2(n436), .A(n438), .ZN(KeyInxD[21]) );
  XOR2_X1 U609 ( .A(StateInxD[5]), .B(KeyOutxD[5]), .Z(n439) );
  XNOR2_X1 U610 ( .A(RCONxD[5]), .B(n439), .ZN(n440) );
  XOR2_X1 U611 ( .A(KeyOutxD[5]), .B(K03xD[5]), .Z(n441) );
  AOI22_X1 U612 ( .A1(n454), .A2(KxDI[5]), .B1(n456), .B2(n441), .ZN(n442) );
  OAI21_X1 U613 ( .B1(n496), .B2(n440), .A(n442), .ZN(KeyInxD[5]) );
  AOI22_X1 U614 ( .A1(n495), .A2(StateInxD[22]), .B1(n456), .B2(K03xD[22]), 
        .ZN(n443) );
  OAI22_X1 U615 ( .A1(n455), .A2(K03xD[22]), .B1(n496), .B2(StateInxD[22]), 
        .ZN(n444) );
  AOI22_X1 U616 ( .A1(n454), .A2(KxDI[22]), .B1(KeyOutxD[22]), .B2(n444), .ZN(
        n445) );
  OAI21_X1 U617 ( .B1(KeyOutxD[22]), .B2(n443), .A(n445), .ZN(KeyInxD[22]) );
  XOR2_X1 U618 ( .A(StateInxD[6]), .B(KeyOutxD[6]), .Z(n446) );
  XNOR2_X1 U619 ( .A(RCONxD[6]), .B(n446), .ZN(n447) );
  XOR2_X1 U620 ( .A(KeyOutxD[6]), .B(K03xD[6]), .Z(n448) );
  AOI22_X1 U621 ( .A1(n454), .A2(KxDI[6]), .B1(n456), .B2(n448), .ZN(n449) );
  OAI21_X1 U622 ( .B1(n496), .B2(n447), .A(n449), .ZN(KeyInxD[6]) );
  AOI22_X1 U623 ( .A1(n495), .A2(StateInxD[23]), .B1(n456), .B2(K03xD[23]), 
        .ZN(n450) );
  OAI22_X1 U624 ( .A1(n455), .A2(K03xD[23]), .B1(n496), .B2(StateInxD[23]), 
        .ZN(n451) );
  AOI22_X1 U625 ( .A1(n454), .A2(KxDI[23]), .B1(KeyOutxD[23]), .B2(n451), .ZN(
        n452) );
  OAI21_X1 U626 ( .B1(KeyOutxD[23]), .B2(n450), .A(n452), .ZN(KeyInxD[23]) );
  INV_X1 U627 ( .A(ClkxCI), .ZN(n462) );
  INV_X8 U628 ( .A(n464), .ZN(n170) );
  OAI21_X4 U629 ( .B1(n494), .B2(KeyInxD[16]), .A(n493), .ZN(CxDO[16]) );
  OAI21_X4 U630 ( .B1(n467), .B2(KeyInxD[0]), .A(n466), .ZN(CxDO[0]) );
  OAI21_X4 U631 ( .B1(n482), .B2(KeyInxD[8]), .A(n481), .ZN(CxDO[8]) );
  NOR2_X1 U632 ( .A1(n454), .A2(n170), .ZN(n497) );
  NOR2_X1 U633 ( .A1(n330), .A2(n462), .ZN(ClkKeyRegxC) );
  OAI22_X1 U634 ( .A1(StateOutxD[0]), .A2(n458), .B1(PTxDI[0]), .B2(n460), 
        .ZN(n465) );
  AOI22_X1 U635 ( .A1(n497), .A2(StateOutxD[1]), .B1(n461), .B2(PTxDI[1]), 
        .ZN(n470) );
  OAI22_X1 U636 ( .A1(StateOutxD[1]), .A2(n458), .B1(PTxDI[1]), .B2(n498), 
        .ZN(n468) );
  AOI22_X1 U637 ( .A1(n497), .A2(StateOutxD[5]), .B1(n461), .B2(PTxDI[5]), 
        .ZN(n479) );
  OAI22_X1 U638 ( .A1(StateOutxD[8]), .A2(n458), .B1(PTxDI[8]), .B2(n498), 
        .ZN(n480) );
  AOI22_X1 U639 ( .A1(n497), .A2(StateOutxD[9]), .B1(n461), .B2(PTxDI[9]), 
        .ZN(n485) );
  AOI22_X1 U640 ( .A1(n497), .A2(StateOutxD[11]), .B1(n461), .B2(PTxDI[11]), 
        .ZN(n488) );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U31 ( .A1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n7), .ZN(aes_ctrl_lsfr_23_cycles_1_n17)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U30 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n9), .ZN(aes_ctrl_lsfr_23_cycles_1_n19)
         );
  NOR2_X4 aes_ctrl_lsfr_23_cycles_1_U29 ( .A1(aes_ctrl_lsfr_23_cycles_1_n23), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n17), .ZN(n453) );
  OAI22_X1 aes_ctrl_lsfr_23_cycles_1_U28 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n23), .B1(aes_ctrl_lsfr_23_cycles_1_n3), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n24), .ZN(aes_ctrl_lsfr_23_cycles_1_n39)
         );
  AOI221_X1 aes_ctrl_lsfr_23_cycles_1_U27 ( .B1(StartxSI), .B2(
        aes_ctrl_lsfr_23_cycles_1_n22), .C1(aes_ctrl_lsfr_23_cycles_1_n21), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n22), .A(aes_ctrl_lsfr_23_cycles_1_n8), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n3) );
  XNOR2_X1 aes_ctrl_lsfr_23_cycles_1_U26 ( .A(aes_ctrl_lsfr_23_cycles_1_n1), 
        .B(aes_ctrl_lsfr_23_cycles_1_n5), .ZN(aes_ctrl_lsfr_23_cycles_1_n36)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U25 ( .A1(aes_ctrl_lsfr_23_cycles_1_n22), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n19), .ZN(aes_ctrl_lsfr_23_cycles_1_n1)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U24 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_N16)
         );
  AOI211_X1 aes_ctrl_lsfr_23_cycles_1_U23 ( .C1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n11), .A(aes_ctrl_lsfr_23_cycles_1_n13), 
        .B(aes_ctrl_lsfr_23_cycles_1_n7), .ZN(aes_ctrl_lsfr_23_cycles_1_N66)
         );
  OAI22_X1 aes_ctrl_lsfr_23_cycles_1_U22 ( .A1(aes_ctrl_lsfr_23_cycles_1_n7), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n15), .B1(aes_ctrl_lsfr_23_cycles_1_n17), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_N83)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U21 ( .A1(aes_ctrl_lsfr_23_cycles_1_n6), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n17), .ZN(disableKeyRegsxS) );
  AOI22_X1 aes_ctrl_lsfr_23_cycles_1_U20 ( .A1(aes_ctrl_lsfr_23_cycles_1_n20), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .B1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n23), .ZN(aes_ctrl_lsfr_23_cycles_1_n37)
         );
  OAI221_X1 aes_ctrl_lsfr_23_cycles_1_U19 ( .B1(aes_ctrl_lsfr_23_cycles_1_n20), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n4), .C1(aes_ctrl_lsfr_23_cycles_1_n23), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n18), .A(aes_ctrl_lsfr_23_cycles_1_n22), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n35) );
  XNOR2_X1 aes_ctrl_lsfr_23_cycles_1_U18 ( .A(aes_ctrl_lsfr_23_cycles_1_n24), 
        .B(aes_ctrl_lsfr_23_cycles_1_n9), .ZN(aes_ctrl_lsfr_23_cycles_1_n38)
         );
  NOR4_X2 aes_ctrl_lsfr_23_cycles_1_U17 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(LastRoundxS), .A3(aes_ctrl_lsfr_23_cycles_1_n7), .A4(
        aes_ctrl_lsfr_23_cycles_1_n10), .ZN(doMixColumnsxS) );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U16 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .ZN(aes_ctrl_lsfr_23_cycles_1_n18)
         );
  NAND3_X1 aes_ctrl_lsfr_23_cycles_1_U15 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n9), .A3(aes_ctrl_lsfr_23_cycles_1_n6), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n14) );
  OAI21_X1 aes_ctrl_lsfr_23_cycles_1_U14 ( .B1(aes_ctrl_lsfr_23_cycles_1_n10), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n8), .A(aes_ctrl_lsfr_23_cycles_1_n5), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n11) );
  NOR2_X2 aes_ctrl_lsfr_23_cycles_1_U13 ( .A1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n11), .ZN(aes_ctrl_lsfr_23_cycles_1_n13)
         );
  INV_X1 aes_ctrl_lsfr_23_cycles_1_U12 ( .A(aes_ctrl_lsfr_23_cycles_1_n13), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n15) );
  AND2_X1 aes_ctrl_lsfr_23_cycles_1_U11 ( .A1(aes_ctrl_lsfr_23_cycles_1_n8), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n22), .ZN(aes_ctrl_lsfr_23_cycles_1_n24)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U10 ( .A1(aes_ctrl_lsfr_23_cycles_1_n19), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n5), .ZN(aes_ctrl_lsfr_23_cycles_1_n23)
         );
  OR2_X1 aes_ctrl_lsfr_23_cycles_1_U9 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .ZN(aes_ctrl_lsfr_23_cycles_1_n22)
         );
  OR3_X1 aes_ctrl_lsfr_23_cycles_1_U8 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n10), .A3(aes_ctrl_lsfr_23_cycles_1_n5), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n21) );
  INV_X1 aes_ctrl_lsfr_23_cycles_1_U7 ( .A(aes_ctrl_lsfr_23_cycles_1_n23), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n20) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U6 ( .A1(aes_ctrl_lsfr_23_cycles_1_n17), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n16), .ZN(StateKEYSCHEDULExS) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U5 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n21), .ZN(showRCONxS) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U4 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n16), .ZN(StateKEYADDITION1o3xS) );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U3 ( .A1(aes_ctrl_lsfr_23_cycles_1_n11), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_n16)
         );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_2_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n36), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n5), .QN(aes_ctrl_lsfr_23_cycles_1_n6) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_1_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n38), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n10), .QN(aes_ctrl_lsfr_23_cycles_1_n9) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_3_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n35), .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(
        aes_ctrl_lsfr_23_cycles_1_n4) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_4_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n37), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n7), .QN(aes_ctrl_lsfr_23_cycles_1_n2) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_0_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n39), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n8), .QN(aes_ctrl_lsfr_23_cycles_1_n12) );
  OAI22_X1 rcon_1_U34 ( .A1(rcon_1_n26), .A2(n453), .B1(rcon_1_n28), .B2(
        rcon_1_n39), .ZN(rcon_1_n19) );
  MUX2_X1 rcon_1_U33 ( .A(rcon_1_n35), .B(rcon_1_n36), .S(n453), .Z(rcon_1_n18) );
  INV_X2 rcon_1_U32 ( .A(rcon_1_n43), .ZN(n454) );
  AOI211_X1 rcon_1_U31 ( .C1(rcon_1_n37), .C2(rcon_1_n29), .A(rcon_1_n41), .B(
        rcon_1_n16), .ZN(rcon_1_n24) );
  AOI22_X1 rcon_1_U30 ( .A1(rcon_1_n34), .A2(rcon_1_n42), .B1(rcon_1_n40), 
        .B2(rcon_1_n17), .ZN(rcon_1_n16) );
  NOR2_X1 rcon_1_U29 ( .A1(rcon_1_n26), .A2(rcon_1_n38), .ZN(RCONxD[6]) );
  AOI211_X1 rcon_1_U28 ( .C1(rcon_1_n9), .C2(rcon_1_n14), .A(rcon_1_n41), .B(
        rcon_1_n15), .ZN(rcon_1_n22) );
  OAI22_X1 rcon_1_U27 ( .A1(n453), .A2(rcon_1_n4), .B1(rcon_1_n9), .B2(
        rcon_1_n40), .ZN(rcon_1_n15) );
  INV_X1 rcon_1_U26 ( .A(rcon_1_n42), .ZN(rcon_1_n14) );
  NOR2_X1 rcon_1_U25 ( .A1(rcon_1_n28), .A2(rcon_1_n38), .ZN(RCONxD[5]) );
  OAI211_X1 rcon_1_U24 ( .C1(n453), .C2(rcon_1_n17), .A(rcon_1_n42), .B(
        rcon_1_n13), .ZN(rcon_1_n25) );
  INV_X1 rcon_1_U23 ( .A(rcon_1_n41), .ZN(rcon_1_n13) );
  NOR2_X1 rcon_1_U22 ( .A1(rcon_1_n38), .A2(rcon_1_n32), .ZN(RCONxD[4]) );
  OAI21_X1 rcon_1_U21 ( .B1(n453), .B2(rcon_1_n32), .A(rcon_1_n12), .ZN(
        rcon_1_n21) );
  OAI211_X1 rcon_1_U20 ( .C1(rcon_1_n35), .C2(rcon_1_n4), .A(n453), .B(
        rcon_1_n11), .ZN(rcon_1_n12) );
  OAI21_X1 rcon_1_U19 ( .B1(rcon_1_n35), .B2(rcon_1_n33), .A(rcon_1_n4), .ZN(
        rcon_1_n11) );
  NOR2_X1 rcon_1_U18 ( .A1(rcon_1_n31), .A2(rcon_1_n38), .ZN(RCONxD[2]) );
  NOR2_X1 rcon_1_U17 ( .A1(rcon_1_n38), .A2(rcon_1_n30), .ZN(RCONxD[7]) );
  AND2_X1 rcon_1_U16 ( .A1(rcon_1_n4), .A2(showRCONxS), .ZN(RCONxD[3]) );
  NOR2_X1 rcon_1_U15 ( .A1(rcon_1_n38), .A2(rcon_1_n29), .ZN(RCONxD[1]) );
  NOR2_X1 rcon_1_U14 ( .A1(rcon_1_n17), .A2(rcon_1_n38), .ZN(RCONxD[0]) );
  OAI22_X1 rcon_1_U13 ( .A1(n453), .A2(rcon_1_n28), .B1(rcon_1_n32), .B2(
        rcon_1_n39), .ZN(rcon_1_n20) );
  OAI22_X1 rcon_1_U12 ( .A1(n453), .A2(rcon_1_n31), .B1(rcon_1_n29), .B2(
        rcon_1_n39), .ZN(rcon_1_n23) );
  NOR2_X1 rcon_1_U11 ( .A1(rcon_1_n26), .A2(rcon_1_n4), .ZN(rcon_1_n36) );
  NAND2_X1 rcon_1_U10 ( .A1(n453), .A2(rcon_1_n43), .ZN(rcon_1_n39) );
  NOR2_X1 rcon_1_U9 ( .A1(rcon_1_n43), .A2(rcon_1_n37), .ZN(rcon_1_n41) );
  NAND2_X1 rcon_1_U8 ( .A1(n453), .A2(rcon_1_n30), .ZN(rcon_1_n40) );
  NAND2_X1 rcon_1_U7 ( .A1(n453), .A2(rcon_1_n35), .ZN(rcon_1_n42) );
  INV_X1 rcon_1_U6 ( .A(n453), .ZN(rcon_1_n37) );
  INV_X1 rcon_1_U5 ( .A(showRCONxS), .ZN(rcon_1_n38) );
  NOR2_X1 rcon_1_U4 ( .A1(rcon_1_n28), .A2(rcon_1_n31), .ZN(LastRoundxS) );
  NAND2_X1 rcon_1_U3 ( .A1(rcon_1_n33), .A2(rcon_1_n4), .ZN(rcon_1_n43) );
  DFFR_X1 rcon_1_RCONxDP_reg_4_ ( .D(rcon_1_n21), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(rcon_1_n32) );
  DFFR_X1 rcon_1_RCONxDP_reg_1_ ( .D(rcon_1_n24), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(rcon_1_n29) );
  DFFR_X1 rcon_1_RCONxDP_reg_0_ ( .D(rcon_1_n25), .CK(ClkxCI), .RN(RstxBI), 
        .Q(rcon_1_n34), .QN(rcon_1_n17) );
  DFFR_X1 rcon_1_RCONxDP_reg_7_ ( .D(rcon_1_n18), .CK(ClkxCI), .RN(RstxBI), 
        .Q(rcon_1_n35), .QN(rcon_1_n30) );
  DFFS_X1 rcon_1_RCONxDP_reg_3_ ( .D(rcon_1_n22), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n4), .QN() );
  DFFS_X1 rcon_1_RCONxDP_reg_2_ ( .D(rcon_1_n23), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n9), .QN(rcon_1_n31) );
  DFFS_X1 rcon_1_RCONxDP_reg_5_ ( .D(rcon_1_n20), .CK(ClkxCI), .SN(RstxBI), 
        .Q(), .QN(rcon_1_n28) );
  DFFS_X1 rcon_1_RCONxDP_reg_6_ ( .D(rcon_1_n19), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n33), .QN(rcon_1_n26) );
  XOR2_X1 SBOX_Inst_f1_U12 ( .A(SBOX_Zh_f1[9]), .B(SBOX_Zl_f1_9_), .Z(
        SBOX_Inst_f1_sZ[9]) );
  XOR2_X1 SBOX_Inst_f1_U11 ( .A(SBOX_Zh_f1[8]), .B(SBOX_Zl_f1_8_), .Z(
        SBOX_ab2[8]) );
  XOR2_X1 SBOX_Inst_f1_U10 ( .A(SBOX_Zh_f1[5]), .B(SBOX_Zl_f1_5_), .Z(
        SBOX_Inst_f1_sZ[5]) );
  XOR2_X1 SBOX_Inst_f1_U9 ( .A(SBOX_Zh_f1[4]), .B(SBOX_Zl_f1_4_), .Z(
        SBOX_ab2[4]) );
  XOR2_X1 SBOX_Inst_f1_U8 ( .A(SBOX_Zh_f1[1]), .B(SBOX_Zl_f1_1_), .Z(
        SBOX_Inst_f1_sZ[1]) );
  XOR2_X1 SBOX_Inst_f1_U7 ( .A(SBOX_Zh_f1[0]), .B(SBOX_Zl_f1_0_), .Z(
        SBOX_ab2[0]) );
  XOR2_X1 SBOX_Inst_f1_U6 ( .A(SBOX_Zh_f1[2]), .B(CxDO[0]), .Z(
        SBOX_Inst_f1_sZ[2]) );
  XOR2_X1 SBOX_Inst_f1_U5 ( .A(SBOX_Zh_f1[10]), .B(CxDO[16]), .Z(
        SBOX_Inst_f1_sZ[10]) );
  XOR2_X1 SBOX_Inst_f1_U4 ( .A(SBOX_Zh_f1[3]), .B(SBOX_Zl_f1_3_), .Z(
        SBOX_Inst_f1_sZ[3]) );
  XOR2_X1 SBOX_Inst_f1_U3 ( .A(SBOX_Zh_f1[6]), .B(CxDO[8]), .Z(
        SBOX_Inst_f1_sZ[6]) );
  XOR2_X1 SBOX_Inst_f1_U2 ( .A(SBOX_Zh_f1[11]), .B(SBOX_Zl_f1_11_), .Z(
        SBOX_Inst_f1_sZ[11]) );
  XOR2_X1 SBOX_Inst_f1_U1 ( .A(SBOX_Zh_f1[7]), .B(SBOX_Zl_f1_7_), .Z(
        SBOX_Inst_f1_sZ[7]) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U42 ( .A(SBOX_Inst_f1_linearMapping_n25), 
        .B(SBOX_Inst_f1_linearMapping_n24), .ZN(SBOX_Inst_f1_linearMapping_n26) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U41 ( .A(SBOX_Inst_f1_linearMapping_n22), 
        .B(SBOX_Inst_f1_linearMapping_n21), .ZN(SBOX_Inst_f1_linearMapping_n23) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U40 ( .A(SBOX_Inst_f1_linearMapping_n19), 
        .B(SBOX_Inst_f1_linearMapping_n18), .ZN(SBOX_Inst_f1_linearMapping_n20) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U39 ( .A(CxDO[5]), .B(
        SBOX_Inst_f1_linearMapping_n14), .ZN(SBOX_Zl_f1_1_) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U38 ( .A(CxDO[1]), .B(SBOX_Zl_f1_1_), .Z(
        SBOX_Zh_f1[1]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U37 ( .A(CxDO[21]), .B(
        SBOX_Inst_f1_linearMapping_n15), .ZN(SBOX_Zl_f1_9_) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U36 ( .A(CxDO[17]), .B(SBOX_Zl_f1_9_), 
        .Z(SBOX_Zh_f1[9]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U35 ( .A(SBOX_Inst_f1_linearMapping_n30), 
        .B(SBOX_Inst_f1_linearMapping_n16), .ZN(SBOX_Zh_f1[4]) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U34 ( .A(CxDO[20]), .B(SBOX_Zl_f1_9_), 
        .Z(SBOX_Zh_f1[10]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U33 ( .A(SBOX_Inst_f1_linearMapping_n28), 
        .B(SBOX_Inst_f1_linearMapping_n27), .ZN(SBOX_Zh_f1[3]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U32 ( .A(SBOX_Inst_f1_linearMapping_n32), 
        .B(SBOX_Inst_f1_linearMapping_n15), .ZN(SBOX_Zh_f1[8]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U31 ( .A(CxDO[3]), .B(
        SBOX_Inst_f1_linearMapping_n27), .ZN(SBOX_Zl_f1_0_) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U30 ( .A(CxDO[13]), .B(
        SBOX_Inst_f1_linearMapping_n16), .ZN(SBOX_Zl_f1_5_) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U29 ( .A(CxDO[9]), .B(SBOX_Zl_f1_5_), .Z(
        SBOX_Zh_f1[5]) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U28 ( .A(CxDO[9]), .B(
        SBOX_Inst_f1_linearMapping_n20), .Z(SBOX_Zl_f1_7_) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U27 ( .A(CxDO[17]), .B(
        SBOX_Inst_f1_linearMapping_n23), .Z(SBOX_Zl_f1_11_) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U26 ( .A(CxDO[11]), .B(
        SBOX_Inst_f1_linearMapping_n29), .ZN(SBOX_Zl_f1_4_) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U25 ( .A(CxDO[4]), .B(SBOX_Zl_f1_1_), .Z(
        SBOX_Zh_f1[2]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U24 ( .A(CxDO[19]), .B(
        SBOX_Inst_f1_linearMapping_n31), .ZN(SBOX_Zl_f1_8_) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U23 ( .A(SBOX_Inst_f1_linearMapping_n28), 
        .B(SBOX_Inst_f1_linearMapping_n14), .ZN(SBOX_Zh_f1[0]) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U22 ( .A(CxDO[1]), .B(
        SBOX_Inst_f1_linearMapping_n26), .Z(SBOX_Zl_f1_3_) );
  XOR2_X2 SBOX_Inst_f1_linearMapping_U21 ( .A(CxDO[12]), .B(SBOX_Zl_f1_5_), 
        .Z(SBOX_Zh_f1[6]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U20 ( .A(SBOX_Inst_f1_linearMapping_n32), 
        .B(SBOX_Inst_f1_linearMapping_n31), .ZN(SBOX_Zh_f1[11]) );
  XNOR2_X2 SBOX_Inst_f1_linearMapping_U19 ( .A(SBOX_Inst_f1_linearMapping_n30), 
        .B(SBOX_Inst_f1_linearMapping_n29), .ZN(SBOX_Zh_f1[7]) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U18 ( .A(SBOX_Inst_f1_linearMapping_n13), 
        .B(SBOX_Inst_f1_linearMapping_n15), .ZN(SBOX_Inst_f1_linearMapping_n31) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U17 ( .A(CxDO[18]), .B(CxDO[17]), .ZN(
        SBOX_Inst_f1_linearMapping_n13) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U16 ( .A(SBOX_Inst_f1_linearMapping_n12), 
        .B(SBOX_Inst_f1_linearMapping_n14), .ZN(SBOX_Inst_f1_linearMapping_n27) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U15 ( .A(CxDO[2]), .B(CxDO[1]), .ZN(
        SBOX_Inst_f1_linearMapping_n12) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U14 ( .A(CxDO[16]), .B(CxDO[19]), .ZN(
        SBOX_Inst_f1_linearMapping_n21) );
  XOR2_X1 SBOX_Inst_f1_linearMapping_U13 ( .A(CxDO[23]), .B(CxDO[20]), .Z(
        SBOX_Inst_f1_linearMapping_n22) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U12 ( .A(CxDO[8]), .B(CxDO[11]), .ZN(
        SBOX_Inst_f1_linearMapping_n18) );
  XOR2_X1 SBOX_Inst_f1_linearMapping_U11 ( .A(CxDO[15]), .B(CxDO[12]), .Z(
        SBOX_Inst_f1_linearMapping_n19) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U10 ( .A(CxDO[0]), .B(CxDO[3]), .ZN(
        SBOX_Inst_f1_linearMapping_n24) );
  XOR2_X1 SBOX_Inst_f1_linearMapping_U9 ( .A(CxDO[7]), .B(CxDO[4]), .Z(
        SBOX_Inst_f1_linearMapping_n25) );
  XOR2_X1 SBOX_Inst_f1_linearMapping_U8 ( .A(CxDO[23]), .B(CxDO[21]), .Z(
        SBOX_Inst_f1_linearMapping_n32) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U7 ( .A(CxDO[16]), .B(CxDO[22]), .ZN(
        SBOX_Inst_f1_linearMapping_n15) );
  XOR2_X1 SBOX_Inst_f1_linearMapping_U6 ( .A(CxDO[15]), .B(CxDO[13]), .Z(
        SBOX_Inst_f1_linearMapping_n30) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U5 ( .A(CxDO[10]), .B(CxDO[9]), .ZN(
        SBOX_Inst_f1_linearMapping_n17) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U4 ( .A(SBOX_Inst_f1_linearMapping_n17), 
        .B(SBOX_Inst_f1_linearMapping_n16), .ZN(SBOX_Inst_f1_linearMapping_n29) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U3 ( .A(CxDO[14]), .B(CxDO[8]), .ZN(
        SBOX_Inst_f1_linearMapping_n16) );
  XOR2_X1 SBOX_Inst_f1_linearMapping_U2 ( .A(CxDO[7]), .B(CxDO[5]), .Z(
        SBOX_Inst_f1_linearMapping_n28) );
  XNOR2_X1 SBOX_Inst_f1_linearMapping_U1 ( .A(CxDO[0]), .B(CxDO[6]), .ZN(
        SBOX_Inst_f1_linearMapping_n14) );
  XOR2_X1 SBOX_Inst_f1_abSQ_U6 ( .A(SBOX_ab2[0]), .B(SBOX_Inst_f1_sZ[2]), .Z(
        SBOX_ab2[3]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_U5 ( .A(SBOX_Inst_f1_sZ[10]), .B(SBOX_ab2[8]), .Z(
        SBOX_ab2[11]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_U4 ( .A(SBOX_Inst_f1_sZ[1]), .B(SBOX_Inst_f1_sZ[3]), .Z(SBOX_ab2[2]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_U3 ( .A(SBOX_ab2[4]), .B(SBOX_Inst_f1_sZ[6]), .Z(
        SBOX_ab2[7]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_U2 ( .A(SBOX_Inst_f1_sZ[11]), .B(
        SBOX_Inst_f1_sZ[9]), .Z(SBOX_ab2[10]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_U1 ( .A(SBOX_Inst_f1_sZ[5]), .B(SBOX_Inst_f1_sZ[7]), .Z(SBOX_ab2[6]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_NxGamma_U3 ( .A(SBOX_ab2[0]), .B(
        SBOX_Inst_f1_sZ[1]), .Z(SBOX_ab2[1]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_NxGamma_U2 ( .A(SBOX_ab2[8]), .B(
        SBOX_Inst_f1_sZ[9]), .Z(SBOX_ab2[9]) );
  XOR2_X1 SBOX_Inst_f1_abSQ_NxGamma_U1 ( .A(SBOX_ab2[4]), .B(
        SBOX_Inst_f1_sZ[5]), .Z(SBOX_ab2[5]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U12 ( .A(SBOX_Zl_f1_11_), .B(SBOX_Zl_f1_9_), 
        .Z(SBOX_Inst_f1_phpplmul_sB[5]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U11 ( .A(SBOX_Zl_f1_5_), .B(SBOX_Zl_f1_7_), 
        .Z(SBOX_Inst_f1_phpplmul_sB[3]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U10 ( .A(SBOX_Zl_f1_1_), .B(SBOX_Zl_f1_3_), 
        .Z(SBOX_Inst_f1_phpplmul_sB[1]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U9 ( .A(SBOX_Zl_f1_0_), .B(CxDO[0]), .Z(
        SBOX_Inst_f1_phpplmul_sB[0]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U8 ( .A(SBOX_Zh_f1[10]), .B(SBOX_Zh_f1[8]), 
        .Z(SBOX_Inst_f1_phpplmul_sA[4]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U7 ( .A(SBOX_Zh_f1[4]), .B(SBOX_Zh_f1[6]), .Z(
        SBOX_Inst_f1_phpplmul_sA[2]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U6 ( .A(SBOX_Zh_f1[1]), .B(SBOX_Zh_f1[3]), .Z(
        SBOX_Inst_f1_phpplmul_sA[1]) );
  XOR2_X2 SBOX_Inst_f1_phpplmul_U5 ( .A(SBOX_Zh_f1[11]), .B(SBOX_Zh_f1[9]), 
        .Z(SBOX_Inst_f1_phpplmul_sA[5]) );
  XOR2_X2 SBOX_Inst_f1_phpplmul_U4 ( .A(CxDO[16]), .B(SBOX_Zl_f1_8_), .Z(
        SBOX_Inst_f1_phpplmul_sB[4]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U3 ( .A(SBOX_Zh_f1[0]), .B(SBOX_Zh_f1[2]), .Z(
        SBOX_Inst_f1_phpplmul_sA[0]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U2 ( .A(SBOX_Zh_f1[5]), .B(SBOX_Zh_f1[7]), .Z(
        SBOX_Inst_f1_phpplmul_sA[3]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_U1 ( .A(SBOX_Zl_f1_4_), .B(CxDO[8]), .Z(
        SBOX_Inst_f1_phpplmul_sB[2]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U103 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n160), .B(SBOX_Inst_f1_phpplmul_himul_n159), .ZN(SBOX_Inst_f1_phpplmul_himul_n165) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_himul_U102 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n158), .B(SBOX_Inst_f1_phpplmul_himul_n157), .Z(SBOX_Inst_f1_phpplmul_himul_n159) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U101 ( .A1(SBOX_Zh_f1[6]), .A2(
        SBOX_Zh_f1[2]), .B1(SBOX_Inst_f1_phpplmul_himul_n171), .B2(
        SBOX_Inst_f1_phpplmul_himul_n172), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n169) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_himul_U100 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n150), .B(SBOX_Inst_f1_phpplmul_himul_n149), .Z(SBOX_Inst_f1_phpplmul_himul_n153) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U99 ( .A1(SBOX_Zh_f1[10]), .A2(
        SBOX_Zh_f1[11]), .B1(SBOX_Inst_f1_phpplmul_himul_n154), .B2(
        SBOX_Inst_f1_phpplmul_himul_n148), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n155) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_himul_U98 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n146), .B(SBOX_Inst_f1_phpplmul_himul_n147), .Z(SBOX_Inst_f1_phpplmul_himul_n161) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U97 ( .A1(SBOX_Zl_f1_3_), .A2(
        SBOX_Zh_f1[2]), .ZN(SBOX_Inst_f1_phpplmul_himul_n147) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U96 ( .A1(SBOX_Zh_f1[3]), .A2(CxDO[0]), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n146) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U95 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n145), .B(SBOX_Inst_f1_phpplmul_himul_n144), .ZN(SBOX_Inst_f1_phpplmul_Orig_ph[4]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U94 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n161), .B(SBOX_Inst_f1_phpplmul_himul_n141), .ZN(SBOX_Inst_f1_phpplmul_himul_n145) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U93 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n142), .B(SBOX_Inst_f1_phpplmul_himul_n143), .ZN(SBOX_Inst_f1_phpplmul_himul_n144) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U92 ( .A1(SBOX_Zl_f1_7_), .A2(
        SBOX_Inst_f1_phpplmul_himul_n166), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n143) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U91 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n172), .A2(
        SBOX_Inst_f1_phpplmul_himul_n162), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n142) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U90 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n165), .B(SBOX_Inst_f1_phpplmul_himul_n140), .ZN(SBOX_Inst_f1_phpplmul_himul_n141) );
  MUX2_X1 SBOX_Inst_f1_phpplmul_himul_U89 ( .A(CxDO[0]), .B(SBOX_Zl_f1_3_), 
        .S(SBOX_Inst_f1_phpplmul_himul_n139), .Z(
        SBOX_Inst_f1_phpplmul_himul_n140) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U88 ( .A1(SBOX_Zh_f1[7]), .A2(
        SBOX_Zh_f1[3]), .B1(SBOX_Inst_f1_phpplmul_himul_n166), .B2(
        SBOX_Inst_f1_phpplmul_himul_n163), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n139) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U87 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n137), .B(SBOX_Inst_f1_phpplmul_himul_n138), .ZN(SBOX_Inst_f1_phpplmul_Orig_ph[5]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_himul_U86 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n133), .B(SBOX_Inst_f1_phpplmul_himul_n135), .Z(SBOX_Inst_f1_phpplmul_himul_n138) );
  AOI211_X1 SBOX_Inst_f1_phpplmul_himul_U85 ( .C1(CxDO[0]), .C2(SBOX_Zl_f1_7_), 
        .A(SBOX_Inst_f1_phpplmul_himul_n136), .B(
        SBOX_Inst_f1_phpplmul_himul_n163), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n137) );
  AND2_X1 SBOX_Inst_f1_phpplmul_himul_U84 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n168), .A2(
        SBOX_Inst_f1_phpplmul_himul_n164), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n136) );
  AOI211_X1 SBOX_Inst_f1_phpplmul_himul_U83 ( .C1(SBOX_Zh_f1[2]), .C2(
        SBOX_Zh_f1[6]), .A(SBOX_Inst_f1_phpplmul_himul_n170), .B(
        SBOX_Inst_f1_phpplmul_himul_n134), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n135) );
  AND2_X1 SBOX_Inst_f1_phpplmul_himul_U82 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n171), .A2(
        SBOX_Inst_f1_phpplmul_himul_n172), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n134) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U81 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n131), .B(SBOX_Inst_f1_phpplmul_himul_n132), .ZN(SBOX_Inst_f1_phpplmul_himul_n133) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U80 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n167), .A2(
        SBOX_Inst_f1_phpplmul_himul_n166), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n132) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U79 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n165), .B(SBOX_Inst_f1_phpplmul_himul_n130), .ZN(SBOX_Inst_f1_phpplmul_himul_n131) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U78 ( .A1(SBOX_Zh_f1[3]), .A2(
        SBOX_Inst_f1_phpplmul_himul_n168), .B1(CxDO[0]), .B2(
        SBOX_Inst_f1_phpplmul_himul_n169), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n130) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U77 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n129), .B(SBOX_Inst_f1_phpplmul_himul_n128), .ZN(SBOX_Inst_f1_phpplmul_Orig_ph[3]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U76 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n124), .B(SBOX_Inst_f1_phpplmul_himul_n126), .ZN(SBOX_Inst_f1_phpplmul_himul_n129) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_himul_U75 ( .B1(
        SBOX_Inst_f1_phpplmul_himul_n118), .B2(SBOX_Zh_f1[3]), .C1(
        SBOX_Inst_f1_phpplmul_himul_n127), .C2(
        SBOX_Inst_f1_phpplmul_himul_n166), .A(CxDO[16]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n128) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U74 ( .A(SBOX_Inst_f1_phpplmul_himul_n118), .ZN(SBOX_Inst_f1_phpplmul_himul_n127) );
  OAI21_X1 SBOX_Inst_f1_phpplmul_himul_U73 ( .B1(
        SBOX_Inst_f1_phpplmul_himul_n156), .B2(
        SBOX_Inst_f1_phpplmul_himul_n155), .A(SBOX_Inst_f1_phpplmul_himul_n125), .ZN(SBOX_Inst_f1_phpplmul_himul_n126) );
  NAND3_X1 SBOX_Inst_f1_phpplmul_himul_U72 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n156), .A2(SBOX_Zh_f1[10]), .A3(
        SBOX_Inst_f1_phpplmul_himul_n154), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n125) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U71 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n122), .B(SBOX_Inst_f1_phpplmul_himul_n123), .ZN(SBOX_Inst_f1_phpplmul_himul_n124) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U70 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n118), .A2(SBOX_Zl_f1_11_), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n123) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_himul_U69 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n153), .B(SBOX_Inst_f1_phpplmul_himul_n121), .Z(SBOX_Inst_f1_phpplmul_himul_n122) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_himul_U68 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n119), .B(SBOX_Inst_f1_phpplmul_himul_n120), .Z(SBOX_Inst_f1_phpplmul_himul_n121) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U67 ( .A1(CxDO[0]), .A2(SBOX_Zh_f1[10]), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n120) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U66 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n167), .A2(SBOX_Zh_f1[3]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n119) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U65 ( .A1(SBOX_Zh_f1[11]), .A2(
        SBOX_Zh_f1[2]), .B1(SBOX_Inst_f1_phpplmul_himul_n154), .B2(
        SBOX_Inst_f1_phpplmul_himul_n171), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n118) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U64 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n161), .B(SBOX_Inst_f1_phpplmul_himul_n117), .ZN(SBOX_Inst_f1_phpplmul_Orig_ph[2]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U63 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n115), .B(SBOX_Inst_f1_phpplmul_himul_n116), .ZN(SBOX_Inst_f1_phpplmul_himul_n117) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U62 ( .A1(SBOX_Zh_f1[2]), .A2(
        SBOX_Zl_f1_11_), .ZN(SBOX_Inst_f1_phpplmul_himul_n116) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_himul_U61 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n114), .B(SBOX_Inst_f1_phpplmul_himul_n153), .Z(SBOX_Inst_f1_phpplmul_himul_n115) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U60 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n112), .B(SBOX_Inst_f1_phpplmul_himul_n113), .ZN(SBOX_Inst_f1_phpplmul_himul_n114) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U59 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n109), .B(SBOX_Inst_f1_phpplmul_himul_n110), .ZN(SBOX_Inst_f1_phpplmul_himul_n113) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U58 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n106), .A2(
        SBOX_Inst_f1_phpplmul_himul_n111), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n112) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_himul_U57 ( .A1(CxDO[16]), .A2(SBOX_Zl_f1_11_), .B1(SBOX_Inst_f1_phpplmul_himul_n152), .B2(SBOX_Inst_f1_phpplmul_himul_n151), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n111) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U56 ( .A1(SBOX_Zh_f1[3]), .A2(CxDO[0]), 
        .B1(SBOX_Inst_f1_phpplmul_himul_n166), .B2(
        SBOX_Inst_f1_phpplmul_himul_n168), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n110) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U55 ( .A1(SBOX_Zh_f1[11]), .A2(
        SBOX_Inst_f1_phpplmul_himul_n107), .B1(CxDO[16]), .B2(
        SBOX_Inst_f1_phpplmul_himul_n108), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n109) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U54 ( .A(SBOX_Zh_f1[11]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n108) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U53 ( .A1(SBOX_Zl_f1_3_), .A2(
        SBOX_Zl_f1_11_), .B1(SBOX_Inst_f1_phpplmul_himul_n152), .B2(
        SBOX_Inst_f1_phpplmul_himul_n167), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n107) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U52 ( .A(SBOX_Zh_f1[3]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n106) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U51 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n103), .B(SBOX_Inst_f1_phpplmul_himul_n105), .ZN(SBOX_Inst_f1_phpplmul_Orig_ph[1]) );
  AOI211_X1 SBOX_Inst_f1_phpplmul_himul_U50 ( .C1(SBOX_Zh_f1[10]), .C2(
        SBOX_Zh_f1[6]), .A(SBOX_Inst_f1_phpplmul_himul_n162), .B(
        SBOX_Inst_f1_phpplmul_himul_n104), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n105) );
  AND2_X1 SBOX_Inst_f1_phpplmul_himul_U49 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n148), .A2(
        SBOX_Inst_f1_phpplmul_himul_n172), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n104) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U48 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n102), .B(SBOX_Inst_f1_phpplmul_himul_n99), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n103) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U47 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n101), .A2(
        SBOX_Inst_f1_phpplmul_himul_n100), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n102) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_himul_U46 ( .A1(SBOX_Zh_f1[7]), .A2(
        SBOX_Zh_f1[10]), .B1(SBOX_Inst_f1_phpplmul_himul_n148), .B2(
        SBOX_Inst_f1_phpplmul_himul_n163), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n101) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U45 ( .A(CxDO[16]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n100) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U44 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n97), .B(SBOX_Inst_f1_phpplmul_himul_n98), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n99) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U43 ( .A(SBOX_Zh_f1[10]), .B(
        SBOX_Inst_f1_phpplmul_himul_n95), .ZN(SBOX_Inst_f1_phpplmul_himul_n98)
         );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U42 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n90), .A2(SBOX_Inst_f1_phpplmul_himul_n96), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n97) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_himul_U41 ( .A1(CxDO[8]), .A2(SBOX_Zl_f1_7_), 
        .B1(SBOX_Inst_f1_phpplmul_himul_n170), .B2(
        SBOX_Inst_f1_phpplmul_himul_n164), .ZN(SBOX_Inst_f1_phpplmul_himul_n96) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U40 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n94), .B(SBOX_Inst_f1_phpplmul_himul_n93), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n95) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U39 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n91), .A2(SBOX_Inst_f1_phpplmul_himul_n154), .ZN(SBOX_Inst_f1_phpplmul_himul_n94) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_himul_U38 ( .B1(
        SBOX_Inst_f1_phpplmul_himul_n91), .B2(CxDO[16]), .C1(
        SBOX_Inst_f1_phpplmul_himul_n92), .C2(SBOX_Inst_f1_phpplmul_himul_n151), .A(SBOX_Zh_f1[6]), .ZN(SBOX_Inst_f1_phpplmul_himul_n93) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U37 ( .A(SBOX_Inst_f1_phpplmul_himul_n91), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n92) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U36 ( .A1(SBOX_Zl_f1_11_), .A2(CxDO[8]), 
        .B1(SBOX_Inst_f1_phpplmul_himul_n170), .B2(
        SBOX_Inst_f1_phpplmul_himul_n152), .ZN(SBOX_Inst_f1_phpplmul_himul_n91) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U35 ( .A(SBOX_Zh_f1[7]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n90) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U34 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n87), .B(SBOX_Inst_f1_phpplmul_himul_n89), 
        .ZN(SBOX_Inst_f1_phpplmul_Orig_ph[0]) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_himul_U33 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n152), .A2(SBOX_Inst_f1_phpplmul_himul_n88), .B1(SBOX_Inst_f1_phpplmul_himul_n156), .B2(CxDO[16]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n89) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U32 ( .A1(CxDO[16]), .A2(SBOX_Zh_f1[10]), .ZN(SBOX_Inst_f1_phpplmul_himul_n88) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U31 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n86), .B(SBOX_Inst_f1_phpplmul_himul_n85), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n87) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U30 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n155), .A2(SBOX_Zl_f1_7_), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n86) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U29 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n84), .B(SBOX_Inst_f1_phpplmul_himul_n78), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n85) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_himul_U28 ( .A(
        SBOX_Inst_f1_phpplmul_himul_n83), .B(SBOX_Inst_f1_phpplmul_himul_n80), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n84) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U27 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n82), .A2(SBOX_Inst_f1_phpplmul_himul_n81), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n83) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_himul_U26 ( .A1(SBOX_Zh_f1[11]), .A2(
        SBOX_Zh_f1[7]), .B1(SBOX_Inst_f1_phpplmul_himul_n154), .B2(
        SBOX_Inst_f1_phpplmul_himul_n163), .ZN(SBOX_Inst_f1_phpplmul_himul_n82) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U25 ( .A(CxDO[8]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n81) );
  OAI211_X1 SBOX_Inst_f1_phpplmul_himul_U24 ( .C1(CxDO[8]), .C2(SBOX_Zl_f1_11_), .A(SBOX_Zh_f1[6]), .B(SBOX_Inst_f1_phpplmul_himul_n79), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n80) );
  OR2_X1 SBOX_Inst_f1_phpplmul_himul_U23 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n152), .A2(
        SBOX_Inst_f1_phpplmul_himul_n170), .ZN(SBOX_Inst_f1_phpplmul_himul_n79) );
  OAI211_X1 SBOX_Inst_f1_phpplmul_himul_U22 ( .C1(
        SBOX_Inst_f1_phpplmul_himul_n76), .C2(CxDO[16]), .A(SBOX_Zh_f1[7]), 
        .B(SBOX_Inst_f1_phpplmul_himul_n77), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n78) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U21 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n76), .A2(CxDO[16]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n77) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U20 ( .A1(SBOX_Zl_f1_7_), .A2(
        SBOX_Zl_f1_11_), .B1(SBOX_Inst_f1_phpplmul_himul_n152), .B2(
        SBOX_Inst_f1_phpplmul_himul_n164), .ZN(SBOX_Inst_f1_phpplmul_himul_n76) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U19 ( .A(SBOX_Zh_f1[3]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n166) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U18 ( .A(SBOX_Zh_f1[6]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n172) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U17 ( .A1(SBOX_Zh_f1[2]), .A2(
        SBOX_Zl_f1_7_), .ZN(SBOX_Inst_f1_phpplmul_himul_n157) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U16 ( .A1(SBOX_Zh_f1[3]), .A2(CxDO[8]), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n158) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U15 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n169), .A2(SBOX_Zl_f1_3_), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n160) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U14 ( .A(SBOX_Zh_f1[7]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n163) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U13 ( .A(CxDO[0]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n168) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U12 ( .A(SBOX_Zl_f1_7_), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n164) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U11 ( .A(CxDO[8]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n170) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U10 ( .A(SBOX_Zh_f1[2]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n171) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U9 ( .A(SBOX_Zl_f1_3_), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n167) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_himul_U8 ( .A1(SBOX_Zl_f1_7_), .A2(
        SBOX_Inst_f1_phpplmul_himul_n170), .B1(CxDO[8]), .B2(
        SBOX_Inst_f1_phpplmul_himul_n164), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n162) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_himul_U7 ( .A1(
        SBOX_Inst_f1_phpplmul_himul_n148), .A2(
        SBOX_Inst_f1_phpplmul_himul_n152), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n156) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U6 ( .A1(SBOX_Zl_f1_3_), .A2(
        SBOX_Zh_f1[10]), .ZN(SBOX_Inst_f1_phpplmul_himul_n149) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_himul_U5 ( .A1(CxDO[0]), .A2(SBOX_Zh_f1[11]), 
        .ZN(SBOX_Inst_f1_phpplmul_himul_n150) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U4 ( .A(SBOX_Zh_f1[11]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n154) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U3 ( .A(SBOX_Zl_f1_11_), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n152) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U2 ( .A(CxDO[16]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n151) );
  INV_X1 SBOX_Inst_f1_phpplmul_himul_U1 ( .A(SBOX_Zh_f1[10]), .ZN(
        SBOX_Inst_f1_phpplmul_himul_n148) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U8 ( .A(
        SBOX_Inst_f1_phpplmul_AddNewMaskph_n6), .B(PRNGQ[2]), .ZN(SBOX_ph[4])
         );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U7 ( .A(PRNGQ[0]), .B(
        SBOX_Inst_f1_phpplmul_Orig_ph[4]), .ZN(
        SBOX_Inst_f1_phpplmul_AddNewMaskph_n6) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U6 ( .A(
        SBOX_Inst_f1_phpplmul_AddNewMaskph_n5), .B(PRNGQ[3]), .ZN(SBOX_ph[5])
         );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U5 ( .A(PRNGQ[1]), .B(
        SBOX_Inst_f1_phpplmul_Orig_ph[5]), .ZN(
        SBOX_Inst_f1_phpplmul_AddNewMaskph_n5) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U4 ( .A(PRNGQ[3]), .B(
        SBOX_Inst_f1_phpplmul_Orig_ph[3]), .Z(SBOX_ph[3]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U3 ( .A(PRNGQ[2]), .B(
        SBOX_Inst_f1_phpplmul_Orig_ph[2]), .Z(SBOX_ph[2]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U2 ( .A(PRNGQ[1]), .B(
        SBOX_Inst_f1_phpplmul_Orig_ph[1]), .Z(SBOX_ph[1]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskph_U1 ( .A(PRNGQ[0]), .B(
        SBOX_Inst_f1_phpplmul_Orig_ph[0]), .Z(SBOX_ph[0]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U92 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n288), .B(
        SBOX_Inst_f1_phpplmul_summul_n287), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n293) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_summul_U91 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n286), .B(
        SBOX_Inst_f1_phpplmul_summul_n285), .Z(
        SBOX_Inst_f1_phpplmul_summul_n287) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U90 ( .A1(SBOX_Inst_f1_phpplmul_sA[1]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[2]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n286) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U89 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n297), .A2(SBOX_Inst_f1_phpplmul_sB[1]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n288) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U88 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n284), .B(
        SBOX_Inst_f1_phpplmul_summul_n283), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_p[3]) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_summul_U87 ( .B1(SBOX_Inst_f1_phpplmul_sA[1]), .B2(SBOX_Inst_f1_phpplmul_summul_n282), .C1(
        SBOX_Inst_f1_phpplmul_summul_n294), .C2(
        SBOX_Inst_f1_phpplmul_summul_n281), .A(SBOX_Inst_f1_phpplmul_sB[4]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n283) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U86 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n280), .B(
        SBOX_Inst_f1_phpplmul_summul_n279), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n284) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U85 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n275), .B(
        SBOX_Inst_f1_phpplmul_summul_n274), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n280) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U84 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n282), .A2(SBOX_Inst_f1_phpplmul_sB[5]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n274) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_summul_U83 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n271), .B(
        SBOX_Inst_f1_phpplmul_summul_n270), .Z(
        SBOX_Inst_f1_phpplmul_summul_n272) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U82 ( .A1(SBOX_Inst_f1_phpplmul_sA[1]), 
        .A2(SBOX_Inst_f1_phpplmul_summul_n295), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n270) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U81 ( .A1(SBOX_Inst_f1_phpplmul_sB[0]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[4]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n271) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U80 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n269), .B(
        SBOX_Inst_f1_phpplmul_summul_n268), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_p[2]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U79 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n267), .B(
        SBOX_Inst_f1_phpplmul_summul_n266), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n268) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_summul_U78 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n265), .B(
        SBOX_Inst_f1_phpplmul_summul_n264), .Z(
        SBOX_Inst_f1_phpplmul_summul_n267) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U77 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n263), .B(
        SBOX_Inst_f1_phpplmul_summul_n262), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n264) );
  MUX2_X1 SBOX_Inst_f1_phpplmul_summul_U76 ( .A(SBOX_Inst_f1_phpplmul_sB[4]), 
        .B(SBOX_Inst_f1_phpplmul_summul_n261), .S(SBOX_Inst_f1_phpplmul_sA[5]), 
        .Z(SBOX_Inst_f1_phpplmul_summul_n262) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U75 ( .A1(SBOX_Inst_f1_phpplmul_sB[5]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[1]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n295), .B2(
        SBOX_Inst_f1_phpplmul_summul_n260), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n261) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_summul_U74 ( .B1(SBOX_Inst_f1_phpplmul_sB[5]), .B2(SBOX_Inst_f1_phpplmul_sB[4]), .C1(SBOX_Inst_f1_phpplmul_summul_n260), 
        .C2(SBOX_Inst_f1_phpplmul_summul_n259), .A(SBOX_Inst_f1_phpplmul_sA[1]), .ZN(SBOX_Inst_f1_phpplmul_summul_n263) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U73 ( .A1(SBOX_Inst_f1_phpplmul_sA[1]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[0]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n296), .B2(
        SBOX_Inst_f1_phpplmul_summul_n294), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n265) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U72 ( .A(SBOX_Inst_f1_phpplmul_sA[1]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n294) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_summul_U71 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n258), .B(
        SBOX_Inst_f1_phpplmul_summul_n257), .Z(
        SBOX_Inst_f1_phpplmul_summul_n273) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U70 ( .A1(SBOX_Inst_f1_phpplmul_sB[1]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[4]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n257) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U69 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n256), .B(
        SBOX_Inst_f1_phpplmul_summul_n255), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_p[1]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U68 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n254), .B(
        SBOX_Inst_f1_phpplmul_summul_n253), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n255) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_summul_U67 ( .B1(SBOX_Inst_f1_phpplmul_sA[4]), .B2(SBOX_Inst_f1_phpplmul_sA[3]), .C1(SBOX_Inst_f1_phpplmul_summul_n252), 
        .C2(SBOX_Inst_f1_phpplmul_summul_n291), .A(SBOX_Inst_f1_phpplmul_sB[4]), .ZN(SBOX_Inst_f1_phpplmul_summul_n253) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U66 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n251), .B(
        SBOX_Inst_f1_phpplmul_summul_n250), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n254) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_summul_U65 ( .B1(SBOX_Inst_f1_phpplmul_sB[3]), .B2(SBOX_Inst_f1_phpplmul_sB[2]), .C1(SBOX_Inst_f1_phpplmul_summul_n292), 
        .C2(SBOX_Inst_f1_phpplmul_summul_n298), .A(SBOX_Inst_f1_phpplmul_sA[3]), .ZN(SBOX_Inst_f1_phpplmul_summul_n250) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U64 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n249), .B(SBOX_Inst_f1_phpplmul_sA[4]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n251) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U63 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n248), .B(
        SBOX_Inst_f1_phpplmul_summul_n247), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n249) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_summul_U62 ( .B1(SBOX_Inst_f1_phpplmul_sB[4]), .B2(SBOX_Inst_f1_phpplmul_summul_n246), .C1(
        SBOX_Inst_f1_phpplmul_summul_n259), .C2(
        SBOX_Inst_f1_phpplmul_summul_n245), .A(SBOX_Inst_f1_phpplmul_sA[2]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n247) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U61 ( .A1(SBOX_Inst_f1_phpplmul_sB[5]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[2]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n298), .B2(
        SBOX_Inst_f1_phpplmul_summul_n260), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n246) );
  AOI221_X1 SBOX_Inst_f1_phpplmul_summul_U60 ( .B1(SBOX_Inst_f1_phpplmul_sA[4]), .B2(SBOX_Inst_f1_phpplmul_sA[2]), .C1(SBOX_Inst_f1_phpplmul_summul_n252), 
        .C2(SBOX_Inst_f1_phpplmul_summul_n300), .A(
        SBOX_Inst_f1_phpplmul_summul_n290), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n256) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U59 ( .A1(SBOX_Inst_f1_phpplmul_sB[3]), 
        .A2(SBOX_Inst_f1_phpplmul_summul_n298), .B1(
        SBOX_Inst_f1_phpplmul_sB[2]), .B2(SBOX_Inst_f1_phpplmul_summul_n292), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n290) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U58 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n244), .B(
        SBOX_Inst_f1_phpplmul_summul_n243), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_p[0]) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U57 ( .A1(SBOX_Inst_f1_phpplmul_sA[4]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[4]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n242) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U56 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n241), .B(
        SBOX_Inst_f1_phpplmul_summul_n240), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n244) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U55 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n277), .A2(SBOX_Inst_f1_phpplmul_sB[3]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n240) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U54 ( .A1(SBOX_Inst_f1_phpplmul_sA[4]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[5]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n276), .B2(
        SBOX_Inst_f1_phpplmul_summul_n252), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n277) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U53 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n239), .B(
        SBOX_Inst_f1_phpplmul_summul_n238), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n241) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U52 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n237), .B(
        SBOX_Inst_f1_phpplmul_summul_n236), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n238) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U51 ( .A1(SBOX_Inst_f1_phpplmul_sB[5]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[3]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n292), .B2(
        SBOX_Inst_f1_phpplmul_summul_n260), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n235) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_summul_U50 ( .B1(SBOX_Inst_f1_phpplmul_sB[5]), .B2(SBOX_Inst_f1_phpplmul_sB[2]), .C1(SBOX_Inst_f1_phpplmul_summul_n260), 
        .C2(SBOX_Inst_f1_phpplmul_summul_n298), .A(SBOX_Inst_f1_phpplmul_sA[2]), .ZN(SBOX_Inst_f1_phpplmul_summul_n237) );
  OAI21_X1 SBOX_Inst_f1_phpplmul_summul_U49 ( .B1(
        SBOX_Inst_f1_phpplmul_summul_n278), .B2(
        SBOX_Inst_f1_phpplmul_summul_n277), .A(
        SBOX_Inst_f1_phpplmul_summul_n233), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n279) );
  NAND3_X1 SBOX_Inst_f1_phpplmul_summul_U48 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n278), .A2(
        SBOX_Inst_f1_phpplmul_summul_n276), .A3(SBOX_Inst_f1_phpplmul_sA[4]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n233) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_summul_U47 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n231), .B(
        SBOX_Inst_f1_phpplmul_summul_n232), .Z(
        SBOX_Inst_f1_phpplmul_summul_n289) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U46 ( .A1(SBOX_Inst_f1_phpplmul_sB[1]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[0]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n232) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U45 ( .A1(SBOX_Inst_f1_phpplmul_sA[1]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[0]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n231) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U44 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n229), .B(
        SBOX_Inst_f1_phpplmul_summul_n230), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_p[5]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_summul_U43 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n225), .B(
        SBOX_Inst_f1_phpplmul_summul_n227), .Z(
        SBOX_Inst_f1_phpplmul_summul_n230) );
  AOI211_X1 SBOX_Inst_f1_phpplmul_summul_U42 ( .C1(SBOX_Inst_f1_phpplmul_sB[0]), .C2(SBOX_Inst_f1_phpplmul_sB[3]), .A(SBOX_Inst_f1_phpplmul_summul_n228), .B(
        SBOX_Inst_f1_phpplmul_summul_n291), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n229) );
  AND2_X1 SBOX_Inst_f1_phpplmul_summul_U41 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n296), .A2(
        SBOX_Inst_f1_phpplmul_summul_n292), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n228) );
  AOI211_X1 SBOX_Inst_f1_phpplmul_summul_U40 ( .C1(SBOX_Inst_f1_phpplmul_sA[0]), .C2(SBOX_Inst_f1_phpplmul_sA[2]), .A(SBOX_Inst_f1_phpplmul_summul_n298), .B(
        SBOX_Inst_f1_phpplmul_summul_n226), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n227) );
  AND2_X1 SBOX_Inst_f1_phpplmul_summul_U39 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n299), .A2(
        SBOX_Inst_f1_phpplmul_summul_n300), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n226) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U38 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n223), .B(
        SBOX_Inst_f1_phpplmul_summul_n224), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n225) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_summul_U37 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n295), .A2(
        SBOX_Inst_f1_phpplmul_summul_n294), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n224) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U36 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n293), .B(
        SBOX_Inst_f1_phpplmul_summul_n222), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n223) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U35 ( .A1(SBOX_Inst_f1_phpplmul_sA[1]), 
        .A2(SBOX_Inst_f1_phpplmul_summul_n296), .B1(
        SBOX_Inst_f1_phpplmul_sB[0]), .B2(SBOX_Inst_f1_phpplmul_summul_n297), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n222) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U34 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n221), .B(
        SBOX_Inst_f1_phpplmul_summul_n220), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_p[4]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U33 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n289), .B(
        SBOX_Inst_f1_phpplmul_summul_n217), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n221) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U32 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n218), .B(
        SBOX_Inst_f1_phpplmul_summul_n219), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n220) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_summul_U31 ( .A1(SBOX_Inst_f1_phpplmul_sB[3]), 
        .A2(SBOX_Inst_f1_phpplmul_summul_n294), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n219) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_summul_U30 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n300), .A2(
        SBOX_Inst_f1_phpplmul_summul_n290), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n218) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U29 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n293), .B(
        SBOX_Inst_f1_phpplmul_summul_n216), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n217) );
  MUX2_X1 SBOX_Inst_f1_phpplmul_summul_U28 ( .A(SBOX_Inst_f1_phpplmul_sB[0]), 
        .B(SBOX_Inst_f1_phpplmul_sB[1]), .S(SBOX_Inst_f1_phpplmul_summul_n215), 
        .Z(SBOX_Inst_f1_phpplmul_summul_n216) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U27 ( .A1(SBOX_Inst_f1_phpplmul_sA[3]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[1]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n294), .B2(
        SBOX_Inst_f1_phpplmul_summul_n291), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n215) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U26 ( .A1(SBOX_Inst_f1_phpplmul_sA[0]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[5]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n266) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_summul_U25 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n289), .B(
        SBOX_Inst_f1_phpplmul_summul_n273), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n269) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U24 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n246), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n245) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_summul_U23 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n246), .A2(
        SBOX_Inst_f1_phpplmul_summul_n276), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n248) );
  OAI21_X1 SBOX_Inst_f1_phpplmul_summul_U22 ( .B1(SBOX_Inst_f1_phpplmul_sB[4]), 
        .B2(SBOX_Inst_f1_phpplmul_summul_n235), .A(SBOX_Inst_f1_phpplmul_sA[3]), .ZN(SBOX_Inst_f1_phpplmul_summul_n234) );
  AOI21_X1 SBOX_Inst_f1_phpplmul_summul_U21 ( .B1(SBOX_Inst_f1_phpplmul_sB[4]), 
        .B2(SBOX_Inst_f1_phpplmul_summul_n235), .A(
        SBOX_Inst_f1_phpplmul_summul_n234), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n236) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_summul_U20 ( .B1(SBOX_Inst_f1_phpplmul_sA[3]), .B2(SBOX_Inst_f1_phpplmul_sA[5]), .C1(SBOX_Inst_f1_phpplmul_summul_n291), 
        .C2(SBOX_Inst_f1_phpplmul_summul_n276), .A(SBOX_Inst_f1_phpplmul_sB[2]), .ZN(SBOX_Inst_f1_phpplmul_summul_n239) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_summul_U19 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n278), .A2(SBOX_Inst_f1_phpplmul_sB[4]), 
        .B1(SBOX_Inst_f1_phpplmul_summul_n260), .B2(
        SBOX_Inst_f1_phpplmul_summul_n242), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n243) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U18 ( .A(SBOX_Inst_f1_phpplmul_sA[2]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n300) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U17 ( .A1(SBOX_Inst_f1_phpplmul_sA[0]), 
        .A2(SBOX_Inst_f1_phpplmul_sB[3]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n285) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U16 ( .A(SBOX_Inst_f1_phpplmul_sA[3]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n291) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U15 ( .A(SBOX_Inst_f1_phpplmul_sB[0]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n296) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U14 ( .A(SBOX_Inst_f1_phpplmul_sB[3]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n292) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U13 ( .A(SBOX_Inst_f1_phpplmul_sB[2]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n298) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U12 ( .A1(SBOX_Inst_f1_phpplmul_sA[2]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[0]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n299), .B2(
        SBOX_Inst_f1_phpplmul_summul_n300), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n297) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U11 ( .A(SBOX_Inst_f1_phpplmul_sA[0]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n299) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U10 ( .A(SBOX_Inst_f1_phpplmul_sB[1]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n295) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U9 ( .A(SBOX_Inst_f1_phpplmul_sB[5]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n260) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_summul_U8 ( .A1(SBOX_Inst_f1_phpplmul_sB[0]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[5]), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n258) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U7 ( .A(SBOX_Inst_f1_phpplmul_sB[4]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n259) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U6 ( .A(SBOX_Inst_f1_phpplmul_sA[4]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n252) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U5 ( .A(SBOX_Inst_f1_phpplmul_sA[5]), 
        .ZN(SBOX_Inst_f1_phpplmul_summul_n276) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_summul_U4 ( .A1(
        SBOX_Inst_f1_phpplmul_summul_n252), .A2(
        SBOX_Inst_f1_phpplmul_summul_n260), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n278) );
  INV_X1 SBOX_Inst_f1_phpplmul_summul_U3 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n282), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n281) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_summul_U2 ( .A1(SBOX_Inst_f1_phpplmul_sA[5]), 
        .A2(SBOX_Inst_f1_phpplmul_sA[0]), .B1(
        SBOX_Inst_f1_phpplmul_summul_n299), .B2(
        SBOX_Inst_f1_phpplmul_summul_n276), .ZN(
        SBOX_Inst_f1_phpplmul_summul_n282) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_summul_U1 ( .A(
        SBOX_Inst_f1_phpplmul_summul_n273), .B(
        SBOX_Inst_f1_phpplmul_summul_n272), .Z(
        SBOX_Inst_f1_phpplmul_summul_n275) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U8 ( .A(PRNGQ[7]), .B(
        SBOX_Inst_f1_phpplmul_Orig_p[3]), .Z(SBOX_p[3]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U7 ( .A(PRNGQ[6]), .B(
        SBOX_Inst_f1_phpplmul_Orig_p[2]), .Z(SBOX_p[2]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U6 ( .A(PRNGQ[5]), .B(
        SBOX_Inst_f1_phpplmul_Orig_p[1]), .Z(SBOX_p[1]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U5 ( .A(PRNGQ[4]), .B(
        SBOX_Inst_f1_phpplmul_Orig_p[0]), .Z(SBOX_p[0]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U4 ( .A(
        SBOX_Inst_f1_phpplmul_AddNewMaskp_n6), .B(PRNGQ[7]), .ZN(SBOX_p[5]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U3 ( .A(PRNGQ[5]), .B(
        SBOX_Inst_f1_phpplmul_Orig_p[5]), .ZN(
        SBOX_Inst_f1_phpplmul_AddNewMaskp_n6) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U2 ( .A(
        SBOX_Inst_f1_phpplmul_AddNewMaskp_n5), .B(PRNGQ[6]), .ZN(SBOX_p[4]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskp_U1 ( .A(PRNGQ[4]), .B(
        SBOX_Inst_f1_phpplmul_Orig_p[4]), .ZN(
        SBOX_Inst_f1_phpplmul_AddNewMaskp_n5) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U93 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n298), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n297), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_pl[4]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U92 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n296), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n295), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n297) );
  MUX2_X1 SBOX_Inst_f1_phpplmul_lowmul_U91 ( .A(SBOX_Zl_f1_0_), .B(
        SBOX_Zl_f1_1_), .S(SBOX_Inst_f1_phpplmul_lowmul_n294), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n295) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U90 ( .A1(SBOX_Zh_f1[1]), .A2(
        SBOX_Zh_f1[5]), .B1(SBOX_Inst_f1_phpplmul_lowmul_n293), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n292), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n294) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U89 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n291), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n290), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n296) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U88 ( .A1(SBOX_Zh_f1[4]), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n289), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n290) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U87 ( .A1(
        SBOX_Inst_f1_phpplmul_lowmul_n292), .A2(SBOX_Zl_f1_5_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n291) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U86 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n287), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n286), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n302) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U85 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n285), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n284), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n286) );
  AOI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U84 ( .B1(SBOX_Zl_f1_1_), .B2(
        SBOX_Zl_f1_5_), .C1(SBOX_Inst_f1_phpplmul_lowmul_n283), .C2(
        SBOX_Inst_f1_phpplmul_lowmul_n282), .A(
        SBOX_Inst_f1_phpplmul_lowmul_n299), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n287) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U83 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n281), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n280), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_pl[3]) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U82 ( .B1(SBOX_Zh_f1[1]), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n279), .C1(
        SBOX_Inst_f1_phpplmul_lowmul_n292), .C2(
        SBOX_Inst_f1_phpplmul_lowmul_n278), .A(SBOX_Zl_f1_8_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n280) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U81 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n277), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n276), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n281) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U80 ( .A1(SBOX_Zh_f1[8]), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n275), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n276) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U79 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n272), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n271), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n273) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U78 ( .A1(
        SBOX_Inst_f1_phpplmul_lowmul_n279), .A2(SBOX_Zl_f1_9_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n271) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U77 ( .A1(
        SBOX_Inst_f1_phpplmul_lowmul_n274), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n299), .B1(SBOX_Zh_f1[0]), .B2(
        SBOX_Zh_f1[9]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n278) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U76 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n268), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n267), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n269) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U75 ( .A1(SBOX_Zh_f1[8]), .A2(
        SBOX_Zl_f1_0_), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n268) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U74 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n266), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n265), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_pl[2]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U73 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n263), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n262), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n288) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U72 ( .A1(SBOX_Zl_f1_1_), .A2(
        SBOX_Zh_f1[0]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n262) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U71 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n261), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n260), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n264) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U70 ( .A1(SBOX_Zl_f1_0_), .A2(
        SBOX_Zh_f1[1]), .B1(SBOX_Inst_f1_phpplmul_lowmul_n292), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n259), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n260) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U69 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n257), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n256), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n270) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U68 ( .A1(SBOX_Zh_f1[8]), .A2(
        SBOX_Zl_f1_1_), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n257) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U67 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n255), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n254), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n258) );
  OAI21_X1 SBOX_Inst_f1_phpplmul_lowmul_U66 ( .B1(
        SBOX_Inst_f1_phpplmul_lowmul_n253), .B2(SBOX_Zl_f1_8_), .A(
        SBOX_Zh_f1[9]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n252) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U65 ( .A1(SBOX_Zl_f1_1_), .A2(
        SBOX_Zl_f1_9_), .B1(SBOX_Inst_f1_phpplmul_lowmul_n275), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n283), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n253) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U64 ( .A1(SBOX_Zh_f1[1]), .A2(
        SBOX_Zl_f1_9_), .B1(SBOX_Zl_f1_8_), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n292), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n255) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U63 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n251), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n250), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_pl[1]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U62 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n249), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n248), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n250) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U61 ( .B1(SBOX_Zl_f1_5_), .B2(
        SBOX_Zl_f1_4_), .C1(SBOX_Inst_f1_phpplmul_lowmul_n282), .C2(
        SBOX_Inst_f1_phpplmul_lowmul_n247), .A(SBOX_Zh_f1[5]), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n248) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U60 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n246), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n245), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n249) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U59 ( .B1(SBOX_Zh_f1[4]), .B2(
        SBOX_Zh_f1[5]), .C1(SBOX_Inst_f1_phpplmul_lowmul_n300), .C2(
        SBOX_Inst_f1_phpplmul_lowmul_n293), .A(SBOX_Zl_f1_8_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n245) );
  OAI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U58 ( .B1(SBOX_Zh_f1[8]), .B2(
        SBOX_Zh_f1[4]), .C1(SBOX_Inst_f1_phpplmul_lowmul_n244), .C2(
        SBOX_Inst_f1_phpplmul_lowmul_n300), .A(
        SBOX_Inst_f1_phpplmul_lowmul_n289), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n246) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U57 ( .A1(SBOX_Zl_f1_5_), .A2(
        SBOX_Zl_f1_4_), .B1(SBOX_Inst_f1_phpplmul_lowmul_n247), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n282), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n289) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U56 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n243), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n242), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n251) );
  AOI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U55 ( .B1(SBOX_Zh_f1[9]), .B2(
        SBOX_Zh_f1[4]), .C1(SBOX_Zl_f1_4_), .C2(SBOX_Zl_f1_9_), .A(
        SBOX_Inst_f1_phpplmul_lowmul_n237), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n243) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U54 ( .A1(SBOX_Zh_f1[9]), .A2(
        SBOX_Zh_f1[4]), .B1(SBOX_Zl_f1_9_), .B2(SBOX_Zl_f1_4_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n237) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U53 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n236), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n235), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_pl[0]) );
  OAI21_X1 SBOX_Inst_f1_phpplmul_lowmul_U52 ( .B1(SBOX_Zh_f1[8]), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n274), .A(
        SBOX_Inst_f1_phpplmul_lowmul_n240), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n239) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U51 ( .A1(SBOX_Zh_f1[8]), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n274), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n240) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U50 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n234), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n233), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n236) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U49 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n232), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n231), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n233) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U48 ( .A1(SBOX_Zh_f1[5]), .A2(
        SBOX_Zl_f1_9_), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n231) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U47 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n229), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n228), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n230) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U46 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n227), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n226), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n301) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U45 ( .A1(SBOX_Zh_f1[4]), .A2(
        SBOX_Zl_f1_4_), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n226) );
  AOI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U44 ( .B1(SBOX_Zh_f1[9]), .B2(
        SBOX_Zh_f1[5]), .C1(SBOX_Inst_f1_phpplmul_lowmul_n274), .C2(
        SBOX_Inst_f1_phpplmul_lowmul_n293), .A(
        SBOX_Inst_f1_phpplmul_lowmul_n247), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n234) );
  AOI221_X1 SBOX_Inst_f1_phpplmul_lowmul_U43 ( .B1(SBOX_Zh_f1[8]), .B2(
        SBOX_Zh_f1[4]), .C1(SBOX_Inst_f1_phpplmul_lowmul_n244), .C2(
        SBOX_Inst_f1_phpplmul_lowmul_n300), .A(
        SBOX_Inst_f1_phpplmul_lowmul_n275), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n228) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U42 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n302), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n225), .ZN(
        SBOX_Inst_f1_phpplmul_Orig_pl[5]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U41 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n218), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n224), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n225) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U40 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n223), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n222), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n224) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U39 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n221), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n301), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n223) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U38 ( .A1(SBOX_Zl_f1_0_), .A2(
        SBOX_Zh_f1[5]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n222) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U37 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n219), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n220), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n221) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U36 ( .A1(SBOX_Zl_f1_4_), .A2(
        SBOX_Zh_f1[0]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n220) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U35 ( .A1(SBOX_Zl_f1_1_), .A2(
        SBOX_Zh_f1[1]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n219) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U34 ( .A1(SBOX_Zl_f1_0_), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n216), .B1(SBOX_Zh_f1[1]), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n217), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n218) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U33 ( .A(SBOX_Zl_f1_0_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n217) );
  OAI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U32 ( .A1(SBOX_Zh_f1[0]), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n300), .B1(SBOX_Zh_f1[4]), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n299), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n216) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U31 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n288), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n302), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n298) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U30 ( .A1(SBOX_Zh_f1[1]), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n283), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n267) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U29 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n278), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n279) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U28 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n270), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n269), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n272) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U27 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n274), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n273), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n277) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U26 ( .A(SBOX_Zl_f1_0_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n259) );
  AOI21_X1 SBOX_Inst_f1_phpplmul_lowmul_U25 ( .B1(
        SBOX_Inst_f1_phpplmul_lowmul_n253), .B2(SBOX_Zl_f1_8_), .A(
        SBOX_Inst_f1_phpplmul_lowmul_n252), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n254) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U24 ( .A1(SBOX_Zh_f1[0]), .A2(
        SBOX_Zl_f1_9_), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n261) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U23 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n258), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n270), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n266) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U22 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n264), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n288), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n265) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U21 ( .A1(SBOX_Zh_f1[8]), .A2(
        SBOX_Zl_f1_8_), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n238) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U20 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n238), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n241) );
  AOI22_X1 SBOX_Inst_f1_phpplmul_lowmul_U19 ( .A1(
        SBOX_Inst_f1_phpplmul_lowmul_n241), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n240), .B1(
        SBOX_Inst_f1_phpplmul_lowmul_n239), .B2(
        SBOX_Inst_f1_phpplmul_lowmul_n238), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n242) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U18 ( .A1(
        SBOX_Inst_f1_phpplmul_lowmul_n293), .A2(SBOX_Zl_f1_8_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n229) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U17 ( .A(
        SBOX_Inst_f1_phpplmul_lowmul_n301), .B(
        SBOX_Inst_f1_phpplmul_lowmul_n230), .Z(
        SBOX_Inst_f1_phpplmul_lowmul_n232) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U16 ( .A1(SBOX_Zl_f1_5_), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n239), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n235) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U15 ( .A1(SBOX_Zl_f1_4_), .A2(
        SBOX_Zh_f1[1]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n285) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U14 ( .A1(SBOX_Zh_f1[4]), .A2(
        SBOX_Zl_f1_1_), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n284) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U13 ( .A(SBOX_Zh_f1[4]), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n300) );
  NOR2_X1 SBOX_Inst_f1_phpplmul_lowmul_U12 ( .A1(
        SBOX_Inst_f1_phpplmul_lowmul_n282), .A2(
        SBOX_Inst_f1_phpplmul_lowmul_n293), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n227) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U11 ( .A(SBOX_Zh_f1[0]), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n299) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U10 ( .A(SBOX_Zh_f1[1]), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n292) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U9 ( .A1(SBOX_Zl_f1_0_), .A2(
        SBOX_Zh_f1[1]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n263) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U8 ( .A(SBOX_Zh_f1[5]), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n293) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U7 ( .A(SBOX_Zh_f1[9]), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n274) );
  NAND2_X1 SBOX_Inst_f1_phpplmul_lowmul_U6 ( .A1(SBOX_Zl_f1_0_), .A2(
        SBOX_Zh_f1[9]), .ZN(SBOX_Inst_f1_phpplmul_lowmul_n256) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U5 ( .A(SBOX_Zl_f1_9_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n275) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U4 ( .A(SBOX_Zl_f1_1_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n283) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U3 ( .A(SBOX_Zl_f1_4_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n247) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U2 ( .A(SBOX_Zl_f1_5_), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n282) );
  INV_X1 SBOX_Inst_f1_phpplmul_lowmul_U1 ( .A(SBOX_Zh_f1[8]), .ZN(
        SBOX_Inst_f1_phpplmul_lowmul_n244) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U8 ( .A(PRNGQ[8]), .B(
        SBOX_Inst_f1_phpplmul_Orig_pl[4]), .ZN(
        SBOX_Inst_f1_phpplmul_AddNewMaskpl_n6) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U7 ( .A(PRNGQ[11]), .B(
        SBOX_Inst_f1_phpplmul_Orig_pl[3]), .Z(SBOX_pl[3]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U6 ( .A(PRNGQ[10]), .B(
        SBOX_Inst_f1_phpplmul_Orig_pl[2]), .Z(SBOX_pl[2]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U5 ( .A(PRNGQ[9]), .B(
        SBOX_Inst_f1_phpplmul_Orig_pl[1]), .Z(SBOX_pl[1]) );
  XOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U4 ( .A(PRNGQ[8]), .B(
        SBOX_Inst_f1_phpplmul_Orig_pl[0]), .Z(SBOX_pl[0]) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U3 ( .A(
        SBOX_Inst_f1_phpplmul_AddNewMaskpl_n5), .B(PRNGQ[11]), .ZN(SBOX_pl[5])
         );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U2 ( .A(PRNGQ[9]), .B(
        SBOX_Inst_f1_phpplmul_Orig_pl[5]), .ZN(
        SBOX_Inst_f1_phpplmul_AddNewMaskpl_n5) );
  XNOR2_X1 SBOX_Inst_f1_phpplmul_AddNewMaskpl_U1 ( .A(
        SBOX_Inst_f1_phpplmul_AddNewMaskpl_n6), .B(PRNGQ[10]), .ZN(SBOX_pl[4])
         );
  OAI21_X1 SBOX_PL_1_U109 ( .B1(1'b1), .B2(SBOX_PL_1_n107), .A(SBOX_PL_1_n54), 
        .ZN(SBOX_PL_1_n161) );
  NAND2_X1 SBOX_PL_1_U108 ( .A1(1'b1), .A2(SBOX_Zh_f1[10]), .ZN(SBOX_PL_1_n54)
         );
  OAI21_X1 SBOX_PL_1_U107 ( .B1(1'b1), .B2(SBOX_PL_1_n101), .A(SBOX_PL_1_n53), 
        .ZN(SBOX_PL_1_n155) );
  NAND2_X1 SBOX_PL_1_U106 ( .A1(1'b1), .A2(SBOX_Zh_f1[4]), .ZN(SBOX_PL_1_n53)
         );
  OAI21_X1 SBOX_PL_1_U105 ( .B1(1'b1), .B2(SBOX_PL_1_n100), .A(SBOX_PL_1_n52), 
        .ZN(SBOX_PL_1_n154) );
  NAND2_X1 SBOX_PL_1_U104 ( .A1(1'b1), .A2(SBOX_Zh_f1[3]), .ZN(SBOX_PL_1_n52)
         );
  OAI21_X1 SBOX_PL_1_U103 ( .B1(1'b1), .B2(SBOX_PL_1_n99), .A(SBOX_PL_1_n51), 
        .ZN(SBOX_PL_1_n153) );
  NAND2_X1 SBOX_PL_1_U102 ( .A1(1'b1), .A2(SBOX_Zh_f1[2]), .ZN(SBOX_PL_1_n51)
         );
  OAI21_X1 SBOX_PL_1_U101 ( .B1(1'b1), .B2(SBOX_PL_1_n98), .A(SBOX_PL_1_n50), 
        .ZN(SBOX_PL_1_n152) );
  NAND2_X1 SBOX_PL_1_U100 ( .A1(1'b1), .A2(SBOX_Zh_f1[1]), .ZN(SBOX_PL_1_n50)
         );
  OAI21_X1 SBOX_PL_1_U99 ( .B1(1'b1), .B2(SBOX_PL_1_n96), .A(SBOX_PL_1_n49), 
        .ZN(SBOX_PL_1_n150) );
  NAND2_X1 SBOX_PL_1_U98 ( .A1(1'b1), .A2(SBOX_Zl_f1_11_), .ZN(SBOX_PL_1_n49)
         );
  OAI21_X1 SBOX_PL_1_U97 ( .B1(1'b1), .B2(SBOX_PL_1_n89), .A(SBOX_PL_1_n48), 
        .ZN(SBOX_PL_1_n143) );
  NAND2_X1 SBOX_PL_1_U96 ( .A1(1'b1), .A2(SBOX_Zl_f1_4_), .ZN(SBOX_PL_1_n48)
         );
  OAI21_X1 SBOX_PL_1_U95 ( .B1(1'b1), .B2(SBOX_PL_1_n86), .A(SBOX_PL_1_n47), 
        .ZN(SBOX_PL_1_n140) );
  NAND2_X1 SBOX_PL_1_U94 ( .A1(1'b1), .A2(SBOX_Zl_f1_1_), .ZN(SBOX_PL_1_n47)
         );
  OAI21_X1 SBOX_PL_1_U93 ( .B1(1'b1), .B2(SBOX_PL_1_n85), .A(SBOX_PL_1_n46), 
        .ZN(SBOX_PL_1_n139) );
  NAND2_X1 SBOX_PL_1_U92 ( .A1(1'b1), .A2(SBOX_Zl_f1_0_), .ZN(SBOX_PL_1_n46)
         );
  OAI21_X1 SBOX_PL_1_U91 ( .B1(1'b1), .B2(SBOX_PL_1_n64), .A(SBOX_PL_1_n45), 
        .ZN(SBOX_PL_1_n118) );
  NAND2_X1 SBOX_PL_1_U90 ( .A1(1'b1), .A2(SBOX_p[3]), .ZN(SBOX_PL_1_n45) );
  OAI21_X1 SBOX_PL_1_U89 ( .B1(1'b1), .B2(SBOX_PL_1_n63), .A(SBOX_PL_1_n44), 
        .ZN(SBOX_PL_1_n117) );
  NAND2_X1 SBOX_PL_1_U88 ( .A1(1'b1), .A2(SBOX_p[2]), .ZN(SBOX_PL_1_n44) );
  OAI21_X1 SBOX_PL_1_U87 ( .B1(1'b1), .B2(SBOX_PL_1_n62), .A(SBOX_PL_1_n43), 
        .ZN(SBOX_PL_1_n116) );
  NAND2_X1 SBOX_PL_1_U86 ( .A1(1'b1), .A2(SBOX_p[1]), .ZN(SBOX_PL_1_n43) );
  OAI21_X1 SBOX_PL_1_U85 ( .B1(1'b1), .B2(SBOX_PL_1_n61), .A(SBOX_PL_1_n42), 
        .ZN(SBOX_PL_1_n115) );
  NAND2_X1 SBOX_PL_1_U84 ( .A1(1'b1), .A2(SBOX_p[0]), .ZN(SBOX_PL_1_n42) );
  OAI21_X1 SBOX_PL_1_U83 ( .B1(1'b1), .B2(SBOX_PL_1_n59), .A(SBOX_PL_1_n41), 
        .ZN(SBOX_PL_1_n113) );
  NAND2_X1 SBOX_PL_1_U82 ( .A1(1'b1), .A2(SBOX_pl[4]), .ZN(SBOX_PL_1_n41) );
  OAI21_X1 SBOX_PL_1_U81 ( .B1(1'b1), .B2(SBOX_PL_1_n58), .A(SBOX_PL_1_n40), 
        .ZN(SBOX_PL_1_n112) );
  NAND2_X1 SBOX_PL_1_U80 ( .A1(1'b1), .A2(SBOX_pl[3]), .ZN(SBOX_PL_1_n40) );
  OAI21_X1 SBOX_PL_1_U79 ( .B1(1'b1), .B2(SBOX_PL_1_n57), .A(SBOX_PL_1_n39), 
        .ZN(SBOX_PL_1_n111) );
  NAND2_X1 SBOX_PL_1_U78 ( .A1(1'b1), .A2(SBOX_pl[2]), .ZN(SBOX_PL_1_n39) );
  OAI21_X1 SBOX_PL_1_U77 ( .B1(1'b1), .B2(SBOX_PL_1_n56), .A(SBOX_PL_1_n38), 
        .ZN(SBOX_PL_1_n110) );
  NAND2_X1 SBOX_PL_1_U76 ( .A1(1'b1), .A2(SBOX_pl[1]), .ZN(SBOX_PL_1_n38) );
  OAI21_X1 SBOX_PL_1_U75 ( .B1(1'b1), .B2(SBOX_PL_1_n55), .A(SBOX_PL_1_n37), 
        .ZN(SBOX_PL_1_n109) );
  NAND2_X1 SBOX_PL_1_U74 ( .A1(1'b1), .A2(SBOX_pl[0]), .ZN(SBOX_PL_1_n37) );
  OAI21_X1 SBOX_PL_1_U73 ( .B1(1'b1), .B2(SBOX_PL_1_n108), .A(SBOX_PL_1_n36), 
        .ZN(SBOX_PL_1_n162) );
  NAND2_X1 SBOX_PL_1_U72 ( .A1(1'b1), .A2(SBOX_Zh_f1[11]), .ZN(SBOX_PL_1_n36)
         );
  OAI21_X1 SBOX_PL_1_U71 ( .B1(1'b1), .B2(SBOX_PL_1_n106), .A(SBOX_PL_1_n35), 
        .ZN(SBOX_PL_1_n160) );
  NAND2_X1 SBOX_PL_1_U70 ( .A1(1'b1), .A2(SBOX_Zh_f1[9]), .ZN(SBOX_PL_1_n35)
         );
  OAI21_X1 SBOX_PL_1_U69 ( .B1(1'b1), .B2(SBOX_PL_1_n104), .A(SBOX_PL_1_n34), 
        .ZN(SBOX_PL_1_n158) );
  NAND2_X1 SBOX_PL_1_U68 ( .A1(1'b1), .A2(SBOX_Zh_f1[7]), .ZN(SBOX_PL_1_n34)
         );
  OAI21_X1 SBOX_PL_1_U67 ( .B1(1'b1), .B2(SBOX_PL_1_n103), .A(SBOX_PL_1_n33), 
        .ZN(SBOX_PL_1_n157) );
  NAND2_X1 SBOX_PL_1_U66 ( .A1(1'b1), .A2(SBOX_Zh_f1[6]), .ZN(SBOX_PL_1_n33)
         );
  OAI21_X1 SBOX_PL_1_U65 ( .B1(1'b1), .B2(SBOX_PL_1_n97), .A(SBOX_PL_1_n32), 
        .ZN(SBOX_PL_1_n151) );
  NAND2_X1 SBOX_PL_1_U64 ( .A1(1'b1), .A2(SBOX_Zh_f1[0]), .ZN(SBOX_PL_1_n32)
         );
  OAI21_X1 SBOX_PL_1_U63 ( .B1(1'b1), .B2(SBOX_PL_1_n95), .A(SBOX_PL_1_n31), 
        .ZN(SBOX_PL_1_n149) );
  NAND2_X1 SBOX_PL_1_U62 ( .A1(1'b1), .A2(CxDO[16]), .ZN(SBOX_PL_1_n31) );
  OAI21_X1 SBOX_PL_1_U61 ( .B1(1'b1), .B2(SBOX_PL_1_n92), .A(SBOX_PL_1_n30), 
        .ZN(SBOX_PL_1_n146) );
  NAND2_X1 SBOX_PL_1_U60 ( .A1(1'b1), .A2(SBOX_Zl_f1_7_), .ZN(SBOX_PL_1_n30)
         );
  OAI21_X1 SBOX_PL_1_U59 ( .B1(1'b1), .B2(SBOX_PL_1_n91), .A(SBOX_PL_1_n29), 
        .ZN(SBOX_PL_1_n145) );
  NAND2_X1 SBOX_PL_1_U58 ( .A1(1'b1), .A2(CxDO[8]), .ZN(SBOX_PL_1_n29) );
  OAI21_X1 SBOX_PL_1_U57 ( .B1(1'b1), .B2(SBOX_PL_1_n88), .A(SBOX_PL_1_n28), 
        .ZN(SBOX_PL_1_n142) );
  NAND2_X1 SBOX_PL_1_U56 ( .A1(1'b1), .A2(SBOX_Zl_f1_3_), .ZN(SBOX_PL_1_n28)
         );
  OAI21_X1 SBOX_PL_1_U55 ( .B1(1'b1), .B2(SBOX_PL_1_n87), .A(SBOX_PL_1_n27), 
        .ZN(SBOX_PL_1_n141) );
  NAND2_X1 SBOX_PL_1_U54 ( .A1(1'b1), .A2(CxDO[0]), .ZN(SBOX_PL_1_n27) );
  OAI21_X1 SBOX_PL_1_U53 ( .B1(1'b1), .B2(SBOX_PL_1_n81), .A(SBOX_PL_1_n26), 
        .ZN(SBOX_PL_1_n135) );
  NAND2_X1 SBOX_PL_1_U52 ( .A1(1'b1), .A2(SBOX_ab2[8]), .ZN(SBOX_PL_1_n26) );
  OAI21_X1 SBOX_PL_1_U51 ( .B1(1'b1), .B2(SBOX_PL_1_n77), .A(SBOX_PL_1_n25), 
        .ZN(SBOX_PL_1_n131) );
  NAND2_X1 SBOX_PL_1_U50 ( .A1(1'b1), .A2(SBOX_ab2[4]), .ZN(SBOX_PL_1_n25) );
  OAI21_X1 SBOX_PL_1_U49 ( .B1(1'b1), .B2(SBOX_PL_1_n105), .A(SBOX_PL_1_n24), 
        .ZN(SBOX_PL_1_n159) );
  NAND2_X1 SBOX_PL_1_U48 ( .A1(1'b1), .A2(SBOX_Zh_f1[8]), .ZN(SBOX_PL_1_n24)
         );
  OAI21_X1 SBOX_PL_1_U47 ( .B1(1'b1), .B2(SBOX_PL_1_n102), .A(SBOX_PL_1_n23), 
        .ZN(SBOX_PL_1_n156) );
  NAND2_X1 SBOX_PL_1_U46 ( .A1(1'b1), .A2(SBOX_Zh_f1[5]), .ZN(SBOX_PL_1_n23)
         );
  OAI21_X1 SBOX_PL_1_U45 ( .B1(1'b1), .B2(SBOX_PL_1_n93), .A(SBOX_PL_1_n22), 
        .ZN(SBOX_PL_1_n147) );
  NAND2_X1 SBOX_PL_1_U44 ( .A1(1'b1), .A2(SBOX_Zl_f1_8_), .ZN(SBOX_PL_1_n22)
         );
  OAI21_X1 SBOX_PL_1_U43 ( .B1(1'b1), .B2(SBOX_PL_1_n76), .A(SBOX_PL_1_n21), 
        .ZN(SBOX_PL_1_n130) );
  NAND2_X1 SBOX_PL_1_U42 ( .A1(1'b1), .A2(SBOX_ab2[3]), .ZN(SBOX_PL_1_n21) );
  OAI21_X1 SBOX_PL_1_U41 ( .B1(1'b1), .B2(SBOX_PL_1_n90), .A(SBOX_PL_1_n20), 
        .ZN(SBOX_PL_1_n144) );
  NAND2_X1 SBOX_PL_1_U40 ( .A1(1'b1), .A2(SBOX_Zl_f1_5_), .ZN(SBOX_PL_1_n20)
         );
  OAI21_X1 SBOX_PL_1_U39 ( .B1(1'b1), .B2(SBOX_PL_1_n84), .A(SBOX_PL_1_n19), 
        .ZN(SBOX_PL_1_n138) );
  NAND2_X1 SBOX_PL_1_U38 ( .A1(1'b1), .A2(SBOX_ab2[11]), .ZN(SBOX_PL_1_n19) );
  OAI21_X1 SBOX_PL_1_U37 ( .B1(1'b1), .B2(SBOX_PL_1_n75), .A(SBOX_PL_1_n18), 
        .ZN(SBOX_PL_1_n129) );
  NAND2_X1 SBOX_PL_1_U36 ( .A1(1'b1), .A2(SBOX_ab2[2]), .ZN(SBOX_PL_1_n18) );
  OAI21_X1 SBOX_PL_1_U35 ( .B1(1'b1), .B2(SBOX_PL_1_n73), .A(SBOX_PL_1_n17), 
        .ZN(SBOX_PL_1_n127) );
  NAND2_X1 SBOX_PL_1_U34 ( .A1(1'b1), .A2(SBOX_ab2[0]), .ZN(SBOX_PL_1_n17) );
  OAI21_X1 SBOX_PL_1_U33 ( .B1(1'b1), .B2(SBOX_PL_1_n94), .A(SBOX_PL_1_n16), 
        .ZN(SBOX_PL_1_n148) );
  NAND2_X1 SBOX_PL_1_U32 ( .A1(1'b1), .A2(SBOX_Zl_f1_9_), .ZN(SBOX_PL_1_n16)
         );
  OAI21_X1 SBOX_PL_1_U31 ( .B1(1'b1), .B2(SBOX_PL_1_n80), .A(SBOX_PL_1_n15), 
        .ZN(SBOX_PL_1_n134) );
  NAND2_X1 SBOX_PL_1_U30 ( .A1(1'b1), .A2(SBOX_ab2[7]), .ZN(SBOX_PL_1_n15) );
  OAI21_X1 SBOX_PL_1_U29 ( .B1(1'b1), .B2(SBOX_PL_1_n74), .A(SBOX_PL_1_n14), 
        .ZN(SBOX_PL_1_n128) );
  NAND2_X1 SBOX_PL_1_U28 ( .A1(1'b1), .A2(SBOX_ab2[1]), .ZN(SBOX_PL_1_n14) );
  OAI21_X1 SBOX_PL_1_U27 ( .B1(1'b1), .B2(SBOX_PL_1_n83), .A(SBOX_PL_1_n13), 
        .ZN(SBOX_PL_1_n137) );
  NAND2_X1 SBOX_PL_1_U26 ( .A1(1'b1), .A2(SBOX_ab2[10]), .ZN(SBOX_PL_1_n13) );
  OAI21_X1 SBOX_PL_1_U25 ( .B1(1'b1), .B2(SBOX_PL_1_n79), .A(SBOX_PL_1_n12), 
        .ZN(SBOX_PL_1_n133) );
  NAND2_X1 SBOX_PL_1_U24 ( .A1(1'b1), .A2(SBOX_ab2[6]), .ZN(SBOX_PL_1_n12) );
  OAI21_X1 SBOX_PL_1_U23 ( .B1(1'b1), .B2(SBOX_PL_1_n82), .A(SBOX_PL_1_n11), 
        .ZN(SBOX_PL_1_n136) );
  NAND2_X1 SBOX_PL_1_U22 ( .A1(1'b1), .A2(SBOX_ab2[9]), .ZN(SBOX_PL_1_n11) );
  OAI21_X1 SBOX_PL_1_U21 ( .B1(1'b1), .B2(SBOX_PL_1_n78), .A(SBOX_PL_1_n10), 
        .ZN(SBOX_PL_1_n132) );
  NAND2_X1 SBOX_PL_1_U20 ( .A1(1'b1), .A2(SBOX_ab2[5]), .ZN(SBOX_PL_1_n10) );
  OAI21_X1 SBOX_PL_1_U19 ( .B1(1'b1), .B2(SBOX_PL_1_n71), .A(SBOX_PL_1_n9), 
        .ZN(SBOX_PL_1_n125) );
  NAND2_X1 SBOX_PL_1_U18 ( .A1(1'b1), .A2(SBOX_ph[4]), .ZN(SBOX_PL_1_n9) );
  OAI21_X1 SBOX_PL_1_U17 ( .B1(1'b1), .B2(SBOX_PL_1_n60), .A(SBOX_PL_1_n8), 
        .ZN(SBOX_PL_1_n114) );
  NAND2_X1 SBOX_PL_1_U16 ( .A1(1'b1), .A2(SBOX_pl[5]), .ZN(SBOX_PL_1_n8) );
  OAI21_X1 SBOX_PL_1_U15 ( .B1(1'b1), .B2(SBOX_PL_1_n72), .A(SBOX_PL_1_n7), 
        .ZN(SBOX_PL_1_n126) );
  NAND2_X1 SBOX_PL_1_U14 ( .A1(1'b1), .A2(SBOX_ph[5]), .ZN(SBOX_PL_1_n7) );
  OAI21_X1 SBOX_PL_1_U13 ( .B1(1'b1), .B2(SBOX_PL_1_n70), .A(SBOX_PL_1_n6), 
        .ZN(SBOX_PL_1_n124) );
  NAND2_X1 SBOX_PL_1_U12 ( .A1(1'b1), .A2(SBOX_ph[3]), .ZN(SBOX_PL_1_n6) );
  OAI21_X1 SBOX_PL_1_U11 ( .B1(1'b1), .B2(SBOX_PL_1_n69), .A(SBOX_PL_1_n5), 
        .ZN(SBOX_PL_1_n123) );
  NAND2_X1 SBOX_PL_1_U10 ( .A1(1'b1), .A2(SBOX_ph[2]), .ZN(SBOX_PL_1_n5) );
  OAI21_X1 SBOX_PL_1_U9 ( .B1(1'b1), .B2(SBOX_PL_1_n68), .A(SBOX_PL_1_n4), 
        .ZN(SBOX_PL_1_n122) );
  NAND2_X1 SBOX_PL_1_U8 ( .A1(1'b1), .A2(SBOX_ph[1]), .ZN(SBOX_PL_1_n4) );
  OAI21_X1 SBOX_PL_1_U7 ( .B1(1'b1), .B2(SBOX_PL_1_n67), .A(SBOX_PL_1_n3), 
        .ZN(SBOX_PL_1_n121) );
  NAND2_X1 SBOX_PL_1_U6 ( .A1(1'b1), .A2(SBOX_ph[0]), .ZN(SBOX_PL_1_n3) );
  OAI21_X1 SBOX_PL_1_U5 ( .B1(1'b1), .B2(SBOX_PL_1_n66), .A(SBOX_PL_1_n2), 
        .ZN(SBOX_PL_1_n120) );
  NAND2_X1 SBOX_PL_1_U4 ( .A1(1'b1), .A2(SBOX_p[5]), .ZN(SBOX_PL_1_n2) );
  OAI21_X1 SBOX_PL_1_U3 ( .B1(1'b1), .B2(SBOX_PL_1_n65), .A(SBOX_PL_1_n1), 
        .ZN(SBOX_PL_1_n119) );
  NAND2_X1 SBOX_PL_1_U2 ( .A1(1'b1), .A2(SBOX_p[4]), .ZN(SBOX_PL_1_n1) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_0_ ( .D(SBOX_PL_1_n109), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[0]), .QN(SBOX_PL_1_n55) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_1_ ( .D(SBOX_PL_1_n110), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[1]), .QN(SBOX_PL_1_n56) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_2_ ( .D(SBOX_PL_1_n111), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[2]), .QN(SBOX_PL_1_n57) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_3_ ( .D(SBOX_PL_1_n112), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[3]), .QN(SBOX_PL_1_n58) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_4_ ( .D(SBOX_PL_1_n113), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[4]), .QN(SBOX_PL_1_n59) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_5_ ( .D(SBOX_PL_1_n114), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[5]), .QN(SBOX_PL_1_n60) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_6_ ( .D(SBOX_PL_1_n115), .CK(ClkxCI), 
        .Q(SBOX_Inst_f2_abmul_pw2_1_), .QN(SBOX_PL_1_n61) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_7_ ( .D(SBOX_PL_1_n116), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[7]), .QN(SBOX_PL_1_n62) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_8_ ( .D(SBOX_PL_1_n117), .CK(ClkxCI), 
        .Q(SBOX_Inst_f2_abmul_pw2_3_), .QN(SBOX_PL_1_n63) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_9_ ( .D(SBOX_PL_1_n118), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[9]), .QN(SBOX_PL_1_n64) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_10_ ( .D(SBOX_PL_1_n119), .CK(ClkxCI), 
        .Q(SBOX_Inst_f2_abmul_pw2_5_), .QN(SBOX_PL_1_n65) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_11_ ( .D(SBOX_PL_1_n120), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[11]), .QN(SBOX_PL_1_n66) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_12_ ( .D(SBOX_PL_1_n121), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[12]), .QN(SBOX_PL_1_n67) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_13_ ( .D(SBOX_PL_1_n122), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[13]), .QN(SBOX_PL_1_n68) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_14_ ( .D(SBOX_PL_1_n123), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[14]), .QN(SBOX_PL_1_n69) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_15_ ( .D(SBOX_PL_1_n124), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[15]), .QN(SBOX_PL_1_n70) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_16_ ( .D(SBOX_PL_1_n125), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[16]), .QN(SBOX_PL_1_n71) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_17_ ( .D(SBOX_PL_1_n126), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[17]), .QN(SBOX_PL_1_n72) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_18_ ( .D(SBOX_PL_1_n127), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[18]), .QN(SBOX_PL_1_n73) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_19_ ( .D(SBOX_PL_1_n128), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[19]), .QN(SBOX_PL_1_n74) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_20_ ( .D(SBOX_PL_1_n129), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[20]), .QN(SBOX_PL_1_n75) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_21_ ( .D(SBOX_PL_1_n130), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[21]), .QN(SBOX_PL_1_n76) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_22_ ( .D(SBOX_PL_1_n131), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[22]), .QN(SBOX_PL_1_n77) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_23_ ( .D(SBOX_PL_1_n132), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[23]), .QN(SBOX_PL_1_n78) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_24_ ( .D(SBOX_PL_1_n133), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[24]), .QN(SBOX_PL_1_n79) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_25_ ( .D(SBOX_PL_1_n134), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[25]), .QN(SBOX_PL_1_n80) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_26_ ( .D(SBOX_PL_1_n135), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[26]), .QN(SBOX_PL_1_n81) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_27_ ( .D(SBOX_PL_1_n136), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[27]), .QN(SBOX_PL_1_n82) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_28_ ( .D(SBOX_PL_1_n137), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[28]), .QN(SBOX_PL_1_n83) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_29_ ( .D(SBOX_PL_1_n138), .CK(ClkxCI), 
        .Q(SBOX_FF1_out[29]), .QN(SBOX_PL_1_n84) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_30_ ( .D(SBOX_PL_1_n139), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[0]), .QN(SBOX_PL_1_n85) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_31_ ( .D(SBOX_PL_1_n140), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[1]), .QN(SBOX_PL_1_n86) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_32_ ( .D(SBOX_PL_1_n141), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[2]), .QN(SBOX_PL_1_n87) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_33_ ( .D(SBOX_PL_1_n142), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[3]), .QN(SBOX_PL_1_n88) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_34_ ( .D(SBOX_PL_1_n143), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[4]), .QN(SBOX_PL_1_n89) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_35_ ( .D(SBOX_PL_1_n144), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[5]), .QN(SBOX_PL_1_n90) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_36_ ( .D(SBOX_PL_1_n145), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[6]), .QN(SBOX_PL_1_n91) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_37_ ( .D(SBOX_PL_1_n146), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[7]), .QN(SBOX_PL_1_n92) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_38_ ( .D(SBOX_PL_1_n147), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[8]), .QN(SBOX_PL_1_n93) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_39_ ( .D(SBOX_PL_1_n148), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[9]), .QN(SBOX_PL_1_n94) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_40_ ( .D(SBOX_PL_1_n149), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[10]), .QN(SBOX_PL_1_n95) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_41_ ( .D(SBOX_PL_1_n150), .CK(ClkxCI), 
        .Q(SBOX_Zl_f2[11]), .QN(SBOX_PL_1_n96) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_42_ ( .D(SBOX_PL_1_n151), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[0]), .QN(SBOX_PL_1_n97) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_43_ ( .D(SBOX_PL_1_n152), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[1]), .QN(SBOX_PL_1_n98) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_44_ ( .D(SBOX_PL_1_n153), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[2]), .QN(SBOX_PL_1_n99) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_45_ ( .D(SBOX_PL_1_n154), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[3]), .QN(SBOX_PL_1_n100) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_46_ ( .D(SBOX_PL_1_n155), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[4]), .QN(SBOX_PL_1_n101) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_47_ ( .D(SBOX_PL_1_n156), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[5]), .QN(SBOX_PL_1_n102) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_48_ ( .D(SBOX_PL_1_n157), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[6]), .QN(SBOX_PL_1_n103) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_49_ ( .D(SBOX_PL_1_n158), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[7]), .QN(SBOX_PL_1_n104) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_50_ ( .D(SBOX_PL_1_n159), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[8]), .QN(SBOX_PL_1_n105) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_51_ ( .D(SBOX_PL_1_n160), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[9]), .QN(SBOX_PL_1_n106) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_52_ ( .D(SBOX_PL_1_n161), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[10]), .QN(SBOX_PL_1_n107) );
  DFF_X1 SBOX_PL_1_s_current_state_reg_53_ ( .D(SBOX_PL_1_n162), .CK(ClkxCI), 
        .Q(SBOX_Zh_f2[11]), .QN(SBOX_PL_1_n108) );
  XOR2_X2 SBOX_Inst_f2_U12 ( .A(SBOX_FF1_out[26]), .B(SBOX_Inst_f2_abin[8]), 
        .Z(SBOX_gamma0[4]) );
  XOR2_X2 SBOX_Inst_f2_U11 ( .A(SBOX_FF1_out[28]), .B(SBOX_Inst_f2_abin[10]), 
        .Z(SBOX_gamma1[4]) );
  XOR2_X2 SBOX_Inst_f2_U10 ( .A(SBOX_FF1_out[21]), .B(SBOX_Inst_f2_abin[3]), 
        .Z(SBOX_gamma1[1]) );
  XOR2_X1 SBOX_Inst_f2_U9 ( .A(SBOX_FF1_out[18]), .B(SBOX_Inst_f2_abin[0]), 
        .Z(SBOX_gamma0[0]) );
  XOR2_X1 SBOX_Inst_f2_U8 ( .A(SBOX_FF1_out[24]), .B(SBOX_Inst_f2_abin[6]), 
        .Z(SBOX_gamma1[2]) );
  XOR2_X1 SBOX_Inst_f2_U7 ( .A(SBOX_FF1_out[19]), .B(SBOX_Inst_f2_abin[1]), 
        .Z(SBOX_gamma0[1]) );
  XOR2_X1 SBOX_Inst_f2_U6 ( .A(SBOX_FF1_out[29]), .B(SBOX_Inst_f2_abin[11]), 
        .Z(SBOX_gamma1[5]) );
  XOR2_X1 SBOX_Inst_f2_U5 ( .A(SBOX_FF1_out[27]), .B(SBOX_Inst_f2_abin[9]), 
        .Z(SBOX_gamma0[5]) );
  XOR2_X1 SBOX_Inst_f2_U4 ( .A(SBOX_FF1_out[25]), .B(SBOX_Inst_f2_abin[7]), 
        .Z(SBOX_gamma1[3]) );
  XOR2_X1 SBOX_Inst_f2_U3 ( .A(SBOX_FF1_out[22]), .B(SBOX_Inst_f2_abin[4]), 
        .Z(SBOX_gamma0[2]) );
  XOR2_X1 SBOX_Inst_f2_U2 ( .A(SBOX_FF1_out[20]), .B(SBOX_Inst_f2_abin[2]), 
        .Z(SBOX_gamma1[0]) );
  XOR2_X1 SBOX_Inst_f2_U1 ( .A(SBOX_FF1_out[23]), .B(SBOX_Inst_f2_abin[5]), 
        .Z(SBOX_gamma0[3]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U12 ( .A(SBOX_Inst_f2_abmul_pw2_0_), .B(
        SBOX_FF1_out[0]), .Z(SBOX_Inst_f2_abin[0]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U11 ( .A(SBOX_Inst_f2_abmul_pw2_2_), .B(
        SBOX_FF1_out[14]), .Z(SBOX_Inst_f2_abin[6]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U10 ( .A(SBOX_Inst_f2_abmul_pw2_1_), .B(
        SBOX_FF1_out[1]), .Z(SBOX_Inst_f2_abin[1]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U9 ( .A(SBOX_Inst_f2_abmul_pw2_5_), .B(
        SBOX_FF1_out[17]), .Z(SBOX_Inst_f2_abin[11]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U8 ( .A(SBOX_Inst_f2_abmul_pw2_5_), .B(
        SBOX_FF1_out[5]), .Z(SBOX_Inst_f2_abin[9]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U7 ( .A(SBOX_Inst_f2_abmul_pw2_3_), .B(
        SBOX_FF1_out[15]), .Z(SBOX_Inst_f2_abin[7]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U6 ( .A(SBOX_Inst_f2_abmul_pw2_2_), .B(
        SBOX_FF1_out[2]), .Z(SBOX_Inst_f2_abin[4]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U5 ( .A(SBOX_Inst_f2_abmul_pw2_0_), .B(
        SBOX_FF1_out[12]), .Z(SBOX_Inst_f2_abin[2]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U4 ( .A(SBOX_Inst_f2_abmul_pw2_3_), .B(
        SBOX_FF1_out[3]), .Z(SBOX_Inst_f2_abin[5]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U3 ( .A(SBOX_Inst_f2_abmul_pw2_4_), .B(
        SBOX_FF1_out[16]), .Z(SBOX_Inst_f2_abin[10]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U2 ( .A(SBOX_Inst_f2_abmul_pw2_1_), .B(
        SBOX_FF1_out[13]), .Z(SBOX_Inst_f2_abin[3]) );
  XOR2_X1 SBOX_Inst_f2_abmul_U1 ( .A(SBOX_Inst_f2_abmul_pw2_4_), .B(
        SBOX_FF1_out[4]), .Z(SBOX_Inst_f2_abin[8]) );
  XOR2_X1 SBOX_Inst_f2_abmul_NxGAMMA_U3 ( .A(SBOX_Inst_f2_abmul_pw2_5_), .B(
        SBOX_FF1_out[11]), .Z(SBOX_Inst_f2_abmul_pw2_4_) );
  XOR2_X1 SBOX_Inst_f2_abmul_NxGAMMA_U2 ( .A(SBOX_Inst_f2_abmul_pw2_3_), .B(
        SBOX_FF1_out[9]), .Z(SBOX_Inst_f2_abmul_pw2_2_) );
  XOR2_X1 SBOX_Inst_f2_abmul_NxGAMMA_U1 ( .A(SBOX_Inst_f2_abmul_pw2_1_), .B(
        SBOX_FF1_out[7]), .Z(SBOX_Inst_f2_abmul_pw2_0_) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_U6 ( .A(SBOX_gamma1[5]), .B(SBOX_gamma0[5]), .Z(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[5]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_U5 ( .A(SBOX_gamma0[3]), .B(SBOX_gamma1[3]), .Z(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[3]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_U4 ( .A(SBOX_gamma0[1]), .B(SBOX_gamma1[1]), .Z(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[1]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_U3 ( .A(SBOX_gamma1[4]), .B(SBOX_gamma0[4]), .Z(
        SBOX_Inst_f2_dinv_1_sA2[5]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_U2 ( .A(SBOX_gamma0[2]), .B(SBOX_gamma1[2]), .Z(
        SBOX_Inst_f2_dinv_1_sA2[3]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_U1 ( .A(SBOX_gamma0[0]), .B(SBOX_gamma1[0]), .Z(
        SBOX_Inst_f2_dinv_1_sA2[1]) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U95 ( .A1(SBOX_gamma1[2]), .A2(
        SBOX_gamma1[0]), .B1(SBOX_Inst_f2_dinv_1_mul_n302), .B2(
        SBOX_Inst_f2_dinv_1_mul_n303), .ZN(SBOX_Inst_f2_dinv_1_mul_n300) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U94 ( .A(SBOX_gamma1[0]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n302) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U93 ( .A(SBOX_Inst_f2_dinv_1_mul_n287), .B(
        SBOX_Inst_f2_dinv_1_mul_n286), .ZN(SBOX_Inst_f2_dinv_1_Orig_ab[2]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U92 ( .A(SBOX_Inst_f2_dinv_1_mul_n285), .B(
        SBOX_Inst_f2_dinv_1_mul_n284), .ZN(SBOX_Inst_f2_dinv_1_mul_n286) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U91 ( .A1(SBOX_gamma1[0]), .A2(
        SBOX_gamma0[5]), .ZN(SBOX_Inst_f2_dinv_1_mul_n284) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_mul_U90 ( .A(SBOX_Inst_f2_dinv_1_mul_n283), .B(
        SBOX_Inst_f2_dinv_1_mul_n282), .Z(SBOX_Inst_f2_dinv_1_mul_n285) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U89 ( .A(SBOX_Inst_f2_dinv_1_mul_n281), .B(
        SBOX_Inst_f2_dinv_1_mul_n280), .ZN(SBOX_Inst_f2_dinv_1_mul_n282) );
  MUX2_X1 SBOX_Inst_f2_dinv_1_mul_U88 ( .A(SBOX_gamma0[4]), .B(
        SBOX_Inst_f2_dinv_1_mul_n279), .S(SBOX_gamma1[5]), .Z(
        SBOX_Inst_f2_dinv_1_mul_n280) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U87 ( .A1(SBOX_gamma0[5]), .A2(
        SBOX_gamma0[1]), .B1(SBOX_Inst_f2_dinv_1_mul_n298), .B2(
        SBOX_Inst_f2_dinv_1_mul_n278), .ZN(SBOX_Inst_f2_dinv_1_mul_n279) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U86 ( .A(SBOX_gamma0[1]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n298) );
  OAI221_X1 SBOX_Inst_f2_dinv_1_mul_U85 ( .B1(SBOX_gamma0[5]), .B2(
        SBOX_gamma0[4]), .C1(SBOX_Inst_f2_dinv_1_mul_n278), .C2(
        SBOX_Inst_f2_dinv_1_mul_n277), .A(SBOX_gamma1[1]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n281) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U84 ( .A1(SBOX_gamma1[1]), .A2(
        SBOX_gamma0[0]), .B1(SBOX_Inst_f2_dinv_1_mul_n299), .B2(
        SBOX_Inst_f2_dinv_1_mul_n297), .ZN(SBOX_Inst_f2_dinv_1_mul_n283) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U83 ( .A(SBOX_gamma0[0]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n299) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_mul_U82 ( .A(SBOX_Inst_f2_dinv_1_mul_n276), .B(
        SBOX_Inst_f2_dinv_1_mul_n275), .Z(SBOX_Inst_f2_dinv_1_mul_n288) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U81 ( .A1(SBOX_gamma0[1]), .A2(
        SBOX_gamma1[4]), .ZN(SBOX_Inst_f2_dinv_1_mul_n275) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U80 ( .A1(SBOX_gamma0[0]), .A2(
        SBOX_gamma1[5]), .ZN(SBOX_Inst_f2_dinv_1_mul_n276) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_mul_U79 ( .A(SBOX_Inst_f2_dinv_1_mul_n274), .B(
        SBOX_Inst_f2_dinv_1_mul_n273), .Z(SBOX_Inst_f2_dinv_1_mul_n292) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U78 ( .A1(SBOX_gamma0[1]), .A2(
        SBOX_gamma1[0]), .ZN(SBOX_Inst_f2_dinv_1_mul_n273) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U77 ( .A1(SBOX_gamma1[1]), .A2(
        SBOX_gamma0[0]), .ZN(SBOX_Inst_f2_dinv_1_mul_n274) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U76 ( .A(SBOX_Inst_f2_dinv_1_mul_n272), .B(
        SBOX_Inst_f2_dinv_1_mul_n271), .ZN(SBOX_Inst_f2_dinv_1_Orig_ab[1]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U75 ( .A(SBOX_Inst_f2_dinv_1_mul_n270), .B(
        SBOX_Inst_f2_dinv_1_mul_n269), .ZN(SBOX_Inst_f2_dinv_1_mul_n271) );
  OAI221_X1 SBOX_Inst_f2_dinv_1_mul_U74 ( .B1(SBOX_gamma1[4]), .B2(
        SBOX_gamma1[3]), .C1(SBOX_Inst_f2_dinv_1_mul_n268), .C2(
        SBOX_Inst_f2_dinv_1_mul_n294), .A(SBOX_gamma0[4]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n269) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U73 ( .A(SBOX_Inst_f2_dinv_1_mul_n267), .B(
        SBOX_Inst_f2_dinv_1_mul_n266), .ZN(SBOX_Inst_f2_dinv_1_mul_n270) );
  OAI221_X1 SBOX_Inst_f2_dinv_1_mul_U72 ( .B1(SBOX_gamma0[3]), .B2(
        SBOX_gamma0[2]), .C1(SBOX_Inst_f2_dinv_1_mul_n295), .C2(
        SBOX_Inst_f2_dinv_1_mul_n301), .A(SBOX_gamma1[3]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n266) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U71 ( .A(SBOX_Inst_f2_dinv_1_mul_n265), .B(
        SBOX_gamma1[4]), .ZN(SBOX_Inst_f2_dinv_1_mul_n267) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U70 ( .A(SBOX_Inst_f2_dinv_1_mul_n264), .B(
        SBOX_Inst_f2_dinv_1_mul_n263), .ZN(SBOX_Inst_f2_dinv_1_mul_n265) );
  OAI221_X1 SBOX_Inst_f2_dinv_1_mul_U69 ( .B1(SBOX_gamma0[4]), .B2(
        SBOX_Inst_f2_dinv_1_mul_n262), .C1(SBOX_Inst_f2_dinv_1_mul_n277), .C2(
        SBOX_Inst_f2_dinv_1_mul_n261), .A(SBOX_gamma1[2]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n263) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U68 ( .A1(SBOX_gamma0[5]), .A2(
        SBOX_gamma0[2]), .B1(SBOX_Inst_f2_dinv_1_mul_n301), .B2(
        SBOX_Inst_f2_dinv_1_mul_n278), .ZN(SBOX_Inst_f2_dinv_1_mul_n262) );
  AOI221_X1 SBOX_Inst_f2_dinv_1_mul_U67 ( .B1(SBOX_gamma1[4]), .B2(
        SBOX_gamma1[2]), .C1(SBOX_Inst_f2_dinv_1_mul_n268), .C2(
        SBOX_Inst_f2_dinv_1_mul_n303), .A(SBOX_Inst_f2_dinv_1_mul_n293), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n272) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U66 ( .A1(SBOX_gamma0[3]), .A2(
        SBOX_Inst_f2_dinv_1_mul_n301), .B1(SBOX_gamma0[2]), .B2(
        SBOX_Inst_f2_dinv_1_mul_n295), .ZN(SBOX_Inst_f2_dinv_1_mul_n293) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U65 ( .A1(SBOX_gamma1[4]), .A2(
        SBOX_gamma1[5]), .B1(SBOX_Inst_f2_dinv_1_mul_n289), .B2(
        SBOX_Inst_f2_dinv_1_mul_n268), .ZN(SBOX_Inst_f2_dinv_1_mul_n290) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U64 ( .A(SBOX_gamma0[3]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n295) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U63 ( .A(SBOX_gamma0[2]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n301) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U62 ( .A(SBOX_gamma0[5]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n278) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U61 ( .A(SBOX_Inst_f2_dinv_1_mul_n260), .B(
        SBOX_Inst_f2_dinv_1_mul_n259), .ZN(SBOX_Inst_f2_dinv_1_Orig_ab[4]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U60 ( .A(SBOX_Inst_f2_dinv_1_mul_n292), .B(
        SBOX_Inst_f2_dinv_1_mul_n256), .ZN(SBOX_Inst_f2_dinv_1_mul_n260) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U59 ( .A(SBOX_Inst_f2_dinv_1_mul_n257), .B(
        SBOX_Inst_f2_dinv_1_mul_n258), .ZN(SBOX_Inst_f2_dinv_1_mul_n259) );
  NOR2_X1 SBOX_Inst_f2_dinv_1_mul_U58 ( .A1(SBOX_gamma0[3]), .A2(
        SBOX_Inst_f2_dinv_1_mul_n297), .ZN(SBOX_Inst_f2_dinv_1_mul_n258) );
  NOR2_X1 SBOX_Inst_f2_dinv_1_mul_U57 ( .A1(SBOX_Inst_f2_dinv_1_mul_n303), 
        .A2(SBOX_Inst_f2_dinv_1_mul_n293), .ZN(SBOX_Inst_f2_dinv_1_mul_n257)
         );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U56 ( .A(SBOX_Inst_f2_dinv_1_mul_n296), .B(
        SBOX_Inst_f2_dinv_1_mul_n255), .ZN(SBOX_Inst_f2_dinv_1_mul_n256) );
  MUX2_X1 SBOX_Inst_f2_dinv_1_mul_U55 ( .A(SBOX_gamma0[0]), .B(SBOX_gamma0[1]), 
        .S(SBOX_Inst_f2_dinv_1_mul_n254), .Z(SBOX_Inst_f2_dinv_1_mul_n255) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U54 ( .A1(SBOX_gamma1[3]), .A2(
        SBOX_gamma1[1]), .B1(SBOX_Inst_f2_dinv_1_mul_n297), .B2(
        SBOX_Inst_f2_dinv_1_mul_n294), .ZN(SBOX_Inst_f2_dinv_1_mul_n254) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U53 ( .A(SBOX_Inst_f2_dinv_1_mul_n252), .B(
        SBOX_Inst_f2_dinv_1_mul_n253), .ZN(SBOX_Inst_f2_dinv_1_Orig_ab[5]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_mul_U52 ( .A(SBOX_Inst_f2_dinv_1_mul_n248), .B(
        SBOX_Inst_f2_dinv_1_mul_n250), .Z(SBOX_Inst_f2_dinv_1_mul_n253) );
  AOI211_X1 SBOX_Inst_f2_dinv_1_mul_U51 ( .C1(SBOX_gamma0[0]), .C2(
        SBOX_gamma0[3]), .A(SBOX_Inst_f2_dinv_1_mul_n251), .B(
        SBOX_Inst_f2_dinv_1_mul_n294), .ZN(SBOX_Inst_f2_dinv_1_mul_n252) );
  AND2_X1 SBOX_Inst_f2_dinv_1_mul_U50 ( .A1(SBOX_Inst_f2_dinv_1_mul_n299), 
        .A2(SBOX_Inst_f2_dinv_1_mul_n295), .ZN(SBOX_Inst_f2_dinv_1_mul_n251)
         );
  AOI211_X1 SBOX_Inst_f2_dinv_1_mul_U49 ( .C1(SBOX_gamma1[0]), .C2(
        SBOX_gamma1[2]), .A(SBOX_Inst_f2_dinv_1_mul_n301), .B(
        SBOX_Inst_f2_dinv_1_mul_n249), .ZN(SBOX_Inst_f2_dinv_1_mul_n250) );
  AND2_X1 SBOX_Inst_f2_dinv_1_mul_U48 ( .A1(SBOX_Inst_f2_dinv_1_mul_n302), 
        .A2(SBOX_Inst_f2_dinv_1_mul_n303), .ZN(SBOX_Inst_f2_dinv_1_mul_n249)
         );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U47 ( .A(SBOX_Inst_f2_dinv_1_mul_n246), .B(
        SBOX_Inst_f2_dinv_1_mul_n247), .ZN(SBOX_Inst_f2_dinv_1_mul_n248) );
  NOR2_X1 SBOX_Inst_f2_dinv_1_mul_U46 ( .A1(SBOX_Inst_f2_dinv_1_mul_n298), 
        .A2(SBOX_Inst_f2_dinv_1_mul_n297), .ZN(SBOX_Inst_f2_dinv_1_mul_n247)
         );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U45 ( .A(SBOX_Inst_f2_dinv_1_mul_n296), .B(
        SBOX_Inst_f2_dinv_1_mul_n245), .ZN(SBOX_Inst_f2_dinv_1_mul_n246) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U44 ( .A1(SBOX_gamma1[1]), .A2(
        SBOX_Inst_f2_dinv_1_mul_n299), .B1(SBOX_gamma0[0]), .B2(
        SBOX_Inst_f2_dinv_1_mul_n300), .ZN(SBOX_Inst_f2_dinv_1_mul_n245) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U43 ( .A(SBOX_Inst_f2_dinv_1_mul_n244), .B(
        SBOX_Inst_f2_dinv_1_mul_n243), .ZN(SBOX_Inst_f2_dinv_1_Orig_ab[3]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U42 ( .A(SBOX_Inst_f2_dinv_1_mul_n239), .B(
        SBOX_Inst_f2_dinv_1_mul_n241), .ZN(SBOX_Inst_f2_dinv_1_mul_n244) );
  OAI221_X1 SBOX_Inst_f2_dinv_1_mul_U41 ( .B1(SBOX_Inst_f2_dinv_1_mul_n233), 
        .B2(SBOX_gamma1[1]), .C1(SBOX_Inst_f2_dinv_1_mul_n242), .C2(
        SBOX_Inst_f2_dinv_1_mul_n297), .A(SBOX_gamma0[4]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n243) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U40 ( .A(SBOX_Inst_f2_dinv_1_mul_n233), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n242) );
  OAI21_X1 SBOX_Inst_f2_dinv_1_mul_U39 ( .B1(SBOX_Inst_f2_dinv_1_mul_n291), 
        .B2(SBOX_Inst_f2_dinv_1_mul_n290), .A(SBOX_Inst_f2_dinv_1_mul_n240), 
        .ZN(SBOX_Inst_f2_dinv_1_mul_n241) );
  NAND3_X1 SBOX_Inst_f2_dinv_1_mul_U38 ( .A1(SBOX_Inst_f2_dinv_1_mul_n291), 
        .A2(SBOX_gamma1[4]), .A3(SBOX_Inst_f2_dinv_1_mul_n289), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n240) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U37 ( .A(SBOX_Inst_f2_dinv_1_mul_n237), .B(
        SBOX_Inst_f2_dinv_1_mul_n238), .ZN(SBOX_Inst_f2_dinv_1_mul_n239) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U36 ( .A1(SBOX_Inst_f2_dinv_1_mul_n233), 
        .A2(SBOX_gamma0[5]), .ZN(SBOX_Inst_f2_dinv_1_mul_n238) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_mul_U35 ( .A(SBOX_Inst_f2_dinv_1_mul_n288), .B(
        SBOX_Inst_f2_dinv_1_mul_n236), .Z(SBOX_Inst_f2_dinv_1_mul_n237) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_mul_U34 ( .A(SBOX_Inst_f2_dinv_1_mul_n234), .B(
        SBOX_Inst_f2_dinv_1_mul_n235), .Z(SBOX_Inst_f2_dinv_1_mul_n236) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U33 ( .A1(SBOX_gamma0[0]), .A2(
        SBOX_gamma1[4]), .ZN(SBOX_Inst_f2_dinv_1_mul_n235) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U32 ( .A1(SBOX_Inst_f2_dinv_1_mul_n298), 
        .A2(SBOX_gamma1[1]), .ZN(SBOX_Inst_f2_dinv_1_mul_n234) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U31 ( .A1(SBOX_gamma1[5]), .A2(
        SBOX_gamma1[0]), .B1(SBOX_Inst_f2_dinv_1_mul_n289), .B2(
        SBOX_Inst_f2_dinv_1_mul_n302), .ZN(SBOX_Inst_f2_dinv_1_mul_n233) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U30 ( .A(SBOX_Inst_f2_dinv_1_mul_n230), .B(
        SBOX_Inst_f2_dinv_1_mul_n232), .ZN(SBOX_Inst_f2_dinv_1_Orig_ab[0]) );
  OAI22_X1 SBOX_Inst_f2_dinv_1_mul_U29 ( .A1(SBOX_Inst_f2_dinv_1_mul_n278), 
        .A2(SBOX_Inst_f2_dinv_1_mul_n231), .B1(SBOX_Inst_f2_dinv_1_mul_n291), 
        .B2(SBOX_gamma0[4]), .ZN(SBOX_Inst_f2_dinv_1_mul_n232) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U28 ( .A1(SBOX_gamma0[4]), .A2(
        SBOX_gamma1[4]), .ZN(SBOX_Inst_f2_dinv_1_mul_n231) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U27 ( .A(SBOX_Inst_f2_dinv_1_mul_n229), .B(
        SBOX_Inst_f2_dinv_1_mul_n228), .ZN(SBOX_Inst_f2_dinv_1_mul_n230) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U26 ( .A1(SBOX_Inst_f2_dinv_1_mul_n290), 
        .A2(SBOX_gamma0[3]), .ZN(SBOX_Inst_f2_dinv_1_mul_n229) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U25 ( .A(SBOX_Inst_f2_dinv_1_mul_n227), .B(
        SBOX_Inst_f2_dinv_1_mul_n221), .ZN(SBOX_Inst_f2_dinv_1_mul_n228) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U24 ( .A(SBOX_Inst_f2_dinv_1_mul_n226), .B(
        SBOX_Inst_f2_dinv_1_mul_n223), .ZN(SBOX_Inst_f2_dinv_1_mul_n227) );
  NOR2_X1 SBOX_Inst_f2_dinv_1_mul_U23 ( .A1(SBOX_Inst_f2_dinv_1_mul_n225), 
        .A2(SBOX_Inst_f2_dinv_1_mul_n224), .ZN(SBOX_Inst_f2_dinv_1_mul_n226)
         );
  OAI22_X1 SBOX_Inst_f2_dinv_1_mul_U22 ( .A1(SBOX_gamma1[5]), .A2(
        SBOX_gamma1[3]), .B1(SBOX_Inst_f2_dinv_1_mul_n289), .B2(
        SBOX_Inst_f2_dinv_1_mul_n294), .ZN(SBOX_Inst_f2_dinv_1_mul_n225) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U21 ( .A(SBOX_gamma0[2]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n224) );
  OAI211_X1 SBOX_Inst_f2_dinv_1_mul_U20 ( .C1(SBOX_gamma0[2]), .C2(
        SBOX_gamma0[5]), .A(SBOX_gamma1[2]), .B(SBOX_Inst_f2_dinv_1_mul_n222), 
        .ZN(SBOX_Inst_f2_dinv_1_mul_n223) );
  OR2_X1 SBOX_Inst_f2_dinv_1_mul_U19 ( .A1(SBOX_Inst_f2_dinv_1_mul_n278), .A2(
        SBOX_Inst_f2_dinv_1_mul_n301), .ZN(SBOX_Inst_f2_dinv_1_mul_n222) );
  OAI211_X1 SBOX_Inst_f2_dinv_1_mul_U18 ( .C1(SBOX_Inst_f2_dinv_1_mul_n219), 
        .C2(SBOX_gamma0[4]), .A(SBOX_gamma1[3]), .B(
        SBOX_Inst_f2_dinv_1_mul_n220), .ZN(SBOX_Inst_f2_dinv_1_mul_n221) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U17 ( .A1(SBOX_Inst_f2_dinv_1_mul_n219), 
        .A2(SBOX_gamma0[4]), .ZN(SBOX_Inst_f2_dinv_1_mul_n220) );
  AOI22_X1 SBOX_Inst_f2_dinv_1_mul_U16 ( .A1(SBOX_gamma0[3]), .A2(
        SBOX_gamma0[5]), .B1(SBOX_Inst_f2_dinv_1_mul_n278), .B2(
        SBOX_Inst_f2_dinv_1_mul_n295), .ZN(SBOX_Inst_f2_dinv_1_mul_n219) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U15 ( .A(SBOX_Inst_f2_dinv_1_mul_n215), .B(
        SBOX_Inst_f2_dinv_1_mul_n218), .ZN(SBOX_Inst_f2_dinv_1_mul_n296) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_mul_U14 ( .A(SBOX_Inst_f2_dinv_1_mul_n216), .B(
        SBOX_Inst_f2_dinv_1_mul_n217), .Z(SBOX_Inst_f2_dinv_1_mul_n218) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U13 ( .A1(SBOX_gamma0[3]), .A2(
        SBOX_gamma1[0]), .ZN(SBOX_Inst_f2_dinv_1_mul_n217) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U12 ( .A1(SBOX_gamma1[1]), .A2(
        SBOX_gamma0[2]), .ZN(SBOX_Inst_f2_dinv_1_mul_n216) );
  NAND2_X1 SBOX_Inst_f2_dinv_1_mul_U11 ( .A1(SBOX_Inst_f2_dinv_1_mul_n300), 
        .A2(SBOX_gamma0[1]), .ZN(SBOX_Inst_f2_dinv_1_mul_n215) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_mul_U10 ( .A(SBOX_Inst_f2_dinv_1_mul_n292), .B(
        SBOX_Inst_f2_dinv_1_mul_n288), .ZN(SBOX_Inst_f2_dinv_1_mul_n287) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U9 ( .A(SBOX_Inst_f2_dinv_1_mul_n262), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n261) );
  NOR2_X1 SBOX_Inst_f2_dinv_1_mul_U8 ( .A1(SBOX_Inst_f2_dinv_1_mul_n262), .A2(
        SBOX_Inst_f2_dinv_1_mul_n289), .ZN(SBOX_Inst_f2_dinv_1_mul_n264) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U7 ( .A(SBOX_gamma1[1]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n297) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U6 ( .A(SBOX_gamma1[2]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n303) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U5 ( .A(SBOX_gamma1[3]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n294) );
  NOR2_X1 SBOX_Inst_f2_dinv_1_mul_U4 ( .A1(SBOX_Inst_f2_dinv_1_mul_n268), .A2(
        SBOX_Inst_f2_dinv_1_mul_n278), .ZN(SBOX_Inst_f2_dinv_1_mul_n291) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U3 ( .A(SBOX_gamma1[5]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n289) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U2 ( .A(SBOX_gamma0[4]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n277) );
  INV_X1 SBOX_Inst_f2_dinv_1_mul_U1 ( .A(SBOX_gamma1[4]), .ZN(
        SBOX_Inst_f2_dinv_1_mul_n268) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U8 ( .A(PRNGQ[14]), .B(
        SBOX_Inst_f2_dinv_1_Orig_ab[2]), .Z(SBOX_ab[2]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U7 ( .A(PRNGQ[13]), .B(
        SBOX_Inst_f2_dinv_1_Orig_ab[1]), .Z(SBOX_ab[1]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U6 ( .A(
        SBOX_Inst_f2_dinv_1_AddNewMaskab_n6), .B(PRNGQ[14]), .ZN(SBOX_ab[4])
         );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U5 ( .A(PRNGQ[12]), .B(
        SBOX_Inst_f2_dinv_1_Orig_ab[4]), .ZN(
        SBOX_Inst_f2_dinv_1_AddNewMaskab_n6) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U4 ( .A(
        SBOX_Inst_f2_dinv_1_AddNewMaskab_n5), .B(PRNGQ[15]), .ZN(SBOX_ab[5])
         );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U3 ( .A(PRNGQ[13]), .B(
        SBOX_Inst_f2_dinv_1_Orig_ab[5]), .ZN(
        SBOX_Inst_f2_dinv_1_AddNewMaskab_n5) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U2 ( .A(PRNGQ[15]), .B(
        SBOX_Inst_f2_dinv_1_Orig_ab[3]), .Z(SBOX_ab[3]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMaskab_U1 ( .A(PRNGQ[12]), .B(
        SBOX_Inst_f2_dinv_1_Orig_ab[0]), .Z(SBOX_ab[0]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_NxGAMMA_U3 ( .A(SBOX_Inst_f2_dinv_1_Orig_sA2N[5]), .B(SBOX_Inst_f2_dinv_1_sA2[5]), .Z(SBOX_Inst_f2_dinv_1_Orig_sA2N[4]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_NxGAMMA_U2 ( .A(SBOX_Inst_f2_dinv_1_Orig_sA2N[3]), .B(SBOX_Inst_f2_dinv_1_sA2[3]), .Z(SBOX_Inst_f2_dinv_1_Orig_sA2N[2]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_NxGAMMA_U1 ( .A(SBOX_Inst_f2_dinv_1_Orig_sA2N[1]), .B(SBOX_Inst_f2_dinv_1_sA2[1]), .Z(SBOX_Inst_f2_dinv_1_Orig_sA2N[0]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U8 ( .A(
        SBOX_Inst_f2_dinv_1_AddNewMasksA2N_n6), .B(PRNGQ[19]), .ZN(
        SBOX_sA2N[5]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U7 ( .A(PRNGQ[17]), .B(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[5]), .ZN(
        SBOX_Inst_f2_dinv_1_AddNewMasksA2N_n6) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U6 ( .A(PRNGQ[19]), .B(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[3]), .Z(SBOX_sA2N[3]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U5 ( .A(PRNGQ[17]), .B(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[1]), .Z(SBOX_sA2N[1]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U4 ( .A(
        SBOX_Inst_f2_dinv_1_AddNewMasksA2N_n5), .B(PRNGQ[18]), .ZN(
        SBOX_sA2N[4]) );
  XNOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U3 ( .A(PRNGQ[16]), .B(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[4]), .ZN(
        SBOX_Inst_f2_dinv_1_AddNewMasksA2N_n5) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U2 ( .A(PRNGQ[18]), .B(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[2]), .Z(SBOX_sA2N[2]) );
  XOR2_X1 SBOX_Inst_f2_dinv_1_AddNewMasksA2N_U1 ( .A(PRNGQ[16]), .B(
        SBOX_Inst_f2_dinv_1_Orig_sA2N[0]), .Z(SBOX_sA2N[0]) );
  OAI21_X1 SBOX_PL_2_U97 ( .B1(1'b1), .B2(SBOX_PL_2_n51), .A(SBOX_PL_2_n48), 
        .ZN(SBOX_PL_2_n99) );
  NAND2_X1 SBOX_PL_2_U96 ( .A1(1'b1), .A2(SBOX_gamma0[2]), .ZN(SBOX_PL_2_n48)
         );
  OAI21_X1 SBOX_PL_2_U95 ( .B1(1'b1), .B2(SBOX_PL_2_n49), .A(SBOX_PL_2_n47), 
        .ZN(SBOX_PL_2_n97) );
  NAND2_X1 SBOX_PL_2_U94 ( .A1(1'b1), .A2(SBOX_gamma0[0]), .ZN(SBOX_PL_2_n47)
         );
  OAI21_X1 SBOX_PL_2_U93 ( .B1(1'b1), .B2(SBOX_PL_2_n96), .A(SBOX_PL_2_n46), 
        .ZN(SBOX_PL_2_n144) );
  NAND2_X1 SBOX_PL_2_U92 ( .A1(1'b1), .A2(SBOX_Zh_f2[11]), .ZN(SBOX_PL_2_n46)
         );
  OAI21_X1 SBOX_PL_2_U91 ( .B1(1'b1), .B2(SBOX_PL_2_n95), .A(SBOX_PL_2_n45), 
        .ZN(SBOX_PL_2_n143) );
  NAND2_X1 SBOX_PL_2_U90 ( .A1(1'b1), .A2(SBOX_Zh_f2[10]), .ZN(SBOX_PL_2_n45)
         );
  OAI21_X1 SBOX_PL_2_U89 ( .B1(1'b1), .B2(SBOX_PL_2_n94), .A(SBOX_PL_2_n44), 
        .ZN(SBOX_PL_2_n142) );
  NAND2_X1 SBOX_PL_2_U88 ( .A1(1'b1), .A2(SBOX_Zh_f2[9]), .ZN(SBOX_PL_2_n44)
         );
  OAI21_X1 SBOX_PL_2_U87 ( .B1(1'b1), .B2(SBOX_PL_2_n93), .A(SBOX_PL_2_n43), 
        .ZN(SBOX_PL_2_n141) );
  NAND2_X1 SBOX_PL_2_U86 ( .A1(1'b1), .A2(SBOX_Zh_f2[8]), .ZN(SBOX_PL_2_n43)
         );
  OAI21_X1 SBOX_PL_2_U85 ( .B1(1'b1), .B2(SBOX_PL_2_n92), .A(SBOX_PL_2_n42), 
        .ZN(SBOX_PL_2_n140) );
  NAND2_X1 SBOX_PL_2_U84 ( .A1(1'b1), .A2(SBOX_Zh_f2[7]), .ZN(SBOX_PL_2_n42)
         );
  OAI21_X1 SBOX_PL_2_U83 ( .B1(1'b1), .B2(SBOX_PL_2_n91), .A(SBOX_PL_2_n41), 
        .ZN(SBOX_PL_2_n139) );
  NAND2_X1 SBOX_PL_2_U82 ( .A1(1'b1), .A2(SBOX_Zh_f2[6]), .ZN(SBOX_PL_2_n41)
         );
  OAI21_X1 SBOX_PL_2_U81 ( .B1(1'b1), .B2(SBOX_PL_2_n90), .A(SBOX_PL_2_n40), 
        .ZN(SBOX_PL_2_n138) );
  NAND2_X1 SBOX_PL_2_U80 ( .A1(1'b1), .A2(SBOX_Zh_f2[5]), .ZN(SBOX_PL_2_n40)
         );
  OAI21_X1 SBOX_PL_2_U79 ( .B1(1'b1), .B2(SBOX_PL_2_n89), .A(SBOX_PL_2_n39), 
        .ZN(SBOX_PL_2_n137) );
  NAND2_X1 SBOX_PL_2_U78 ( .A1(1'b1), .A2(SBOX_Zh_f2[4]), .ZN(SBOX_PL_2_n39)
         );
  OAI21_X1 SBOX_PL_2_U77 ( .B1(1'b1), .B2(SBOX_PL_2_n88), .A(SBOX_PL_2_n38), 
        .ZN(SBOX_PL_2_n136) );
  NAND2_X1 SBOX_PL_2_U76 ( .A1(1'b1), .A2(SBOX_Zh_f2[3]), .ZN(SBOX_PL_2_n38)
         );
  OAI21_X1 SBOX_PL_2_U75 ( .B1(1'b1), .B2(SBOX_PL_2_n87), .A(SBOX_PL_2_n37), 
        .ZN(SBOX_PL_2_n135) );
  NAND2_X1 SBOX_PL_2_U74 ( .A1(1'b1), .A2(SBOX_Zh_f2[2]), .ZN(SBOX_PL_2_n37)
         );
  OAI21_X1 SBOX_PL_2_U73 ( .B1(1'b1), .B2(SBOX_PL_2_n86), .A(SBOX_PL_2_n36), 
        .ZN(SBOX_PL_2_n134) );
  NAND2_X1 SBOX_PL_2_U72 ( .A1(1'b1), .A2(SBOX_Zh_f2[1]), .ZN(SBOX_PL_2_n36)
         );
  OAI21_X1 SBOX_PL_2_U71 ( .B1(1'b1), .B2(SBOX_PL_2_n85), .A(SBOX_PL_2_n35), 
        .ZN(SBOX_PL_2_n133) );
  NAND2_X1 SBOX_PL_2_U70 ( .A1(1'b1), .A2(SBOX_Zh_f2[0]), .ZN(SBOX_PL_2_n35)
         );
  OAI21_X1 SBOX_PL_2_U69 ( .B1(1'b1), .B2(SBOX_PL_2_n84), .A(SBOX_PL_2_n34), 
        .ZN(SBOX_PL_2_n132) );
  NAND2_X1 SBOX_PL_2_U68 ( .A1(1'b1), .A2(SBOX_Zl_f2[11]), .ZN(SBOX_PL_2_n34)
         );
  OAI21_X1 SBOX_PL_2_U67 ( .B1(1'b1), .B2(SBOX_PL_2_n83), .A(SBOX_PL_2_n33), 
        .ZN(SBOX_PL_2_n131) );
  NAND2_X1 SBOX_PL_2_U66 ( .A1(1'b1), .A2(SBOX_Zl_f2[10]), .ZN(SBOX_PL_2_n33)
         );
  OAI21_X1 SBOX_PL_2_U65 ( .B1(1'b1), .B2(SBOX_PL_2_n82), .A(SBOX_PL_2_n32), 
        .ZN(SBOX_PL_2_n130) );
  NAND2_X1 SBOX_PL_2_U64 ( .A1(1'b1), .A2(SBOX_Zl_f2[9]), .ZN(SBOX_PL_2_n32)
         );
  OAI21_X1 SBOX_PL_2_U63 ( .B1(1'b1), .B2(SBOX_PL_2_n81), .A(SBOX_PL_2_n31), 
        .ZN(SBOX_PL_2_n129) );
  NAND2_X1 SBOX_PL_2_U62 ( .A1(1'b1), .A2(SBOX_Zl_f2[8]), .ZN(SBOX_PL_2_n31)
         );
  OAI21_X1 SBOX_PL_2_U61 ( .B1(1'b1), .B2(SBOX_PL_2_n80), .A(SBOX_PL_2_n30), 
        .ZN(SBOX_PL_2_n128) );
  NAND2_X1 SBOX_PL_2_U60 ( .A1(1'b1), .A2(SBOX_Zl_f2[7]), .ZN(SBOX_PL_2_n30)
         );
  OAI21_X1 SBOX_PL_2_U59 ( .B1(1'b1), .B2(SBOX_PL_2_n79), .A(SBOX_PL_2_n29), 
        .ZN(SBOX_PL_2_n127) );
  NAND2_X1 SBOX_PL_2_U58 ( .A1(1'b1), .A2(SBOX_Zl_f2[6]), .ZN(SBOX_PL_2_n29)
         );
  OAI21_X1 SBOX_PL_2_U57 ( .B1(1'b1), .B2(SBOX_PL_2_n78), .A(SBOX_PL_2_n28), 
        .ZN(SBOX_PL_2_n126) );
  NAND2_X1 SBOX_PL_2_U56 ( .A1(1'b1), .A2(SBOX_Zl_f2[5]), .ZN(SBOX_PL_2_n28)
         );
  OAI21_X1 SBOX_PL_2_U55 ( .B1(1'b1), .B2(SBOX_PL_2_n77), .A(SBOX_PL_2_n27), 
        .ZN(SBOX_PL_2_n125) );
  NAND2_X1 SBOX_PL_2_U54 ( .A1(1'b1), .A2(SBOX_Zl_f2[4]), .ZN(SBOX_PL_2_n27)
         );
  OAI21_X1 SBOX_PL_2_U53 ( .B1(1'b1), .B2(SBOX_PL_2_n76), .A(SBOX_PL_2_n26), 
        .ZN(SBOX_PL_2_n124) );
  NAND2_X1 SBOX_PL_2_U52 ( .A1(1'b1), .A2(SBOX_Zl_f2[3]), .ZN(SBOX_PL_2_n26)
         );
  OAI21_X1 SBOX_PL_2_U51 ( .B1(1'b1), .B2(SBOX_PL_2_n75), .A(SBOX_PL_2_n25), 
        .ZN(SBOX_PL_2_n123) );
  NAND2_X1 SBOX_PL_2_U50 ( .A1(1'b1), .A2(SBOX_Zl_f2[2]), .ZN(SBOX_PL_2_n25)
         );
  OAI21_X1 SBOX_PL_2_U49 ( .B1(1'b1), .B2(SBOX_PL_2_n74), .A(SBOX_PL_2_n24), 
        .ZN(SBOX_PL_2_n122) );
  NAND2_X1 SBOX_PL_2_U48 ( .A1(1'b1), .A2(SBOX_Zl_f2[1]), .ZN(SBOX_PL_2_n24)
         );
  OAI21_X1 SBOX_PL_2_U47 ( .B1(1'b1), .B2(SBOX_PL_2_n73), .A(SBOX_PL_2_n23), 
        .ZN(SBOX_PL_2_n121) );
  NAND2_X1 SBOX_PL_2_U46 ( .A1(1'b1), .A2(SBOX_Zl_f2[0]), .ZN(SBOX_PL_2_n23)
         );
  OAI21_X1 SBOX_PL_2_U45 ( .B1(1'b1), .B2(SBOX_PL_2_n71), .A(SBOX_PL_2_n22), 
        .ZN(SBOX_PL_2_n119) );
  NAND2_X1 SBOX_PL_2_U44 ( .A1(1'b1), .A2(SBOX_gamma1[4]), .ZN(SBOX_PL_2_n22)
         );
  OAI21_X1 SBOX_PL_2_U43 ( .B1(1'b1), .B2(SBOX_PL_2_n57), .A(SBOX_PL_2_n21), 
        .ZN(SBOX_PL_2_n105) );
  NAND2_X1 SBOX_PL_2_U42 ( .A1(1'b1), .A2(SBOX_ab[2]), .ZN(SBOX_PL_2_n21) );
  OAI21_X1 SBOX_PL_2_U41 ( .B1(1'b1), .B2(SBOX_PL_2_n56), .A(SBOX_PL_2_n20), 
        .ZN(SBOX_PL_2_n104) );
  NAND2_X1 SBOX_PL_2_U40 ( .A1(1'b1), .A2(SBOX_ab[1]), .ZN(SBOX_PL_2_n20) );
  OAI21_X1 SBOX_PL_2_U39 ( .B1(1'b1), .B2(SBOX_PL_2_n54), .A(SBOX_PL_2_n19), 
        .ZN(SBOX_PL_2_n102) );
  NAND2_X1 SBOX_PL_2_U38 ( .A1(1'b1), .A2(SBOX_gamma0[5]), .ZN(SBOX_PL_2_n19)
         );
  OAI21_X1 SBOX_PL_2_U37 ( .B1(1'b1), .B2(SBOX_PL_2_n52), .A(SBOX_PL_2_n18), 
        .ZN(SBOX_PL_2_n100) );
  NAND2_X1 SBOX_PL_2_U36 ( .A1(1'b1), .A2(SBOX_gamma0[3]), .ZN(SBOX_PL_2_n18)
         );
  OAI21_X1 SBOX_PL_2_U35 ( .B1(1'b1), .B2(SBOX_PL_2_n72), .A(SBOX_PL_2_n17), 
        .ZN(SBOX_PL_2_n120) );
  NAND2_X1 SBOX_PL_2_U34 ( .A1(1'b1), .A2(SBOX_gamma1[5]), .ZN(SBOX_PL_2_n17)
         );
  OAI21_X1 SBOX_PL_2_U33 ( .B1(1'b1), .B2(SBOX_PL_2_n70), .A(SBOX_PL_2_n16), 
        .ZN(SBOX_PL_2_n118) );
  NAND2_X1 SBOX_PL_2_U32 ( .A1(1'b1), .A2(SBOX_gamma1[3]), .ZN(SBOX_PL_2_n16)
         );
  OAI21_X1 SBOX_PL_2_U31 ( .B1(1'b1), .B2(SBOX_PL_2_n69), .A(SBOX_PL_2_n15), 
        .ZN(SBOX_PL_2_n117) );
  NAND2_X1 SBOX_PL_2_U30 ( .A1(1'b1), .A2(SBOX_gamma1[2]), .ZN(SBOX_PL_2_n15)
         );
  OAI21_X1 SBOX_PL_2_U29 ( .B1(1'b1), .B2(SBOX_PL_2_n68), .A(SBOX_PL_2_n14), 
        .ZN(SBOX_PL_2_n116) );
  NAND2_X1 SBOX_PL_2_U28 ( .A1(1'b1), .A2(SBOX_gamma1[1]), .ZN(SBOX_PL_2_n14)
         );
  OAI21_X1 SBOX_PL_2_U27 ( .B1(1'b1), .B2(SBOX_PL_2_n67), .A(SBOX_PL_2_n13), 
        .ZN(SBOX_PL_2_n115) );
  NAND2_X1 SBOX_PL_2_U26 ( .A1(1'b1), .A2(SBOX_gamma1[0]), .ZN(SBOX_PL_2_n13)
         );
  OAI21_X1 SBOX_PL_2_U25 ( .B1(1'b1), .B2(SBOX_PL_2_n50), .A(SBOX_PL_2_n12), 
        .ZN(SBOX_PL_2_n98) );
  NAND2_X1 SBOX_PL_2_U24 ( .A1(1'b1), .A2(SBOX_gamma0[1]), .ZN(SBOX_PL_2_n12)
         );
  OAI21_X1 SBOX_PL_2_U23 ( .B1(1'b1), .B2(SBOX_PL_2_n66), .A(SBOX_PL_2_n11), 
        .ZN(SBOX_PL_2_n114) );
  NAND2_X1 SBOX_PL_2_U22 ( .A1(1'b1), .A2(SBOX_sA2N[5]), .ZN(SBOX_PL_2_n11) );
  OAI21_X1 SBOX_PL_2_U21 ( .B1(1'b1), .B2(SBOX_PL_2_n64), .A(SBOX_PL_2_n10), 
        .ZN(SBOX_PL_2_n112) );
  NAND2_X1 SBOX_PL_2_U20 ( .A1(1'b1), .A2(SBOX_sA2N[3]), .ZN(SBOX_PL_2_n10) );
  OAI21_X1 SBOX_PL_2_U19 ( .B1(1'b1), .B2(SBOX_PL_2_n62), .A(SBOX_PL_2_n9), 
        .ZN(SBOX_PL_2_n110) );
  NAND2_X1 SBOX_PL_2_U18 ( .A1(1'b1), .A2(SBOX_sA2N[1]), .ZN(SBOX_PL_2_n9) );
  OAI21_X1 SBOX_PL_2_U17 ( .B1(1'b1), .B2(SBOX_PL_2_n53), .A(SBOX_PL_2_n8), 
        .ZN(SBOX_PL_2_n101) );
  NAND2_X1 SBOX_PL_2_U16 ( .A1(1'b1), .A2(SBOX_gamma0[4]), .ZN(SBOX_PL_2_n8)
         );
  OAI21_X1 SBOX_PL_2_U15 ( .B1(1'b1), .B2(SBOX_PL_2_n65), .A(SBOX_PL_2_n7), 
        .ZN(SBOX_PL_2_n113) );
  NAND2_X1 SBOX_PL_2_U14 ( .A1(1'b1), .A2(SBOX_sA2N[4]), .ZN(SBOX_PL_2_n7) );
  OAI21_X1 SBOX_PL_2_U13 ( .B1(1'b1), .B2(SBOX_PL_2_n63), .A(SBOX_PL_2_n6), 
        .ZN(SBOX_PL_2_n111) );
  NAND2_X1 SBOX_PL_2_U12 ( .A1(1'b1), .A2(SBOX_sA2N[2]), .ZN(SBOX_PL_2_n6) );
  OAI21_X1 SBOX_PL_2_U11 ( .B1(1'b1), .B2(SBOX_PL_2_n61), .A(SBOX_PL_2_n5), 
        .ZN(SBOX_PL_2_n109) );
  NAND2_X1 SBOX_PL_2_U10 ( .A1(1'b1), .A2(SBOX_sA2N[0]), .ZN(SBOX_PL_2_n5) );
  OAI21_X1 SBOX_PL_2_U9 ( .B1(1'b1), .B2(SBOX_PL_2_n59), .A(SBOX_PL_2_n4), 
        .ZN(SBOX_PL_2_n107) );
  NAND2_X1 SBOX_PL_2_U8 ( .A1(1'b1), .A2(SBOX_ab[4]), .ZN(SBOX_PL_2_n4) );
  OAI21_X1 SBOX_PL_2_U7 ( .B1(1'b1), .B2(SBOX_PL_2_n60), .A(SBOX_PL_2_n3), 
        .ZN(SBOX_PL_2_n108) );
  NAND2_X1 SBOX_PL_2_U6 ( .A1(1'b1), .A2(SBOX_ab[5]), .ZN(SBOX_PL_2_n3) );
  OAI21_X1 SBOX_PL_2_U5 ( .B1(1'b1), .B2(SBOX_PL_2_n58), .A(SBOX_PL_2_n2), 
        .ZN(SBOX_PL_2_n106) );
  NAND2_X1 SBOX_PL_2_U4 ( .A1(1'b1), .A2(SBOX_ab[3]), .ZN(SBOX_PL_2_n2) );
  OAI21_X1 SBOX_PL_2_U3 ( .B1(1'b1), .B2(SBOX_PL_2_n55), .A(SBOX_PL_2_n1), 
        .ZN(SBOX_PL_2_n103) );
  NAND2_X1 SBOX_PL_2_U2 ( .A1(1'b1), .A2(SBOX_ab[0]), .ZN(SBOX_PL_2_n1) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_0_ ( .D(SBOX_PL_2_n97), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[0]), .QN(SBOX_PL_2_n49) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_1_ ( .D(SBOX_PL_2_n98), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[1]), .QN(SBOX_PL_2_n50) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_2_ ( .D(SBOX_PL_2_n99), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[2]), .QN(SBOX_PL_2_n51) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_3_ ( .D(SBOX_PL_2_n100), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[3]), .QN(SBOX_PL_2_n52) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_4_ ( .D(SBOX_PL_2_n101), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[4]), .QN(SBOX_PL_2_n53) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_5_ ( .D(SBOX_PL_2_n102), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[5]), .QN(SBOX_PL_2_n54) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_6_ ( .D(SBOX_PL_2_n103), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[6]), .QN(SBOX_PL_2_n55) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_7_ ( .D(SBOX_PL_2_n104), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[7]), .QN(SBOX_PL_2_n56) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_8_ ( .D(SBOX_PL_2_n105), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[8]), .QN(SBOX_PL_2_n57) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_9_ ( .D(SBOX_PL_2_n106), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[9]), .QN(SBOX_PL_2_n58) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_10_ ( .D(SBOX_PL_2_n107), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[10]), .QN(SBOX_PL_2_n59) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_11_ ( .D(SBOX_PL_2_n108), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[11]), .QN(SBOX_PL_2_n60) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_12_ ( .D(SBOX_PL_2_n109), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[12]), .QN(SBOX_PL_2_n61) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_13_ ( .D(SBOX_PL_2_n110), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[13]), .QN(SBOX_PL_2_n62) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_14_ ( .D(SBOX_PL_2_n111), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[14]), .QN(SBOX_PL_2_n63) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_15_ ( .D(SBOX_PL_2_n112), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[15]), .QN(SBOX_PL_2_n64) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_16_ ( .D(SBOX_PL_2_n113), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[16]), .QN(SBOX_PL_2_n65) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_17_ ( .D(SBOX_PL_2_n114), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[17]), .QN(SBOX_PL_2_n66) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_18_ ( .D(SBOX_PL_2_n115), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[18]), .QN(SBOX_PL_2_n67) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_19_ ( .D(SBOX_PL_2_n116), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[19]), .QN(SBOX_PL_2_n68) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_20_ ( .D(SBOX_PL_2_n117), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[20]), .QN(SBOX_PL_2_n69) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_21_ ( .D(SBOX_PL_2_n118), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[21]), .QN(SBOX_PL_2_n70) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_22_ ( .D(SBOX_PL_2_n119), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[22]), .QN(SBOX_PL_2_n71) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_23_ ( .D(SBOX_PL_2_n120), .CK(ClkxCI), 
        .Q(SBOX_FF2_out[23]), .QN(SBOX_PL_2_n72) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_24_ ( .D(SBOX_PL_2_n121), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[0]), .QN(SBOX_PL_2_n73) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_25_ ( .D(SBOX_PL_2_n122), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[1]), .QN(SBOX_PL_2_n74) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_26_ ( .D(SBOX_PL_2_n123), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[2]), .QN(SBOX_PL_2_n75) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_27_ ( .D(SBOX_PL_2_n124), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[3]), .QN(SBOX_PL_2_n76) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_28_ ( .D(SBOX_PL_2_n125), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[4]), .QN(SBOX_PL_2_n77) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_29_ ( .D(SBOX_PL_2_n126), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[5]), .QN(SBOX_PL_2_n78) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_30_ ( .D(SBOX_PL_2_n127), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[6]), .QN(SBOX_PL_2_n79) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_31_ ( .D(SBOX_PL_2_n128), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[7]), .QN(SBOX_PL_2_n80) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_32_ ( .D(SBOX_PL_2_n129), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[8]), .QN(SBOX_PL_2_n81) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_33_ ( .D(SBOX_PL_2_n130), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[9]), .QN(SBOX_PL_2_n82) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_34_ ( .D(SBOX_PL_2_n131), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[10]), .QN(SBOX_PL_2_n83) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_35_ ( .D(SBOX_PL_2_n132), .CK(ClkxCI), 
        .Q(SBOX_Zl_f3[11]), .QN(SBOX_PL_2_n84) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_36_ ( .D(SBOX_PL_2_n133), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[0]), .QN(SBOX_PL_2_n85) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_37_ ( .D(SBOX_PL_2_n134), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[1]), .QN(SBOX_PL_2_n86) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_38_ ( .D(SBOX_PL_2_n135), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[2]), .QN(SBOX_PL_2_n87) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_39_ ( .D(SBOX_PL_2_n136), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[3]), .QN(SBOX_PL_2_n88) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_40_ ( .D(SBOX_PL_2_n137), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[4]), .QN(SBOX_PL_2_n89) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_41_ ( .D(SBOX_PL_2_n138), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[5]), .QN(SBOX_PL_2_n90) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_42_ ( .D(SBOX_PL_2_n139), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[6]), .QN(SBOX_PL_2_n91) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_43_ ( .D(SBOX_PL_2_n140), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[7]), .QN(SBOX_PL_2_n92) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_44_ ( .D(SBOX_PL_2_n141), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[8]), .QN(SBOX_PL_2_n93) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_45_ ( .D(SBOX_PL_2_n142), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[9]), .QN(SBOX_PL_2_n94) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_46_ ( .D(SBOX_PL_2_n143), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[10]), .QN(SBOX_PL_2_n95) );
  DFF_X1 SBOX_PL_2_s_current_state_reg_47_ ( .D(SBOX_PL_2_n144), .CK(ClkxCI), 
        .Q(SBOX_Zh_f3[11]), .QN(SBOX_PL_2_n96) );
  XOR2_X2 SBOX_Inst_f3_dinv_2_U6 ( .A(SBOX_FF2_out[11]), .B(SBOX_FF2_out[17]), 
        .Z(SBOX_Inst_f3_dinv_2_d_4_) );
  XOR2_X2 SBOX_Inst_f3_dinv_2_U5 ( .A(SBOX_FF2_out[7]), .B(SBOX_FF2_out[13]), 
        .Z(SBOX_Inst_f3_dinv_2_d_0_) );
  XOR2_X2 SBOX_Inst_f3_dinv_2_U4 ( .A(SBOX_FF2_out[6]), .B(SBOX_FF2_out[12]), 
        .Z(SBOX_Inst_f3_dinv_2_d_1_) );
  XOR2_X2 SBOX_Inst_f3_dinv_2_U3 ( .A(SBOX_FF2_out[10]), .B(SBOX_FF2_out[16]), 
        .Z(SBOX_Inst_f3_dinv_2_d_5_) );
  XOR2_X2 SBOX_Inst_f3_dinv_2_U2 ( .A(SBOX_FF2_out[8]), .B(SBOX_FF2_out[14]), 
        .Z(SBOX_Inst_f3_dinv_2_d_3_) );
  XOR2_X2 SBOX_Inst_f3_dinv_2_U1 ( .A(SBOX_FF2_out[9]), .B(SBOX_FF2_out[15]), 
        .Z(SBOX_Inst_f3_dinv_2_d_2_) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U100 ( .A(SBOX_Inst_f3_dinv_2_himul_n296), 
        .B(SBOX_Inst_f3_dinv_2_himul_n295), .ZN(SBOX_Inst_f3_dinv_2_himul_n301) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_himul_U99 ( .A(SBOX_Inst_f3_dinv_2_himul_n294), 
        .B(SBOX_Inst_f3_dinv_2_himul_n293), .Z(SBOX_Inst_f3_dinv_2_himul_n295)
         );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U98 ( .A1(SBOX_Inst_f3_dinv_2_himul_n305), 
        .A2(SBOX_Inst_f3_dinv_2_d_1_), .ZN(SBOX_Inst_f3_dinv_2_himul_n296) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_himul_U97 ( .A(SBOX_Inst_f3_dinv_2_himul_n286), 
        .B(SBOX_Inst_f3_dinv_2_himul_n285), .Z(SBOX_Inst_f3_dinv_2_himul_n289)
         );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U96 ( .A1(SBOX_Inst_f3_dinv_2_d_1_), .A2(
        SBOX_FF2_out[22]), .ZN(SBOX_Inst_f3_dinv_2_himul_n285) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U95 ( .A1(SBOX_Inst_f3_dinv_2_d_0_), .A2(
        SBOX_FF2_out[23]), .ZN(SBOX_Inst_f3_dinv_2_himul_n286) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_himul_U94 ( .A(SBOX_Inst_f3_dinv_2_himul_n284), 
        .B(SBOX_Inst_f3_dinv_2_himul_n283), .Z(SBOX_Inst_f3_dinv_2_himul_n297)
         );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U93 ( .A1(SBOX_Inst_f3_dinv_2_d_1_), .A2(
        SBOX_FF2_out[18]), .ZN(SBOX_Inst_f3_dinv_2_himul_n283) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U92 ( .A1(SBOX_FF2_out[19]), .A2(
        SBOX_Inst_f3_dinv_2_d_0_), .ZN(SBOX_Inst_f3_dinv_2_himul_n284) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U91 ( .A(SBOX_Inst_f3_dinv_2_d_4_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n287) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U90 ( .A1(SBOX_Inst_f3_dinv_2_d_3_), .A2(
        SBOX_Inst_f3_dinv_2_himul_n306), .B1(SBOX_Inst_f3_dinv_2_d_2_), .B2(
        SBOX_Inst_f3_dinv_2_himul_n300), .ZN(SBOX_Inst_f3_dinv_2_himul_n298)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U89 ( .A(SBOX_Inst_f3_dinv_2_himul_n281), 
        .B(SBOX_Inst_f3_dinv_2_himul_n280), .ZN(SBOX_Inst_f3_dinv_2_pl[0]) );
  OAI22_X1 SBOX_Inst_f3_dinv_2_himul_U88 ( .A1(SBOX_Inst_f3_dinv_2_himul_n292), 
        .A2(SBOX_Inst_f3_dinv_2_d_4_), .B1(SBOX_Inst_f3_dinv_2_himul_n288), 
        .B2(SBOX_Inst_f3_dinv_2_himul_n279), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n280) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U87 ( .A1(SBOX_FF2_out[22]), .A2(
        SBOX_Inst_f3_dinv_2_d_4_), .ZN(SBOX_Inst_f3_dinv_2_himul_n279) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U86 ( .A(SBOX_Inst_f3_dinv_2_himul_n278), 
        .B(SBOX_Inst_f3_dinv_2_himul_n277), .ZN(SBOX_Inst_f3_dinv_2_himul_n281) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U85 ( .A1(SBOX_Inst_f3_dinv_2_himul_n291), 
        .A2(SBOX_Inst_f3_dinv_2_d_3_), .ZN(SBOX_Inst_f3_dinv_2_himul_n277) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U84 ( .A(SBOX_Inst_f3_dinv_2_himul_n276), 
        .B(SBOX_Inst_f3_dinv_2_himul_n275), .ZN(SBOX_Inst_f3_dinv_2_himul_n278) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U83 ( .A(SBOX_Inst_f3_dinv_2_himul_n274), 
        .B(SBOX_Inst_f3_dinv_2_himul_n273), .ZN(SBOX_Inst_f3_dinv_2_himul_n275) );
  AOI21_X1 SBOX_Inst_f3_dinv_2_himul_U82 ( .B1(SBOX_Inst_f3_dinv_2_d_4_), .B2(
        SBOX_Inst_f3_dinv_2_himul_n272), .A(SBOX_Inst_f3_dinv_2_himul_n271), 
        .ZN(SBOX_Inst_f3_dinv_2_himul_n273) );
  OAI21_X1 SBOX_Inst_f3_dinv_2_himul_U81 ( .B1(SBOX_Inst_f3_dinv_2_d_4_), .B2(
        SBOX_Inst_f3_dinv_2_himul_n272), .A(SBOX_FF2_out[21]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n271) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U80 ( .A1(SBOX_Inst_f3_dinv_2_d_5_), .A2(
        SBOX_Inst_f3_dinv_2_d_3_), .B1(SBOX_Inst_f3_dinv_2_himul_n300), .B2(
        SBOX_Inst_f3_dinv_2_himul_n288), .ZN(SBOX_Inst_f3_dinv_2_himul_n272)
         );
  OAI221_X1 SBOX_Inst_f3_dinv_2_himul_U79 ( .B1(SBOX_Inst_f3_dinv_2_d_5_), 
        .B2(SBOX_Inst_f3_dinv_2_d_2_), .C1(SBOX_Inst_f3_dinv_2_himul_n288), 
        .C2(SBOX_Inst_f3_dinv_2_himul_n306), .A(SBOX_FF2_out[20]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n274) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U78 ( .A(SBOX_Inst_f3_dinv_2_d_5_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n288) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U77 ( .A(SBOX_Inst_f3_dinv_2_himul_n269), 
        .B(SBOX_Inst_f3_dinv_2_himul_n270), .ZN(SBOX_Inst_f3_dinv_2_pl[5]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_himul_U76 ( .A(SBOX_Inst_f3_dinv_2_himul_n265), 
        .B(SBOX_Inst_f3_dinv_2_himul_n267), .Z(SBOX_Inst_f3_dinv_2_himul_n270)
         );
  AOI211_X1 SBOX_Inst_f3_dinv_2_himul_U75 ( .C1(SBOX_Inst_f3_dinv_2_d_0_), 
        .C2(SBOX_Inst_f3_dinv_2_d_3_), .A(SBOX_Inst_f3_dinv_2_himul_n268), .B(
        SBOX_Inst_f3_dinv_2_himul_n299), .ZN(SBOX_Inst_f3_dinv_2_himul_n269)
         );
  AND2_X1 SBOX_Inst_f3_dinv_2_himul_U74 ( .A1(SBOX_Inst_f3_dinv_2_himul_n304), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n300), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n268) );
  AOI211_X1 SBOX_Inst_f3_dinv_2_himul_U73 ( .C1(SBOX_FF2_out[18]), .C2(
        SBOX_FF2_out[20]), .A(SBOX_Inst_f3_dinv_2_himul_n306), .B(
        SBOX_Inst_f3_dinv_2_himul_n266), .ZN(SBOX_Inst_f3_dinv_2_himul_n267)
         );
  AND2_X1 SBOX_Inst_f3_dinv_2_himul_U72 ( .A1(SBOX_Inst_f3_dinv_2_himul_n307), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n308), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n266) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U71 ( .A(SBOX_Inst_f3_dinv_2_himul_n263), 
        .B(SBOX_Inst_f3_dinv_2_himul_n264), .ZN(SBOX_Inst_f3_dinv_2_himul_n265) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U70 ( .A1(SBOX_Inst_f3_dinv_2_himul_n303), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n302), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n264) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U69 ( .A(SBOX_Inst_f3_dinv_2_himul_n301), 
        .B(SBOX_Inst_f3_dinv_2_himul_n262), .ZN(SBOX_Inst_f3_dinv_2_himul_n263) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U68 ( .A1(SBOX_FF2_out[19]), .A2(
        SBOX_Inst_f3_dinv_2_himul_n304), .B1(SBOX_Inst_f3_dinv_2_d_0_), .B2(
        SBOX_Inst_f3_dinv_2_himul_n305), .ZN(SBOX_Inst_f3_dinv_2_himul_n262)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U67 ( .A(SBOX_Inst_f3_dinv_2_himul_n261), 
        .B(SBOX_Inst_f3_dinv_2_himul_n260), .ZN(SBOX_Inst_f3_dinv_2_pl[4]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U66 ( .A(SBOX_Inst_f3_dinv_2_himul_n297), 
        .B(SBOX_Inst_f3_dinv_2_himul_n257), .ZN(SBOX_Inst_f3_dinv_2_himul_n261) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U65 ( .A(SBOX_Inst_f3_dinv_2_himul_n258), 
        .B(SBOX_Inst_f3_dinv_2_himul_n259), .ZN(SBOX_Inst_f3_dinv_2_himul_n260) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U64 ( .A1(SBOX_Inst_f3_dinv_2_d_3_), .A2(
        SBOX_Inst_f3_dinv_2_himul_n302), .ZN(SBOX_Inst_f3_dinv_2_himul_n259)
         );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U63 ( .A1(SBOX_Inst_f3_dinv_2_himul_n308), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n298), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n258) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U62 ( .A(SBOX_Inst_f3_dinv_2_himul_n301), 
        .B(SBOX_Inst_f3_dinv_2_himul_n256), .ZN(SBOX_Inst_f3_dinv_2_himul_n257) );
  MUX2_X1 SBOX_Inst_f3_dinv_2_himul_U61 ( .A(SBOX_Inst_f3_dinv_2_d_0_), .B(
        SBOX_Inst_f3_dinv_2_d_1_), .S(SBOX_Inst_f3_dinv_2_himul_n255), .Z(
        SBOX_Inst_f3_dinv_2_himul_n256) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U60 ( .A1(SBOX_FF2_out[21]), .A2(
        SBOX_FF2_out[19]), .B1(SBOX_Inst_f3_dinv_2_himul_n302), .B2(
        SBOX_Inst_f3_dinv_2_himul_n299), .ZN(SBOX_Inst_f3_dinv_2_himul_n255)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U59 ( .A(SBOX_Inst_f3_dinv_2_himul_n254), 
        .B(SBOX_Inst_f3_dinv_2_himul_n253), .ZN(SBOX_Inst_f3_dinv_2_pl[3]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U58 ( .A(SBOX_Inst_f3_dinv_2_himul_n249), 
        .B(SBOX_Inst_f3_dinv_2_himul_n251), .ZN(SBOX_Inst_f3_dinv_2_himul_n254) );
  OAI221_X1 SBOX_Inst_f3_dinv_2_himul_U57 ( .B1(SBOX_Inst_f3_dinv_2_himul_n243), .B2(SBOX_FF2_out[19]), .C1(SBOX_Inst_f3_dinv_2_himul_n252), .C2(
        SBOX_Inst_f3_dinv_2_himul_n302), .A(SBOX_Inst_f3_dinv_2_d_4_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n253) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U56 ( .A(SBOX_Inst_f3_dinv_2_himul_n243), 
        .ZN(SBOX_Inst_f3_dinv_2_himul_n252) );
  OAI21_X1 SBOX_Inst_f3_dinv_2_himul_U55 ( .B1(SBOX_Inst_f3_dinv_2_himul_n292), 
        .B2(SBOX_Inst_f3_dinv_2_himul_n291), .A(SBOX_Inst_f3_dinv_2_himul_n250), .ZN(SBOX_Inst_f3_dinv_2_himul_n251) );
  NAND3_X1 SBOX_Inst_f3_dinv_2_himul_U54 ( .A1(SBOX_Inst_f3_dinv_2_himul_n292), 
        .A2(SBOX_FF2_out[22]), .A3(SBOX_Inst_f3_dinv_2_himul_n290), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n250) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U53 ( .A(SBOX_Inst_f3_dinv_2_himul_n247), 
        .B(SBOX_Inst_f3_dinv_2_himul_n248), .ZN(SBOX_Inst_f3_dinv_2_himul_n249) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U52 ( .A1(SBOX_Inst_f3_dinv_2_himul_n243), 
        .A2(SBOX_Inst_f3_dinv_2_d_5_), .ZN(SBOX_Inst_f3_dinv_2_himul_n248) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_himul_U51 ( .A(SBOX_Inst_f3_dinv_2_himul_n289), 
        .B(SBOX_Inst_f3_dinv_2_himul_n246), .Z(SBOX_Inst_f3_dinv_2_himul_n247)
         );
  XOR2_X1 SBOX_Inst_f3_dinv_2_himul_U50 ( .A(SBOX_Inst_f3_dinv_2_himul_n244), 
        .B(SBOX_Inst_f3_dinv_2_himul_n245), .Z(SBOX_Inst_f3_dinv_2_himul_n246)
         );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U49 ( .A1(SBOX_Inst_f3_dinv_2_d_0_), .A2(
        SBOX_FF2_out[22]), .ZN(SBOX_Inst_f3_dinv_2_himul_n245) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U48 ( .A1(SBOX_Inst_f3_dinv_2_himul_n303), 
        .A2(SBOX_FF2_out[19]), .ZN(SBOX_Inst_f3_dinv_2_himul_n244) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U47 ( .A1(SBOX_FF2_out[23]), .A2(
        SBOX_FF2_out[18]), .B1(SBOX_Inst_f3_dinv_2_himul_n290), .B2(
        SBOX_Inst_f3_dinv_2_himul_n307), .ZN(SBOX_Inst_f3_dinv_2_himul_n243)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U46 ( .A(SBOX_Inst_f3_dinv_2_himul_n297), 
        .B(SBOX_Inst_f3_dinv_2_himul_n242), .ZN(SBOX_Inst_f3_dinv_2_pl[2]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U45 ( .A(SBOX_Inst_f3_dinv_2_himul_n240), 
        .B(SBOX_Inst_f3_dinv_2_himul_n241), .ZN(SBOX_Inst_f3_dinv_2_himul_n242) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U44 ( .A1(SBOX_FF2_out[18]), .A2(
        SBOX_Inst_f3_dinv_2_d_5_), .ZN(SBOX_Inst_f3_dinv_2_himul_n241) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_himul_U43 ( .A(SBOX_Inst_f3_dinv_2_himul_n239), 
        .B(SBOX_Inst_f3_dinv_2_himul_n289), .Z(SBOX_Inst_f3_dinv_2_himul_n240)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U42 ( .A(SBOX_Inst_f3_dinv_2_himul_n237), 
        .B(SBOX_Inst_f3_dinv_2_himul_n238), .ZN(SBOX_Inst_f3_dinv_2_himul_n239) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U41 ( .A(SBOX_Inst_f3_dinv_2_himul_n234), 
        .B(SBOX_Inst_f3_dinv_2_himul_n235), .ZN(SBOX_Inst_f3_dinv_2_himul_n238) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U40 ( .A1(SBOX_Inst_f3_dinv_2_himul_n231), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n236), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n237) );
  OAI22_X1 SBOX_Inst_f3_dinv_2_himul_U39 ( .A1(SBOX_Inst_f3_dinv_2_d_4_), .A2(
        SBOX_Inst_f3_dinv_2_d_5_), .B1(SBOX_Inst_f3_dinv_2_himul_n288), .B2(
        SBOX_Inst_f3_dinv_2_himul_n287), .ZN(SBOX_Inst_f3_dinv_2_himul_n236)
         );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U38 ( .A1(SBOX_FF2_out[19]), .A2(
        SBOX_Inst_f3_dinv_2_d_0_), .B1(SBOX_Inst_f3_dinv_2_himul_n302), .B2(
        SBOX_Inst_f3_dinv_2_himul_n304), .ZN(SBOX_Inst_f3_dinv_2_himul_n235)
         );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U37 ( .A1(SBOX_FF2_out[23]), .A2(
        SBOX_Inst_f3_dinv_2_himul_n232), .B1(SBOX_Inst_f3_dinv_2_d_4_), .B2(
        SBOX_Inst_f3_dinv_2_himul_n233), .ZN(SBOX_Inst_f3_dinv_2_himul_n234)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U36 ( .A(SBOX_FF2_out[23]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n233) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U35 ( .A1(SBOX_Inst_f3_dinv_2_d_1_), .A2(
        SBOX_Inst_f3_dinv_2_d_5_), .B1(SBOX_Inst_f3_dinv_2_himul_n288), .B2(
        SBOX_Inst_f3_dinv_2_himul_n303), .ZN(SBOX_Inst_f3_dinv_2_himul_n232)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U34 ( .A(SBOX_FF2_out[19]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n231) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U33 ( .A(SBOX_Inst_f3_dinv_2_himul_n228), 
        .B(SBOX_Inst_f3_dinv_2_himul_n230), .ZN(SBOX_Inst_f3_dinv_2_pl[1]) );
  AOI211_X1 SBOX_Inst_f3_dinv_2_himul_U32 ( .C1(SBOX_FF2_out[22]), .C2(
        SBOX_FF2_out[20]), .A(SBOX_Inst_f3_dinv_2_himul_n298), .B(
        SBOX_Inst_f3_dinv_2_himul_n229), .ZN(SBOX_Inst_f3_dinv_2_himul_n230)
         );
  AND2_X1 SBOX_Inst_f3_dinv_2_himul_U31 ( .A1(SBOX_Inst_f3_dinv_2_himul_n282), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n308), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n229) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U30 ( .A(SBOX_Inst_f3_dinv_2_himul_n227), 
        .B(SBOX_Inst_f3_dinv_2_himul_n224), .ZN(SBOX_Inst_f3_dinv_2_himul_n228) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U29 ( .A1(SBOX_Inst_f3_dinv_2_himul_n226), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n225), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n227) );
  OAI22_X1 SBOX_Inst_f3_dinv_2_himul_U28 ( .A1(SBOX_FF2_out[21]), .A2(
        SBOX_FF2_out[22]), .B1(SBOX_Inst_f3_dinv_2_himul_n282), .B2(
        SBOX_Inst_f3_dinv_2_himul_n299), .ZN(SBOX_Inst_f3_dinv_2_himul_n226)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U27 ( .A(SBOX_Inst_f3_dinv_2_d_4_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n225) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U26 ( .A(SBOX_Inst_f3_dinv_2_himul_n222), 
        .B(SBOX_Inst_f3_dinv_2_himul_n223), .ZN(SBOX_Inst_f3_dinv_2_himul_n224) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U25 ( .A(SBOX_FF2_out[22]), .B(
        SBOX_Inst_f3_dinv_2_himul_n220), .ZN(SBOX_Inst_f3_dinv_2_himul_n223)
         );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U24 ( .A1(SBOX_Inst_f3_dinv_2_himul_n215), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n221), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n222) );
  OAI22_X1 SBOX_Inst_f3_dinv_2_himul_U23 ( .A1(SBOX_Inst_f3_dinv_2_d_2_), .A2(
        SBOX_Inst_f3_dinv_2_d_3_), .B1(SBOX_Inst_f3_dinv_2_himul_n306), .B2(
        SBOX_Inst_f3_dinv_2_himul_n300), .ZN(SBOX_Inst_f3_dinv_2_himul_n221)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_himul_U22 ( .A(SBOX_Inst_f3_dinv_2_himul_n219), 
        .B(SBOX_Inst_f3_dinv_2_himul_n218), .ZN(SBOX_Inst_f3_dinv_2_himul_n220) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U21 ( .A1(SBOX_Inst_f3_dinv_2_himul_n216), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n290), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n219) );
  OAI221_X1 SBOX_Inst_f3_dinv_2_himul_U20 ( .B1(SBOX_Inst_f3_dinv_2_himul_n216), .B2(SBOX_Inst_f3_dinv_2_d_4_), .C1(SBOX_Inst_f3_dinv_2_himul_n217), .C2(
        SBOX_Inst_f3_dinv_2_himul_n287), .A(SBOX_FF2_out[20]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n218) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U19 ( .A(SBOX_Inst_f3_dinv_2_himul_n216), 
        .ZN(SBOX_Inst_f3_dinv_2_himul_n217) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U18 ( .A1(SBOX_Inst_f3_dinv_2_d_5_), .A2(
        SBOX_Inst_f3_dinv_2_d_2_), .B1(SBOX_Inst_f3_dinv_2_himul_n306), .B2(
        SBOX_Inst_f3_dinv_2_himul_n288), .ZN(SBOX_Inst_f3_dinv_2_himul_n216)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U17 ( .A(SBOX_FF2_out[21]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n215) );
  OAI221_X1 SBOX_Inst_f3_dinv_2_himul_U16 ( .B1(SBOX_FF2_out[21]), .B2(
        SBOX_FF2_out[23]), .C1(SBOX_Inst_f3_dinv_2_himul_n299), .C2(
        SBOX_Inst_f3_dinv_2_himul_n290), .A(SBOX_Inst_f3_dinv_2_d_2_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n276) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U15 ( .A(SBOX_FF2_out[19]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n302) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U14 ( .A(SBOX_FF2_out[20]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n308) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U13 ( .A1(SBOX_FF2_out[18]), .A2(
        SBOX_Inst_f3_dinv_2_d_3_), .ZN(SBOX_Inst_f3_dinv_2_himul_n293) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_himul_U12 ( .A1(SBOX_FF2_out[19]), .A2(
        SBOX_Inst_f3_dinv_2_d_2_), .ZN(SBOX_Inst_f3_dinv_2_himul_n294) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U11 ( .A(SBOX_FF2_out[21]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n299) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U10 ( .A(SBOX_Inst_f3_dinv_2_d_0_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n304) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U9 ( .A(SBOX_Inst_f3_dinv_2_d_3_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n300) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U8 ( .A(SBOX_Inst_f3_dinv_2_d_2_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n306) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U7 ( .A1(SBOX_FF2_out[20]), .A2(
        SBOX_FF2_out[18]), .B1(SBOX_Inst_f3_dinv_2_himul_n307), .B2(
        SBOX_Inst_f3_dinv_2_himul_n308), .ZN(SBOX_Inst_f3_dinv_2_himul_n305)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U6 ( .A(SBOX_FF2_out[18]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n307) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U5 ( .A(SBOX_Inst_f3_dinv_2_d_1_), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n303) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_himul_U4 ( .A1(SBOX_Inst_f3_dinv_2_himul_n282), 
        .A2(SBOX_Inst_f3_dinv_2_himul_n288), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n292) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_himul_U3 ( .A1(SBOX_FF2_out[22]), .A2(
        SBOX_FF2_out[23]), .B1(SBOX_Inst_f3_dinv_2_himul_n290), .B2(
        SBOX_Inst_f3_dinv_2_himul_n282), .ZN(SBOX_Inst_f3_dinv_2_himul_n291)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U2 ( .A(SBOX_FF2_out[23]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n290) );
  INV_X1 SBOX_Inst_f3_dinv_2_himul_U1 ( .A(SBOX_FF2_out[22]), .ZN(
        SBOX_Inst_f3_dinv_2_himul_n282) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U100 ( .A1(SBOX_Inst_f3_dinv_2_d_2_), 
        .A2(SBOX_Inst_f3_dinv_2_d_0_), .B1(SBOX_Inst_f3_dinv_2_lowmul_n307), 
        .B2(SBOX_Inst_f3_dinv_2_lowmul_n308), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n305) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U99 ( .A(SBOX_Inst_f3_dinv_2_d_0_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n307) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U98 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n292), .B(SBOX_Inst_f3_dinv_2_lowmul_n291), .ZN(SBOX_Inst_f3_dinv_2_ph[2]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U97 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n290), .B(SBOX_Inst_f3_dinv_2_lowmul_n289), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n291) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U96 ( .A1(SBOX_Inst_f3_dinv_2_d_0_), 
        .A2(SBOX_FF2_out[5]), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n289) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U95 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n288), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n287), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n290) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U94 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n286), .B(SBOX_Inst_f3_dinv_2_lowmul_n285), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n287) );
  MUX2_X1 SBOX_Inst_f3_dinv_2_lowmul_U93 ( .A(SBOX_FF2_out[4]), .B(
        SBOX_Inst_f3_dinv_2_lowmul_n284), .S(SBOX_Inst_f3_dinv_2_d_5_), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n285) );
  OAI221_X1 SBOX_Inst_f3_dinv_2_lowmul_U92 ( .B1(SBOX_FF2_out[5]), .B2(
        SBOX_FF2_out[4]), .C1(SBOX_Inst_f3_dinv_2_lowmul_n283), .C2(
        SBOX_Inst_f3_dinv_2_lowmul_n282), .A(SBOX_Inst_f3_dinv_2_d_1_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n286) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U91 ( .A1(SBOX_Inst_f3_dinv_2_d_1_), 
        .A2(SBOX_FF2_out[0]), .B1(SBOX_Inst_f3_dinv_2_lowmul_n304), .B2(
        SBOX_Inst_f3_dinv_2_lowmul_n302), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n288)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U90 ( .A(SBOX_Inst_f3_dinv_2_d_1_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n302) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U89 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n281), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n280), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n293) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U88 ( .A1(SBOX_FF2_out[1]), .A2(
        SBOX_Inst_f3_dinv_2_d_4_), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n280) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U87 ( .A1(SBOX_FF2_out[0]), .A2(
        SBOX_Inst_f3_dinv_2_d_5_), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n281) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U86 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n279), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n278), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n297) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U85 ( .A1(SBOX_FF2_out[1]), .A2(
        SBOX_Inst_f3_dinv_2_d_0_), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n278) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U84 ( .A1(SBOX_Inst_f3_dinv_2_d_1_), 
        .A2(SBOX_FF2_out[0]), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n279) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U83 ( .A(SBOX_Inst_f3_dinv_2_d_2_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n308) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U82 ( .A1(SBOX_Inst_f3_dinv_2_d_4_), 
        .A2(SBOX_Inst_f3_dinv_2_d_5_), .B1(SBOX_Inst_f3_dinv_2_lowmul_n294), 
        .B2(SBOX_Inst_f3_dinv_2_lowmul_n277), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n295) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U81 ( .A(SBOX_Inst_f3_dinv_2_d_4_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n277) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U80 ( .A(SBOX_Inst_f3_dinv_2_d_3_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n299) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U79 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n274), .B(SBOX_Inst_f3_dinv_2_lowmul_n276), .ZN(SBOX_Inst_f3_dinv_2_ph[1]) );
  AOI211_X1 SBOX_Inst_f3_dinv_2_lowmul_U78 ( .C1(SBOX_Inst_f3_dinv_2_d_4_), 
        .C2(SBOX_Inst_f3_dinv_2_d_2_), .A(SBOX_Inst_f3_dinv_2_lowmul_n298), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n275), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n276) );
  AND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U77 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n277), .A2(SBOX_Inst_f3_dinv_2_lowmul_n308), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n275)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U76 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n273), .B(SBOX_Inst_f3_dinv_2_lowmul_n270), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n274) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U75 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n272), .A2(SBOX_Inst_f3_dinv_2_lowmul_n271), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n273)
         );
  OAI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U74 ( .A1(SBOX_Inst_f3_dinv_2_d_3_), 
        .A2(SBOX_Inst_f3_dinv_2_d_4_), .B1(SBOX_Inst_f3_dinv_2_lowmul_n277), 
        .B2(SBOX_Inst_f3_dinv_2_lowmul_n299), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n272) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U73 ( .A(SBOX_FF2_out[4]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n271) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U72 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n268), .B(SBOX_Inst_f3_dinv_2_lowmul_n269), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n270) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U71 ( .A(SBOX_Inst_f3_dinv_2_d_4_), .B(
        SBOX_Inst_f3_dinv_2_lowmul_n266), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n269)
         );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U70 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n261), .A2(SBOX_Inst_f3_dinv_2_lowmul_n267), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n268)
         );
  OAI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U69 ( .A1(SBOX_FF2_out[2]), .A2(
        SBOX_FF2_out[3]), .B1(SBOX_Inst_f3_dinv_2_lowmul_n306), .B2(
        SBOX_Inst_f3_dinv_2_lowmul_n300), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n267)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U68 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n265), .B(SBOX_Inst_f3_dinv_2_lowmul_n264), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n266) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U67 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n262), .A2(SBOX_Inst_f3_dinv_2_lowmul_n294), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n265)
         );
  OAI221_X1 SBOX_Inst_f3_dinv_2_lowmul_U66 ( .B1(
        SBOX_Inst_f3_dinv_2_lowmul_n262), .B2(SBOX_FF2_out[4]), .C1(
        SBOX_Inst_f3_dinv_2_lowmul_n263), .C2(SBOX_Inst_f3_dinv_2_lowmul_n282), 
        .A(SBOX_Inst_f3_dinv_2_d_2_), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n264) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U65 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n262), 
        .ZN(SBOX_Inst_f3_dinv_2_lowmul_n263) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U64 ( .A1(SBOX_FF2_out[5]), .A2(
        SBOX_FF2_out[2]), .B1(SBOX_Inst_f3_dinv_2_lowmul_n306), .B2(
        SBOX_Inst_f3_dinv_2_lowmul_n283), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n262)
         );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U63 ( .A(SBOX_Inst_f3_dinv_2_d_3_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n261) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U62 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n260), .B(SBOX_Inst_f3_dinv_2_lowmul_n259), .ZN(SBOX_Inst_f3_dinv_2_ph[4]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U61 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n297), .B(SBOX_Inst_f3_dinv_2_lowmul_n256), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n260) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U60 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n257), .B(SBOX_Inst_f3_dinv_2_lowmul_n258), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n259) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U59 ( .A1(SBOX_FF2_out[3]), .A2(
        SBOX_Inst_f3_dinv_2_lowmul_n302), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n258)
         );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U58 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n308), .A2(SBOX_Inst_f3_dinv_2_lowmul_n298), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n257)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U57 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n301), .B(SBOX_Inst_f3_dinv_2_lowmul_n255), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n256) );
  MUX2_X1 SBOX_Inst_f3_dinv_2_lowmul_U56 ( .A(SBOX_FF2_out[0]), .B(
        SBOX_FF2_out[1]), .S(SBOX_Inst_f3_dinv_2_lowmul_n254), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n255) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U55 ( .A1(SBOX_Inst_f3_dinv_2_d_3_), 
        .A2(SBOX_Inst_f3_dinv_2_d_1_), .B1(SBOX_Inst_f3_dinv_2_lowmul_n302), 
        .B2(SBOX_Inst_f3_dinv_2_lowmul_n299), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n254) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U54 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n252), .B(SBOX_Inst_f3_dinv_2_lowmul_n253), .ZN(SBOX_Inst_f3_dinv_2_ph[5]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U53 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n248), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n250), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n253) );
  AOI211_X1 SBOX_Inst_f3_dinv_2_lowmul_U52 ( .C1(SBOX_FF2_out[0]), .C2(
        SBOX_FF2_out[3]), .A(SBOX_Inst_f3_dinv_2_lowmul_n251), .B(
        SBOX_Inst_f3_dinv_2_lowmul_n299), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n252)
         );
  AND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U51 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n304), .A2(SBOX_Inst_f3_dinv_2_lowmul_n300), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n251)
         );
  AOI211_X1 SBOX_Inst_f3_dinv_2_lowmul_U50 ( .C1(SBOX_Inst_f3_dinv_2_d_0_), 
        .C2(SBOX_Inst_f3_dinv_2_d_2_), .A(SBOX_Inst_f3_dinv_2_lowmul_n306), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n249), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n250) );
  AND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U49 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n307), .A2(SBOX_Inst_f3_dinv_2_lowmul_n308), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n249)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U48 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n246), .B(SBOX_Inst_f3_dinv_2_lowmul_n247), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n248) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U47 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n303), .A2(SBOX_Inst_f3_dinv_2_lowmul_n302), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n247)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U46 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n301), .B(SBOX_Inst_f3_dinv_2_lowmul_n245), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n246) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U45 ( .A1(SBOX_Inst_f3_dinv_2_d_1_), 
        .A2(SBOX_Inst_f3_dinv_2_lowmul_n304), .B1(SBOX_FF2_out[0]), .B2(
        SBOX_Inst_f3_dinv_2_lowmul_n305), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n245)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U44 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n241), .B(SBOX_Inst_f3_dinv_2_lowmul_n244), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n301) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U43 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n242), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n243), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n244) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U42 ( .A1(SBOX_FF2_out[3]), .A2(
        SBOX_Inst_f3_dinv_2_d_0_), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n243) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U41 ( .A1(SBOX_Inst_f3_dinv_2_d_1_), 
        .A2(SBOX_FF2_out[2]), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n242) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U40 ( .A1(
        SBOX_Inst_f3_dinv_2_lowmul_n305), .A2(SBOX_FF2_out[1]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n241) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U39 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n240), .B(SBOX_Inst_f3_dinv_2_lowmul_n239), .ZN(SBOX_Inst_f3_dinv_2_ph[3]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U38 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n235), .B(SBOX_Inst_f3_dinv_2_lowmul_n237), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n240) );
  OAI221_X1 SBOX_Inst_f3_dinv_2_lowmul_U37 ( .B1(
        SBOX_Inst_f3_dinv_2_lowmul_n229), .B2(SBOX_Inst_f3_dinv_2_d_1_), .C1(
        SBOX_Inst_f3_dinv_2_lowmul_n238), .C2(SBOX_Inst_f3_dinv_2_lowmul_n302), 
        .A(SBOX_FF2_out[4]), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n239) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U36 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n229), 
        .ZN(SBOX_Inst_f3_dinv_2_lowmul_n238) );
  OAI21_X1 SBOX_Inst_f3_dinv_2_lowmul_U35 ( .B1(
        SBOX_Inst_f3_dinv_2_lowmul_n296), .B2(SBOX_Inst_f3_dinv_2_lowmul_n295), 
        .A(SBOX_Inst_f3_dinv_2_lowmul_n236), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n237) );
  NAND3_X1 SBOX_Inst_f3_dinv_2_lowmul_U34 ( .A1(
        SBOX_Inst_f3_dinv_2_lowmul_n296), .A2(SBOX_Inst_f3_dinv_2_d_4_), .A3(
        SBOX_Inst_f3_dinv_2_lowmul_n294), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n236)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U33 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n233), .B(SBOX_Inst_f3_dinv_2_lowmul_n234), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n235) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U32 ( .A1(
        SBOX_Inst_f3_dinv_2_lowmul_n229), .A2(SBOX_FF2_out[5]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n234) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U31 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n293), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n232), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n233) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U30 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n230), 
        .B(SBOX_Inst_f3_dinv_2_lowmul_n231), .Z(
        SBOX_Inst_f3_dinv_2_lowmul_n232) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U29 ( .A1(SBOX_FF2_out[0]), .A2(
        SBOX_Inst_f3_dinv_2_d_4_), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n231) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U28 ( .A1(
        SBOX_Inst_f3_dinv_2_lowmul_n303), .A2(SBOX_Inst_f3_dinv_2_d_1_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n230) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U27 ( .A1(SBOX_Inst_f3_dinv_2_d_5_), 
        .A2(SBOX_Inst_f3_dinv_2_d_0_), .B1(SBOX_Inst_f3_dinv_2_lowmul_n294), 
        .B2(SBOX_Inst_f3_dinv_2_lowmul_n307), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n229) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U26 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n226), .B(SBOX_Inst_f3_dinv_2_lowmul_n228), .ZN(SBOX_Inst_f3_dinv_2_ph[0]) );
  OAI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U25 ( .A1(
        SBOX_Inst_f3_dinv_2_lowmul_n283), .A2(SBOX_Inst_f3_dinv_2_lowmul_n227), 
        .B1(SBOX_Inst_f3_dinv_2_lowmul_n296), .B2(SBOX_FF2_out[4]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n228) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U24 ( .A1(SBOX_FF2_out[4]), .A2(
        SBOX_Inst_f3_dinv_2_d_4_), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n227) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U23 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n225), .B(SBOX_Inst_f3_dinv_2_lowmul_n224), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n226) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U22 ( .A1(
        SBOX_Inst_f3_dinv_2_lowmul_n295), .A2(SBOX_FF2_out[3]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n225) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U21 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n223), .B(SBOX_Inst_f3_dinv_2_lowmul_n217), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n224) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U20 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n222), .B(SBOX_Inst_f3_dinv_2_lowmul_n219), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n223) );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U19 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n221), .A2(SBOX_Inst_f3_dinv_2_lowmul_n220), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n222)
         );
  OAI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U18 ( .A1(SBOX_Inst_f3_dinv_2_d_5_), 
        .A2(SBOX_Inst_f3_dinv_2_d_3_), .B1(SBOX_Inst_f3_dinv_2_lowmul_n294), 
        .B2(SBOX_Inst_f3_dinv_2_lowmul_n299), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n221) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U17 ( .A(SBOX_FF2_out[2]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n220) );
  OAI211_X1 SBOX_Inst_f3_dinv_2_lowmul_U16 ( .C1(SBOX_FF2_out[2]), .C2(
        SBOX_FF2_out[5]), .A(SBOX_Inst_f3_dinv_2_d_2_), .B(
        SBOX_Inst_f3_dinv_2_lowmul_n218), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n219)
         );
  OR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U15 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n283), 
        .A2(SBOX_Inst_f3_dinv_2_lowmul_n306), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n218) );
  OAI211_X1 SBOX_Inst_f3_dinv_2_lowmul_U14 ( .C1(
        SBOX_Inst_f3_dinv_2_lowmul_n215), .C2(SBOX_FF2_out[4]), .A(
        SBOX_Inst_f3_dinv_2_d_3_), .B(SBOX_Inst_f3_dinv_2_lowmul_n216), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n217) );
  NAND2_X1 SBOX_Inst_f3_dinv_2_lowmul_U13 ( .A1(
        SBOX_Inst_f3_dinv_2_lowmul_n215), .A2(SBOX_FF2_out[4]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n216) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U12 ( .A1(SBOX_FF2_out[3]), .A2(
        SBOX_FF2_out[5]), .B1(SBOX_Inst_f3_dinv_2_lowmul_n283), .B2(
        SBOX_Inst_f3_dinv_2_lowmul_n300), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n215)
         );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U11 ( .A1(SBOX_FF2_out[5]), .A2(
        SBOX_FF2_out[1]), .B1(SBOX_Inst_f3_dinv_2_lowmul_n303), .B2(
        SBOX_Inst_f3_dinv_2_lowmul_n283), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n284)
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U10 ( .A(SBOX_Inst_f3_dinv_2_lowmul_n297), .B(SBOX_Inst_f3_dinv_2_lowmul_n293), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n292) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U9 ( .A(SBOX_FF2_out[3]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n300) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U8 ( .A(SBOX_FF2_out[2]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n306) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U7 ( .A(SBOX_FF2_out[0]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n304) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U6 ( .A(SBOX_FF2_out[1]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n303) );
  AOI22_X1 SBOX_Inst_f3_dinv_2_lowmul_U5 ( .A1(SBOX_FF2_out[3]), .A2(
        SBOX_Inst_f3_dinv_2_lowmul_n306), .B1(SBOX_FF2_out[2]), .B2(
        SBOX_Inst_f3_dinv_2_lowmul_n300), .ZN(SBOX_Inst_f3_dinv_2_lowmul_n298)
         );
  NOR2_X1 SBOX_Inst_f3_dinv_2_lowmul_U4 ( .A1(SBOX_Inst_f3_dinv_2_lowmul_n277), 
        .A2(SBOX_Inst_f3_dinv_2_lowmul_n283), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n296) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U3 ( .A(SBOX_Inst_f3_dinv_2_d_5_), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n294) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U2 ( .A(SBOX_FF2_out[5]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n283) );
  INV_X1 SBOX_Inst_f3_dinv_2_lowmul_U1 ( .A(SBOX_FF2_out[4]), .ZN(
        SBOX_Inst_f3_dinv_2_lowmul_n282) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U16 ( .A(PRNGQ[26]), .B(
        SBOX_Inst_f3_dinv_2_ph[2]), .Z(SBOX_muld[6]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U15 ( .A(PRNGQ[20]), .B(
        SBOX_Inst_f3_dinv_2_pl[0]), .Z(SBOX_muld[0]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U14 ( .A(PRNGQ[25]), .B(
        SBOX_Inst_f3_dinv_2_ph[1]), .Z(SBOX_muld[3]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U13 ( .A(
        SBOX_Inst_f3_dinv_2_AddNewMaskQ_n4), .B(SBOX_Inst_f3_dinv_2_ph[4]), 
        .ZN(SBOX_muld[10]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U12 ( .A(PRNGQ[26]), .B(PRNGQ[24]), 
        .ZN(SBOX_Inst_f3_dinv_2_AddNewMaskQ_n4) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U11 ( .A(
        SBOX_Inst_f3_dinv_2_AddNewMaskQ_n3), .B(SBOX_Inst_f3_dinv_2_ph[5]), 
        .ZN(SBOX_muld[11]) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U10 ( .A(PRNGQ[27]), .B(PRNGQ[25]), 
        .ZN(SBOX_Inst_f3_dinv_2_AddNewMaskQ_n3) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U9 ( .A(
        SBOX_Inst_f3_dinv_2_AddNewMaskQ_n2), .B(PRNGQ[23]), .ZN(SBOX_muld[9])
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U8 ( .A(PRNGQ[21]), .B(
        SBOX_Inst_f3_dinv_2_pl[5]), .ZN(SBOX_Inst_f3_dinv_2_AddNewMaskQ_n2) );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U7 ( .A(
        SBOX_Inst_f3_dinv_2_AddNewMaskQ_n1), .B(PRNGQ[22]), .ZN(SBOX_muld[8])
         );
  XNOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U6 ( .A(PRNGQ[20]), .B(
        SBOX_Inst_f3_dinv_2_pl[4]), .ZN(SBOX_Inst_f3_dinv_2_AddNewMaskQ_n1) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U5 ( .A(PRNGQ[27]), .B(
        SBOX_Inst_f3_dinv_2_ph[3]), .Z(SBOX_muld[7]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U4 ( .A(PRNGQ[23]), .B(
        SBOX_Inst_f3_dinv_2_pl[3]), .Z(SBOX_muld[5]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U3 ( .A(PRNGQ[22]), .B(
        SBOX_Inst_f3_dinv_2_pl[2]), .Z(SBOX_muld[4]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U2 ( .A(PRNGQ[24]), .B(
        SBOX_Inst_f3_dinv_2_ph[0]), .Z(SBOX_muld[2]) );
  XOR2_X1 SBOX_Inst_f3_dinv_2_AddNewMaskQ_U1 ( .A(PRNGQ[21]), .B(
        SBOX_Inst_f3_dinv_2_pl[1]), .Z(SBOX_muld[1]) );
  OAI21_X1 SBOX_PL_3_U73 ( .B1(1'b1), .B2(SBOX_PL_3_n180), .A(SBOX_PL_3_n252), 
        .ZN(SBOX_PL_3_n144) );
  NAND2_X1 SBOX_PL_3_U72 ( .A1(1'b1), .A2(SBOX_muld[0]), .ZN(SBOX_PL_3_n252)
         );
  OAI21_X1 SBOX_PL_3_U71 ( .B1(1'b1), .B2(SBOX_PL_3_n174), .A(SBOX_PL_3_n251), 
        .ZN(SBOX_PL_3_n138) );
  NAND2_X1 SBOX_PL_3_U70 ( .A1(1'b1), .A2(SBOX_muld[6]), .ZN(SBOX_PL_3_n251)
         );
  OAI21_X1 SBOX_PL_3_U69 ( .B1(1'b1), .B2(SBOX_PL_3_n168), .A(SBOX_PL_3_n250), 
        .ZN(SBOX_PL_3_n132) );
  NAND2_X1 SBOX_PL_3_U68 ( .A1(1'b1), .A2(SBOX_Zl_f3[0]), .ZN(SBOX_PL_3_n250)
         );
  OAI21_X1 SBOX_PL_3_U67 ( .B1(1'b1), .B2(SBOX_PL_3_n167), .A(SBOX_PL_3_n249), 
        .ZN(SBOX_PL_3_n131) );
  NAND2_X1 SBOX_PL_3_U66 ( .A1(1'b1), .A2(SBOX_Zl_f3[1]), .ZN(SBOX_PL_3_n249)
         );
  OAI21_X1 SBOX_PL_3_U65 ( .B1(1'b1), .B2(SBOX_PL_3_n166), .A(SBOX_PL_3_n248), 
        .ZN(SBOX_PL_3_n130) );
  NAND2_X1 SBOX_PL_3_U64 ( .A1(1'b1), .A2(SBOX_Zl_f3[2]), .ZN(SBOX_PL_3_n248)
         );
  OAI21_X1 SBOX_PL_3_U63 ( .B1(1'b1), .B2(SBOX_PL_3_n165), .A(SBOX_PL_3_n247), 
        .ZN(SBOX_PL_3_n129) );
  NAND2_X1 SBOX_PL_3_U62 ( .A1(1'b1), .A2(SBOX_Zl_f3[3]), .ZN(SBOX_PL_3_n247)
         );
  OAI21_X1 SBOX_PL_3_U61 ( .B1(1'b1), .B2(SBOX_PL_3_n164), .A(SBOX_PL_3_n246), 
        .ZN(SBOX_PL_3_n128) );
  NAND2_X1 SBOX_PL_3_U60 ( .A1(1'b1), .A2(SBOX_Zl_f3[4]), .ZN(SBOX_PL_3_n246)
         );
  OAI21_X1 SBOX_PL_3_U59 ( .B1(1'b1), .B2(SBOX_PL_3_n163), .A(SBOX_PL_3_n245), 
        .ZN(SBOX_PL_3_n127) );
  NAND2_X1 SBOX_PL_3_U58 ( .A1(1'b1), .A2(SBOX_Zl_f3[5]), .ZN(SBOX_PL_3_n245)
         );
  OAI21_X1 SBOX_PL_3_U57 ( .B1(1'b1), .B2(SBOX_PL_3_n162), .A(SBOX_PL_3_n244), 
        .ZN(SBOX_PL_3_n126) );
  NAND2_X1 SBOX_PL_3_U56 ( .A1(1'b1), .A2(SBOX_Zl_f3[6]), .ZN(SBOX_PL_3_n244)
         );
  OAI21_X1 SBOX_PL_3_U55 ( .B1(1'b1), .B2(SBOX_PL_3_n161), .A(SBOX_PL_3_n243), 
        .ZN(SBOX_PL_3_n125) );
  NAND2_X1 SBOX_PL_3_U54 ( .A1(1'b1), .A2(SBOX_Zl_f3[7]), .ZN(SBOX_PL_3_n243)
         );
  OAI21_X1 SBOX_PL_3_U53 ( .B1(1'b1), .B2(SBOX_PL_3_n160), .A(SBOX_PL_3_n242), 
        .ZN(SBOX_PL_3_n124) );
  NAND2_X1 SBOX_PL_3_U52 ( .A1(1'b1), .A2(SBOX_Zl_f3[8]), .ZN(SBOX_PL_3_n242)
         );
  OAI21_X1 SBOX_PL_3_U51 ( .B1(1'b1), .B2(SBOX_PL_3_n159), .A(SBOX_PL_3_n241), 
        .ZN(SBOX_PL_3_n123) );
  NAND2_X1 SBOX_PL_3_U50 ( .A1(1'b1), .A2(SBOX_Zl_f3[9]), .ZN(SBOX_PL_3_n241)
         );
  OAI21_X1 SBOX_PL_3_U49 ( .B1(1'b1), .B2(SBOX_PL_3_n158), .A(SBOX_PL_3_n240), 
        .ZN(SBOX_PL_3_n122) );
  NAND2_X1 SBOX_PL_3_U48 ( .A1(1'b1), .A2(SBOX_Zl_f3[10]), .ZN(SBOX_PL_3_n240)
         );
  OAI21_X1 SBOX_PL_3_U47 ( .B1(1'b1), .B2(SBOX_PL_3_n157), .A(SBOX_PL_3_n239), 
        .ZN(SBOX_PL_3_n121) );
  NAND2_X1 SBOX_PL_3_U46 ( .A1(1'b1), .A2(SBOX_Zl_f3[11]), .ZN(SBOX_PL_3_n239)
         );
  OAI21_X1 SBOX_PL_3_U45 ( .B1(1'b1), .B2(SBOX_PL_3_n156), .A(SBOX_PL_3_n238), 
        .ZN(SBOX_PL_3_n120) );
  NAND2_X1 SBOX_PL_3_U44 ( .A1(1'b1), .A2(SBOX_Zh_f3[0]), .ZN(SBOX_PL_3_n238)
         );
  OAI21_X1 SBOX_PL_3_U43 ( .B1(1'b1), .B2(SBOX_PL_3_n155), .A(SBOX_PL_3_n237), 
        .ZN(SBOX_PL_3_n119) );
  NAND2_X1 SBOX_PL_3_U42 ( .A1(1'b1), .A2(SBOX_Zh_f3[1]), .ZN(SBOX_PL_3_n237)
         );
  OAI21_X1 SBOX_PL_3_U41 ( .B1(1'b1), .B2(SBOX_PL_3_n154), .A(SBOX_PL_3_n236), 
        .ZN(SBOX_PL_3_n118) );
  NAND2_X1 SBOX_PL_3_U40 ( .A1(1'b1), .A2(SBOX_Zh_f3[2]), .ZN(SBOX_PL_3_n236)
         );
  OAI21_X1 SBOX_PL_3_U39 ( .B1(1'b1), .B2(SBOX_PL_3_n153), .A(SBOX_PL_3_n235), 
        .ZN(SBOX_PL_3_n117) );
  NAND2_X1 SBOX_PL_3_U38 ( .A1(1'b1), .A2(SBOX_Zh_f3[3]), .ZN(SBOX_PL_3_n235)
         );
  OAI21_X1 SBOX_PL_3_U37 ( .B1(1'b1), .B2(SBOX_PL_3_n152), .A(SBOX_PL_3_n234), 
        .ZN(SBOX_PL_3_n116) );
  NAND2_X1 SBOX_PL_3_U36 ( .A1(1'b1), .A2(SBOX_Zh_f3[4]), .ZN(SBOX_PL_3_n234)
         );
  OAI21_X1 SBOX_PL_3_U35 ( .B1(1'b1), .B2(SBOX_PL_3_n151), .A(SBOX_PL_3_n233), 
        .ZN(SBOX_PL_3_n115) );
  NAND2_X1 SBOX_PL_3_U34 ( .A1(1'b1), .A2(SBOX_Zh_f3[5]), .ZN(SBOX_PL_3_n233)
         );
  OAI21_X1 SBOX_PL_3_U33 ( .B1(1'b1), .B2(SBOX_PL_3_n150), .A(SBOX_PL_3_n232), 
        .ZN(SBOX_PL_3_n114) );
  NAND2_X1 SBOX_PL_3_U32 ( .A1(1'b1), .A2(SBOX_Zh_f3[6]), .ZN(SBOX_PL_3_n232)
         );
  OAI21_X1 SBOX_PL_3_U31 ( .B1(1'b1), .B2(SBOX_PL_3_n149), .A(SBOX_PL_3_n231), 
        .ZN(SBOX_PL_3_n113) );
  NAND2_X1 SBOX_PL_3_U30 ( .A1(1'b1), .A2(SBOX_Zh_f3[7]), .ZN(SBOX_PL_3_n231)
         );
  OAI21_X1 SBOX_PL_3_U29 ( .B1(1'b1), .B2(SBOX_PL_3_n148), .A(SBOX_PL_3_n230), 
        .ZN(SBOX_PL_3_n112) );
  NAND2_X1 SBOX_PL_3_U28 ( .A1(1'b1), .A2(SBOX_Zh_f3[8]), .ZN(SBOX_PL_3_n230)
         );
  OAI21_X1 SBOX_PL_3_U27 ( .B1(1'b1), .B2(SBOX_PL_3_n147), .A(SBOX_PL_3_n229), 
        .ZN(SBOX_PL_3_n111) );
  NAND2_X1 SBOX_PL_3_U26 ( .A1(1'b1), .A2(SBOX_Zh_f3[9]), .ZN(SBOX_PL_3_n229)
         );
  OAI21_X1 SBOX_PL_3_U25 ( .B1(1'b1), .B2(SBOX_PL_3_n146), .A(SBOX_PL_3_n228), 
        .ZN(SBOX_PL_3_n110) );
  NAND2_X1 SBOX_PL_3_U24 ( .A1(1'b1), .A2(SBOX_Zh_f3[10]), .ZN(SBOX_PL_3_n228)
         );
  OAI21_X1 SBOX_PL_3_U23 ( .B1(1'b1), .B2(SBOX_PL_3_n145), .A(SBOX_PL_3_n227), 
        .ZN(SBOX_PL_3_n109) );
  NAND2_X1 SBOX_PL_3_U22 ( .A1(1'b1), .A2(SBOX_Zh_f3[11]), .ZN(SBOX_PL_3_n227)
         );
  OAI21_X1 SBOX_PL_3_U21 ( .B1(1'b1), .B2(SBOX_PL_3_n177), .A(SBOX_PL_3_n226), 
        .ZN(SBOX_PL_3_n141) );
  NAND2_X1 SBOX_PL_3_U20 ( .A1(1'b1), .A2(SBOX_muld[3]), .ZN(SBOX_PL_3_n226)
         );
  OAI21_X1 SBOX_PL_3_U19 ( .B1(1'b1), .B2(SBOX_PL_3_n170), .A(SBOX_PL_3_n225), 
        .ZN(SBOX_PL_3_n134) );
  NAND2_X1 SBOX_PL_3_U18 ( .A1(1'b1), .A2(SBOX_muld[10]), .ZN(SBOX_PL_3_n225)
         );
  OAI21_X1 SBOX_PL_3_U17 ( .B1(1'b1), .B2(SBOX_PL_3_n169), .A(SBOX_PL_3_n224), 
        .ZN(SBOX_PL_3_n133) );
  NAND2_X1 SBOX_PL_3_U16 ( .A1(1'b1), .A2(SBOX_muld[11]), .ZN(SBOX_PL_3_n224)
         );
  OAI21_X1 SBOX_PL_3_U15 ( .B1(1'b1), .B2(SBOX_PL_3_n171), .A(SBOX_PL_3_n223), 
        .ZN(SBOX_PL_3_n135) );
  NAND2_X1 SBOX_PL_3_U14 ( .A1(1'b1), .A2(SBOX_muld[9]), .ZN(SBOX_PL_3_n223)
         );
  OAI21_X1 SBOX_PL_3_U13 ( .B1(1'b1), .B2(SBOX_PL_3_n172), .A(SBOX_PL_3_n222), 
        .ZN(SBOX_PL_3_n136) );
  NAND2_X1 SBOX_PL_3_U12 ( .A1(1'b1), .A2(SBOX_muld[8]), .ZN(SBOX_PL_3_n222)
         );
  OAI21_X1 SBOX_PL_3_U11 ( .B1(1'b1), .B2(SBOX_PL_3_n173), .A(SBOX_PL_3_n221), 
        .ZN(SBOX_PL_3_n137) );
  NAND2_X1 SBOX_PL_3_U10 ( .A1(1'b1), .A2(SBOX_muld[7]), .ZN(SBOX_PL_3_n221)
         );
  OAI21_X1 SBOX_PL_3_U9 ( .B1(1'b1), .B2(SBOX_PL_3_n175), .A(SBOX_PL_3_n220), 
        .ZN(SBOX_PL_3_n139) );
  NAND2_X1 SBOX_PL_3_U8 ( .A1(1'b1), .A2(SBOX_muld[5]), .ZN(SBOX_PL_3_n220) );
  OAI21_X1 SBOX_PL_3_U7 ( .B1(1'b1), .B2(SBOX_PL_3_n176), .A(SBOX_PL_3_n219), 
        .ZN(SBOX_PL_3_n140) );
  NAND2_X1 SBOX_PL_3_U6 ( .A1(1'b1), .A2(SBOX_muld[4]), .ZN(SBOX_PL_3_n219) );
  OAI21_X1 SBOX_PL_3_U5 ( .B1(1'b1), .B2(SBOX_PL_3_n178), .A(SBOX_PL_3_n218), 
        .ZN(SBOX_PL_3_n142) );
  NAND2_X1 SBOX_PL_3_U4 ( .A1(1'b1), .A2(SBOX_muld[2]), .ZN(SBOX_PL_3_n218) );
  OAI21_X1 SBOX_PL_3_U3 ( .B1(1'b1), .B2(SBOX_PL_3_n179), .A(SBOX_PL_3_n217), 
        .ZN(SBOX_PL_3_n143) );
  NAND2_X1 SBOX_PL_3_U2 ( .A1(1'b1), .A2(SBOX_muld[1]), .ZN(SBOX_PL_3_n217) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_0_ ( .D(SBOX_PL_3_n144), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[0]), .QN(SBOX_PL_3_n180) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_1_ ( .D(SBOX_PL_3_n143), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[1]), .QN(SBOX_PL_3_n179) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_2_ ( .D(SBOX_PL_3_n142), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[2]), .QN(SBOX_PL_3_n178) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_3_ ( .D(SBOX_PL_3_n141), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[3]), .QN(SBOX_PL_3_n177) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_4_ ( .D(SBOX_PL_3_n140), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[4]), .QN(SBOX_PL_3_n176) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_5_ ( .D(SBOX_PL_3_n139), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[5]), .QN(SBOX_PL_3_n175) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_6_ ( .D(SBOX_PL_3_n138), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[6]), .QN(SBOX_PL_3_n174) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_7_ ( .D(SBOX_PL_3_n137), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[7]), .QN(SBOX_PL_3_n173) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_8_ ( .D(SBOX_PL_3_n136), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[8]), .QN(SBOX_PL_3_n172) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_9_ ( .D(SBOX_PL_3_n135), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[9]), .QN(SBOX_PL_3_n171) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_10_ ( .D(SBOX_PL_3_n134), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[10]), .QN(SBOX_PL_3_n170) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_11_ ( .D(SBOX_PL_3_n133), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[11]), .QN(SBOX_PL_3_n169) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_12_ ( .D(SBOX_PL_3_n132), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[12]), .QN(SBOX_PL_3_n168) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_13_ ( .D(SBOX_PL_3_n131), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[13]), .QN(SBOX_PL_3_n167) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_14_ ( .D(SBOX_PL_3_n130), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[14]), .QN(SBOX_PL_3_n166) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_15_ ( .D(SBOX_PL_3_n129), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[15]), .QN(SBOX_PL_3_n165) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_16_ ( .D(SBOX_PL_3_n128), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[16]), .QN(SBOX_PL_3_n164) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_17_ ( .D(SBOX_PL_3_n127), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[17]), .QN(SBOX_PL_3_n163) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_18_ ( .D(SBOX_PL_3_n126), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[18]), .QN(SBOX_PL_3_n162) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_19_ ( .D(SBOX_PL_3_n125), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[19]), .QN(SBOX_PL_3_n161) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_20_ ( .D(SBOX_PL_3_n124), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[20]), .QN(SBOX_PL_3_n160) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_21_ ( .D(SBOX_PL_3_n123), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[21]), .QN(SBOX_PL_3_n159) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_22_ ( .D(SBOX_PL_3_n122), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[22]), .QN(SBOX_PL_3_n158) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_23_ ( .D(SBOX_PL_3_n121), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[23]), .QN(SBOX_PL_3_n157) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_24_ ( .D(SBOX_PL_3_n120), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[24]), .QN(SBOX_PL_3_n156) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_25_ ( .D(SBOX_PL_3_n119), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[25]), .QN(SBOX_PL_3_n155) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_26_ ( .D(SBOX_PL_3_n118), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[26]), .QN(SBOX_PL_3_n154) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_27_ ( .D(SBOX_PL_3_n117), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[27]), .QN(SBOX_PL_3_n153) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_28_ ( .D(SBOX_PL_3_n116), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[28]), .QN(SBOX_PL_3_n152) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_29_ ( .D(SBOX_PL_3_n115), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[29]), .QN(SBOX_PL_3_n151) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_30_ ( .D(SBOX_PL_3_n114), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[30]), .QN(SBOX_PL_3_n150) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_31_ ( .D(SBOX_PL_3_n113), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[31]), .QN(SBOX_PL_3_n149) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_32_ ( .D(SBOX_PL_3_n112), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[32]), .QN(SBOX_PL_3_n148) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_33_ ( .D(SBOX_PL_3_n111), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[33]), .QN(SBOX_PL_3_n147) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_34_ ( .D(SBOX_PL_3_n110), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[34]), .QN(SBOX_PL_3_n146) );
  DFF_X1 SBOX_PL_3_s_current_state_reg_35_ ( .D(SBOX_PL_3_n109), .CK(ClkxCI), 
        .Q(SBOX_FF3_out[35]), .QN(SBOX_PL_3_n145) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U12 ( .A(SBOX_FF3_out[11]), .B(SBOX_FF3_out[9]), 
        .Z(SBOX_Inst_f4_multd_L_sB[5]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U11 ( .A(SBOX_FF3_out[10]), .B(SBOX_FF3_out[8]), 
        .Z(SBOX_Inst_f4_multd_L_sB[4]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U10 ( .A(SBOX_FF3_out[4]), .B(SBOX_FF3_out[6]), 
        .Z(SBOX_Inst_f4_multd_L_sB[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U9 ( .A(SBOX_FF3_out[1]), .B(SBOX_FF3_out[3]), 
        .Z(SBOX_Inst_f4_multd_L_sB[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U8 ( .A(SBOX_FF3_out[0]), .B(SBOX_FF3_out[2]), 
        .Z(SBOX_Inst_f4_multd_L_sB[0]) );
  XOR2_X2 SBOX_Inst_f4_multd_L_U7 ( .A(SBOX_FF3_out[34]), .B(SBOX_FF3_out[32]), 
        .Z(SBOX_Inst_f4_multd_L_sA[4]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U6 ( .A(SBOX_FF3_out[28]), .B(SBOX_FF3_out[30]), 
        .Z(SBOX_Inst_f4_multd_L_sA[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U5 ( .A(SBOX_FF3_out[5]), .B(SBOX_FF3_out[7]), 
        .Z(SBOX_Inst_f4_multd_L_sB[3]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U4 ( .A(SBOX_FF3_out[25]), .B(SBOX_FF3_out[27]), 
        .Z(SBOX_Inst_f4_multd_L_sA[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U3 ( .A(SBOX_FF3_out[24]), .B(SBOX_FF3_out[26]), 
        .Z(SBOX_Inst_f4_multd_L_sA[0]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U2 ( .A(SBOX_FF3_out[29]), .B(SBOX_FF3_out[31]), 
        .Z(SBOX_Inst_f4_multd_L_sA[3]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_U1 ( .A(SBOX_FF3_out[35]), .B(SBOX_FF3_out[33]), 
        .Z(SBOX_Inst_f4_multd_L_sA[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U93 ( .A(SBOX_Inst_f4_multd_L_himul_n294), .B(SBOX_Inst_f4_multd_L_himul_n293), .ZN(SBOX_Inst_f4_multd_L_himul_n302) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U92 ( .A(SBOX_Inst_f4_multd_L_himul_n292), .B(SBOX_Inst_f4_multd_L_himul_n291), .ZN(SBOX_Inst_f4_multd_L_himul_n293) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U91 ( .A1(SBOX_FF3_out[30]), .A2(
        SBOX_FF3_out[3]), .ZN(SBOX_Inst_f4_multd_L_himul_n291) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U90 ( .A1(SBOX_FF3_out[6]), .A2(
        SBOX_FF3_out[27]), .ZN(SBOX_Inst_f4_multd_L_himul_n292) );
  AOI221_X1 SBOX_Inst_f4_multd_L_himul_U89 ( .B1(SBOX_FF3_out[3]), .B2(
        SBOX_FF3_out[7]), .C1(SBOX_Inst_f4_multd_L_himul_n290), .C2(
        SBOX_Inst_f4_multd_L_himul_n289), .A(SBOX_Inst_f4_multd_L_himul_n299), 
        .ZN(SBOX_Inst_f4_multd_L_himul_n294) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U88 ( .A(SBOX_Inst_f4_multd_L_himul_n285), 
        .B(SBOX_Inst_f4_multd_L_himul_n284), .Z(
        SBOX_Inst_f4_multd_L_himul_n295) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U87 ( .A1(SBOX_FF3_out[3]), .A2(
        SBOX_FF3_out[26]), .ZN(SBOX_Inst_f4_multd_L_himul_n284) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U86 ( .A1(SBOX_FF3_out[2]), .A2(
        SBOX_FF3_out[27]), .ZN(SBOX_Inst_f4_multd_L_himul_n285) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U85 ( .A(SBOX_Inst_f4_multd_L_himul_n283), 
        .B(SBOX_Inst_f4_multd_L_himul_n282), .Z(
        SBOX_Inst_f4_multd_L_himul_n286) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U84 ( .A1(SBOX_FF3_out[2]), .A2(
        SBOX_FF3_out[35]), .ZN(SBOX_Inst_f4_multd_L_himul_n282) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U83 ( .A1(SBOX_FF3_out[34]), .A2(
        SBOX_FF3_out[3]), .ZN(SBOX_Inst_f4_multd_L_himul_n283) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U82 ( .A(SBOX_FF3_out[3]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n290) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U81 ( .A(SBOX_Inst_f4_multd_L_himul_n281), .B(SBOX_Inst_f4_multd_L_himul_n280), .ZN(SBOX_Inst_f4_multd_L_Orig_ph[1]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U80 ( .A(SBOX_Inst_f4_multd_L_himul_n279), .B(SBOX_Inst_f4_multd_L_himul_n278), .ZN(SBOX_Inst_f4_multd_L_himul_n280) );
  OAI221_X1 SBOX_Inst_f4_multd_L_himul_U79 ( .B1(SBOX_FF3_out[7]), .B2(
        SBOX_FF3_out[6]), .C1(SBOX_Inst_f4_multd_L_himul_n289), .C2(
        SBOX_Inst_f4_multd_L_himul_n277), .A(SBOX_FF3_out[31]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n278) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U78 ( .A(SBOX_Inst_f4_multd_L_himul_n276), .B(SBOX_Inst_f4_multd_L_himul_n275), .ZN(SBOX_Inst_f4_multd_L_himul_n279) );
  OAI221_X1 SBOX_Inst_f4_multd_L_himul_U77 ( .B1(SBOX_FF3_out[30]), .B2(
        SBOX_FF3_out[31]), .C1(SBOX_Inst_f4_multd_L_himul_n300), .C2(
        SBOX_Inst_f4_multd_L_himul_n298), .A(SBOX_FF3_out[10]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n275) );
  AOI22_X1 SBOX_Inst_f4_multd_L_himul_U76 ( .A1(SBOX_FF3_out[7]), .A2(
        SBOX_FF3_out[6]), .B1(SBOX_Inst_f4_multd_L_himul_n277), .B2(
        SBOX_Inst_f4_multd_L_himul_n289), .ZN(SBOX_Inst_f4_multd_L_himul_n296)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U75 ( .A(SBOX_Inst_f4_multd_L_himul_n273), .B(SBOX_Inst_f4_multd_L_himul_n272), .ZN(SBOX_Inst_f4_multd_L_himul_n281) );
  AOI221_X1 SBOX_Inst_f4_multd_L_himul_U74 ( .B1(SBOX_FF3_out[35]), .B2(
        SBOX_FF3_out[30]), .C1(SBOX_FF3_out[6]), .C2(SBOX_FF3_out[11]), .A(
        SBOX_Inst_f4_multd_L_himul_n267), .ZN(SBOX_Inst_f4_multd_L_himul_n273)
         );
  OAI22_X1 SBOX_Inst_f4_multd_L_himul_U73 ( .A1(SBOX_FF3_out[35]), .A2(
        SBOX_FF3_out[30]), .B1(SBOX_FF3_out[11]), .B2(SBOX_FF3_out[6]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n267) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U72 ( .A(SBOX_Inst_f4_multd_L_himul_n266), .B(SBOX_Inst_f4_multd_L_himul_n265), .ZN(SBOX_Inst_f4_multd_L_Orig_ph[0]) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U71 ( .A1(SBOX_FF3_out[7]), .A2(
        SBOX_Inst_f4_multd_L_himul_n269), .ZN(SBOX_Inst_f4_multd_L_himul_n265)
         );
  OAI21_X1 SBOX_Inst_f4_multd_L_himul_U70 ( .B1(SBOX_FF3_out[34]), .B2(
        SBOX_Inst_f4_multd_L_himul_n287), .A(SBOX_Inst_f4_multd_L_himul_n270), 
        .ZN(SBOX_Inst_f4_multd_L_himul_n269) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U69 ( .A(SBOX_Inst_f4_multd_L_himul_n264), 
        .B(SBOX_Inst_f4_multd_L_himul_n263), .Z(
        SBOX_Inst_f4_multd_L_himul_n266) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U68 ( .A(SBOX_Inst_f4_multd_L_himul_n262), .B(SBOX_Inst_f4_multd_L_himul_n261), .ZN(SBOX_Inst_f4_multd_L_himul_n263) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U67 ( .A1(SBOX_FF3_out[31]), .A2(
        SBOX_FF3_out[11]), .ZN(SBOX_Inst_f4_multd_L_himul_n261) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U66 ( .A(SBOX_Inst_f4_multd_L_himul_n259), .B(SBOX_Inst_f4_multd_L_himul_n258), .ZN(SBOX_Inst_f4_multd_L_himul_n260) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U65 ( .A1(
        SBOX_Inst_f4_multd_L_himul_n298), .A2(SBOX_FF3_out[10]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n259) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U64 ( .A(SBOX_FF3_out[6]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n277) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U63 ( .A(SBOX_Inst_f4_multd_L_himul_n256), .B(SBOX_Inst_f4_multd_L_himul_n257), .ZN(SBOX_Inst_f4_multd_L_himul_n301) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U62 ( .A1(SBOX_FF3_out[30]), .A2(
        SBOX_FF3_out[6]), .ZN(SBOX_Inst_f4_multd_L_himul_n257) );
  NOR2_X1 SBOX_Inst_f4_multd_L_himul_U61 ( .A1(SBOX_Inst_f4_multd_L_himul_n289), .A2(SBOX_Inst_f4_multd_L_himul_n298), .ZN(SBOX_Inst_f4_multd_L_himul_n256)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U60 ( .A(SBOX_Inst_f4_multd_L_himul_n302), .B(SBOX_Inst_f4_multd_L_himul_n255), .ZN(SBOX_Inst_f4_multd_L_Orig_ph[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U59 ( .A(SBOX_Inst_f4_multd_L_himul_n248), .B(SBOX_Inst_f4_multd_L_himul_n254), .ZN(SBOX_Inst_f4_multd_L_himul_n255) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U58 ( .A(SBOX_Inst_f4_multd_L_himul_n253), .B(SBOX_Inst_f4_multd_L_himul_n252), .ZN(SBOX_Inst_f4_multd_L_himul_n254) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U57 ( .A(SBOX_Inst_f4_multd_L_himul_n251), .B(SBOX_Inst_f4_multd_L_himul_n301), .ZN(SBOX_Inst_f4_multd_L_himul_n253) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U56 ( .A1(SBOX_FF3_out[2]), .A2(
        SBOX_FF3_out[31]), .ZN(SBOX_Inst_f4_multd_L_himul_n252) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U55 ( .A(SBOX_Inst_f4_multd_L_himul_n249), 
        .B(SBOX_Inst_f4_multd_L_himul_n250), .Z(
        SBOX_Inst_f4_multd_L_himul_n251) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U54 ( .A1(SBOX_FF3_out[6]), .A2(
        SBOX_FF3_out[26]), .ZN(SBOX_Inst_f4_multd_L_himul_n250) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U53 ( .A1(SBOX_FF3_out[3]), .A2(
        SBOX_FF3_out[27]), .ZN(SBOX_Inst_f4_multd_L_himul_n249) );
  AOI22_X1 SBOX_Inst_f4_multd_L_himul_U52 ( .A1(SBOX_FF3_out[2]), .A2(
        SBOX_Inst_f4_multd_L_himul_n246), .B1(SBOX_FF3_out[27]), .B2(
        SBOX_Inst_f4_multd_L_himul_n247), .ZN(SBOX_Inst_f4_multd_L_himul_n248)
         );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U51 ( .A(SBOX_FF3_out[2]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n247) );
  OAI22_X1 SBOX_Inst_f4_multd_L_himul_U50 ( .A1(SBOX_FF3_out[26]), .A2(
        SBOX_Inst_f4_multd_L_himul_n300), .B1(SBOX_FF3_out[30]), .B2(
        SBOX_Inst_f4_multd_L_himul_n299), .ZN(SBOX_Inst_f4_multd_L_himul_n246)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U49 ( .A(SBOX_Inst_f4_multd_L_himul_n245), .B(SBOX_Inst_f4_multd_L_himul_n244), .ZN(SBOX_Inst_f4_multd_L_Orig_ph[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U48 ( .A(SBOX_Inst_f4_multd_L_himul_n295), .B(SBOX_Inst_f4_multd_L_himul_n241), .ZN(SBOX_Inst_f4_multd_L_himul_n245) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U47 ( .A(SBOX_Inst_f4_multd_L_himul_n242), 
        .B(SBOX_Inst_f4_multd_L_himul_n243), .Z(
        SBOX_Inst_f4_multd_L_himul_n244) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U46 ( .A1(
        SBOX_Inst_f4_multd_L_himul_n296), .A2(SBOX_FF3_out[30]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n243) );
  NOR2_X1 SBOX_Inst_f4_multd_L_himul_U45 ( .A1(SBOX_FF3_out[7]), .A2(
        SBOX_Inst_f4_multd_L_himul_n297), .ZN(SBOX_Inst_f4_multd_L_himul_n242)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U44 ( .A(SBOX_Inst_f4_multd_L_himul_n302), .B(SBOX_Inst_f4_multd_L_himul_n240), .ZN(SBOX_Inst_f4_multd_L_himul_n241) );
  MUX2_X1 SBOX_Inst_f4_multd_L_himul_U43 ( .A(SBOX_FF3_out[2]), .B(
        SBOX_FF3_out[3]), .S(SBOX_Inst_f4_multd_L_himul_n239), .Z(
        SBOX_Inst_f4_multd_L_himul_n240) );
  AOI22_X1 SBOX_Inst_f4_multd_L_himul_U42 ( .A1(SBOX_FF3_out[31]), .A2(
        SBOX_FF3_out[27]), .B1(SBOX_Inst_f4_multd_L_himul_n297), .B2(
        SBOX_Inst_f4_multd_L_himul_n298), .ZN(SBOX_Inst_f4_multd_L_himul_n239)
         );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U41 ( .A(SBOX_Inst_f4_multd_L_himul_n237), 
        .B(SBOX_Inst_f4_multd_L_himul_n238), .Z(
        SBOX_Inst_f4_multd_L_Orig_ph[3]) );
  OAI221_X1 SBOX_Inst_f4_multd_L_himul_U40 ( .B1(
        SBOX_Inst_f4_multd_L_himul_n228), .B2(SBOX_FF3_out[27]), .C1(
        SBOX_Inst_f4_multd_L_himul_n227), .C2(SBOX_Inst_f4_multd_L_himul_n297), 
        .A(SBOX_FF3_out[10]), .ZN(SBOX_Inst_f4_multd_L_himul_n238) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U39 ( .A(SBOX_Inst_f4_multd_L_himul_n235), .B(SBOX_Inst_f4_multd_L_himul_n236), .ZN(SBOX_Inst_f4_multd_L_himul_n237) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U38 ( .A1(
        SBOX_Inst_f4_multd_L_himul_n288), .A2(SBOX_FF3_out[34]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n236) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U37 ( .A(SBOX_Inst_f4_multd_L_himul_n234), 
        .B(SBOX_Inst_f4_multd_L_himul_n287), .Z(
        SBOX_Inst_f4_multd_L_himul_n235) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U36 ( .A(SBOX_Inst_f4_multd_L_himul_n232), .B(SBOX_Inst_f4_multd_L_himul_n233), .ZN(SBOX_Inst_f4_multd_L_himul_n234) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U35 ( .A1(
        SBOX_Inst_f4_multd_L_himul_n228), .A2(SBOX_FF3_out[11]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n233) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U34 ( .A(SBOX_Inst_f4_multd_L_himul_n231), 
        .B(SBOX_Inst_f4_multd_L_himul_n286), .Z(
        SBOX_Inst_f4_multd_L_himul_n232) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U33 ( .A(SBOX_Inst_f4_multd_L_himul_n229), 
        .B(SBOX_Inst_f4_multd_L_himul_n230), .Z(
        SBOX_Inst_f4_multd_L_himul_n231) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U32 ( .A1(
        SBOX_Inst_f4_multd_L_himul_n290), .A2(SBOX_FF3_out[27]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n230) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U31 ( .A1(SBOX_FF3_out[34]), .A2(
        SBOX_FF3_out[2]), .ZN(SBOX_Inst_f4_multd_L_himul_n229) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U30 ( .A(SBOX_Inst_f4_multd_L_himul_n227), 
        .ZN(SBOX_Inst_f4_multd_L_himul_n228) );
  OAI22_X1 SBOX_Inst_f4_multd_L_himul_U29 ( .A1(SBOX_FF3_out[26]), .A2(
        SBOX_FF3_out[35]), .B1(SBOX_Inst_f4_multd_L_himul_n287), .B2(
        SBOX_Inst_f4_multd_L_himul_n299), .ZN(SBOX_Inst_f4_multd_L_himul_n227)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U28 ( .A(SBOX_Inst_f4_multd_L_himul_n225), .B(SBOX_Inst_f4_multd_L_himul_n226), .ZN(SBOX_Inst_f4_multd_L_Orig_ph[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U27 ( .A(SBOX_Inst_f4_multd_L_himul_n220), 
        .B(SBOX_Inst_f4_multd_L_himul_n286), .Z(
        SBOX_Inst_f4_multd_L_himul_n226) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U26 ( .A(SBOX_Inst_f4_multd_L_himul_n223), .B(SBOX_Inst_f4_multd_L_himul_n224), .ZN(SBOX_Inst_f4_multd_L_himul_n225) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U25 ( .A1(SBOX_FF3_out[26]), .A2(
        SBOX_FF3_out[11]), .ZN(SBOX_Inst_f4_multd_L_himul_n224) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U24 ( .A(SBOX_Inst_f4_multd_L_himul_n222), 
        .B(SBOX_Inst_f4_multd_L_himul_n295), .Z(
        SBOX_Inst_f4_multd_L_himul_n223) );
  AOI22_X1 SBOX_Inst_f4_multd_L_himul_U23 ( .A1(SBOX_FF3_out[2]), .A2(
        SBOX_FF3_out[27]), .B1(SBOX_Inst_f4_multd_L_himul_n297), .B2(
        SBOX_Inst_f4_multd_L_himul_n221), .ZN(SBOX_Inst_f4_multd_L_himul_n222)
         );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U22 ( .A(SBOX_FF3_out[2]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n221) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_himul_U21 ( .A(SBOX_Inst_f4_multd_L_himul_n217), .B(SBOX_Inst_f4_multd_L_himul_n219), .ZN(SBOX_Inst_f4_multd_L_himul_n220) );
  OAI211_X1 SBOX_Inst_f4_multd_L_himul_U20 ( .C1(
        SBOX_Inst_f4_multd_L_himul_n216), .C2(SBOX_FF3_out[10]), .A(
        SBOX_FF3_out[35]), .B(SBOX_Inst_f4_multd_L_himul_n218), .ZN(
        SBOX_Inst_f4_multd_L_himul_n219) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U19 ( .A1(
        SBOX_Inst_f4_multd_L_himul_n216), .A2(SBOX_FF3_out[10]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n218) );
  AOI22_X1 SBOX_Inst_f4_multd_L_himul_U18 ( .A1(SBOX_FF3_out[11]), .A2(
        SBOX_FF3_out[27]), .B1(SBOX_FF3_out[10]), .B2(
        SBOX_Inst_f4_multd_L_himul_n297), .ZN(SBOX_Inst_f4_multd_L_himul_n217)
         );
  AOI22_X1 SBOX_Inst_f4_multd_L_himul_U17 ( .A1(SBOX_FF3_out[3]), .A2(
        SBOX_FF3_out[11]), .B1(SBOX_Inst_f4_multd_L_himul_n290), .B2(
        SBOX_Inst_f4_multd_L_himul_n288), .ZN(SBOX_Inst_f4_multd_L_himul_n216)
         );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U16 ( .A1(SBOX_FF3_out[34]), .A2(
        SBOX_FF3_out[10]), .ZN(SBOX_Inst_f4_multd_L_himul_n268) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U15 ( .A(SBOX_Inst_f4_multd_L_himul_n268), 
        .ZN(SBOX_Inst_f4_multd_L_himul_n271) );
  OAI221_X1 SBOX_Inst_f4_multd_L_himul_U14 ( .B1(SBOX_FF3_out[34]), .B2(
        SBOX_FF3_out[30]), .C1(SBOX_Inst_f4_multd_L_himul_n274), .C2(
        SBOX_Inst_f4_multd_L_himul_n300), .A(SBOX_Inst_f4_multd_L_himul_n296), 
        .ZN(SBOX_Inst_f4_multd_L_himul_n276) );
  AOI22_X1 SBOX_Inst_f4_multd_L_himul_U13 ( .A1(
        SBOX_Inst_f4_multd_L_himul_n271), .A2(SBOX_Inst_f4_multd_L_himul_n270), 
        .B1(SBOX_Inst_f4_multd_L_himul_n269), .B2(
        SBOX_Inst_f4_multd_L_himul_n268), .ZN(SBOX_Inst_f4_multd_L_himul_n272)
         );
  AOI221_X1 SBOX_Inst_f4_multd_L_himul_U12 ( .B1(SBOX_FF3_out[34]), .B2(
        SBOX_FF3_out[30]), .C1(SBOX_Inst_f4_multd_L_himul_n274), .C2(
        SBOX_Inst_f4_multd_L_himul_n300), .A(SBOX_Inst_f4_multd_L_himul_n288), 
        .ZN(SBOX_Inst_f4_multd_L_himul_n258) );
  XOR2_X1 SBOX_Inst_f4_multd_L_himul_U11 ( .A(SBOX_Inst_f4_multd_L_himul_n301), 
        .B(SBOX_Inst_f4_multd_L_himul_n260), .Z(
        SBOX_Inst_f4_multd_L_himul_n262) );
  AOI221_X1 SBOX_Inst_f4_multd_L_himul_U10 ( .B1(SBOX_FF3_out[35]), .B2(
        SBOX_FF3_out[31]), .C1(SBOX_Inst_f4_multd_L_himul_n287), .C2(
        SBOX_Inst_f4_multd_L_himul_n298), .A(SBOX_Inst_f4_multd_L_himul_n277), 
        .ZN(SBOX_Inst_f4_multd_L_himul_n264) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U9 ( .A(SBOX_FF3_out[30]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n300) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U8 ( .A(SBOX_FF3_out[26]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n299) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U7 ( .A(SBOX_FF3_out[27]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n297) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U6 ( .A(SBOX_FF3_out[31]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n298) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U5 ( .A(SBOX_FF3_out[35]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n287) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U4 ( .A(SBOX_FF3_out[11]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n288) );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U3 ( .A(SBOX_FF3_out[7]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n289) );
  NAND2_X1 SBOX_Inst_f4_multd_L_himul_U2 ( .A1(SBOX_FF3_out[34]), .A2(
        SBOX_Inst_f4_multd_L_himul_n287), .ZN(SBOX_Inst_f4_multd_L_himul_n270)
         );
  INV_X1 SBOX_Inst_f4_multd_L_himul_U1 ( .A(SBOX_FF3_out[34]), .ZN(
        SBOX_Inst_f4_multd_L_himul_n274) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U8 ( .A(PRNGQ[41]), .B(
        SBOX_Inst_f4_multd_L_Orig_ph[1]), .Z(SBOX_ph_L[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U7 ( .A(PRNGQ[40]), .B(
        SBOX_Inst_f4_multd_L_Orig_ph[0]), .Z(SBOX_ph_L[0]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U6 ( .A(
        SBOX_Inst_f4_multd_L_AddNewMaskph_n6), .B(PRNGQ[43]), .ZN(SBOX_ph_L[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U5 ( .A(PRNGQ[41]), .B(
        SBOX_Inst_f4_multd_L_Orig_ph[5]), .ZN(
        SBOX_Inst_f4_multd_L_AddNewMaskph_n6) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U4 ( .A(
        SBOX_Inst_f4_multd_L_AddNewMaskph_n5), .B(PRNGQ[42]), .ZN(SBOX_ph_L[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U3 ( .A(PRNGQ[40]), .B(
        SBOX_Inst_f4_multd_L_Orig_ph[4]), .ZN(
        SBOX_Inst_f4_multd_L_AddNewMaskph_n5) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U2 ( .A(PRNGQ[43]), .B(
        SBOX_Inst_f4_multd_L_Orig_ph[3]), .Z(SBOX_ph_L[3]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskph_U1 ( .A(PRNGQ[42]), .B(
        SBOX_Inst_f4_multd_L_Orig_ph[2]), .Z(SBOX_ph_L[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U90 ( .A(
        SBOX_Inst_f4_multd_L_summul_n298), .B(SBOX_Inst_f4_multd_L_summul_n297), .ZN(SBOX_Inst_f4_multd_L_Orig_p[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U89 ( .A(
        SBOX_Inst_f4_multd_L_summul_n296), .B(SBOX_Inst_f4_multd_L_summul_n295), .ZN(SBOX_Inst_f4_multd_L_summul_n297) );
  XOR2_X1 SBOX_Inst_f4_multd_L_summul_U88 ( .A(
        SBOX_Inst_f4_multd_L_summul_n294), .B(SBOX_Inst_f4_multd_L_summul_n293), .Z(SBOX_Inst_f4_multd_L_summul_n295) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U87 ( .A1(SBOX_Inst_f4_multd_L_sB[0]), 
        .A2(SBOX_Inst_f4_multd_L_summul_n289), .B1(SBOX_Inst_f4_multd_L_sA[1]), 
        .B2(SBOX_Inst_f4_multd_L_summul_n288), .ZN(
        SBOX_Inst_f4_multd_L_summul_n294) );
  AOI221_X1 SBOX_Inst_f4_multd_L_summul_U86 ( .B1(SBOX_Inst_f4_multd_L_sB[3]), 
        .B2(SBOX_Inst_f4_multd_L_sB[0]), .C1(SBOX_Inst_f4_multd_L_summul_n283), 
        .C2(SBOX_Inst_f4_multd_L_summul_n288), .A(
        SBOX_Inst_f4_multd_L_summul_n282), .ZN(
        SBOX_Inst_f4_multd_L_summul_n284) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U85 ( .A(
        SBOX_Inst_f4_multd_L_summul_n281), .B(SBOX_Inst_f4_multd_L_summul_n280), .ZN(SBOX_Inst_f4_multd_L_Orig_p[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U84 ( .A(
        SBOX_Inst_f4_multd_L_summul_n279), .B(SBOX_Inst_f4_multd_L_summul_n278), .ZN(SBOX_Inst_f4_multd_L_summul_n280) );
  MUX2_X1 SBOX_Inst_f4_multd_L_summul_U83 ( .A(SBOX_Inst_f4_multd_L_sB[0]), 
        .B(SBOX_Inst_f4_multd_L_sB[1]), .S(SBOX_Inst_f4_multd_L_summul_n277), 
        .Z(SBOX_Inst_f4_multd_L_summul_n278) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U82 ( .A(
        SBOX_Inst_f4_multd_L_summul_n276), .B(SBOX_Inst_f4_multd_L_summul_n275), .ZN(SBOX_Inst_f4_multd_L_summul_n279) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U81 ( .A(
        SBOX_Inst_f4_multd_L_summul_n272), .B(SBOX_Inst_f4_multd_L_summul_n271), .ZN(SBOX_Inst_f4_multd_L_summul_n285) );
  XOR2_X1 SBOX_Inst_f4_multd_L_summul_U80 ( .A(
        SBOX_Inst_f4_multd_L_summul_n270), .B(SBOX_Inst_f4_multd_L_summul_n269), .Z(SBOX_Inst_f4_multd_L_summul_n271) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U79 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n289), .A2(SBOX_Inst_f4_multd_L_sB[1]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n272) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U78 ( .A(
        SBOX_Inst_f4_multd_L_summul_n264), .B(SBOX_Inst_f4_multd_L_summul_n263), .ZN(SBOX_Inst_f4_multd_L_Orig_p[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U77 ( .A(
        SBOX_Inst_f4_multd_L_summul_n262), .B(SBOX_Inst_f4_multd_L_summul_n261), .ZN(SBOX_Inst_f4_multd_L_summul_n263) );
  XOR2_X1 SBOX_Inst_f4_multd_L_summul_U76 ( .A(
        SBOX_Inst_f4_multd_L_summul_n260), .B(SBOX_Inst_f4_multd_L_summul_n259), .Z(SBOX_Inst_f4_multd_L_summul_n262) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U75 ( .A(
        SBOX_Inst_f4_multd_L_summul_n258), .B(SBOX_Inst_f4_multd_L_summul_n257), .ZN(SBOX_Inst_f4_multd_L_summul_n259) );
  MUX2_X1 SBOX_Inst_f4_multd_L_summul_U74 ( .A(SBOX_Inst_f4_multd_L_sB[4]), 
        .B(SBOX_Inst_f4_multd_L_summul_n256), .S(SBOX_Inst_f4_multd_L_sA[5]), 
        .Z(SBOX_Inst_f4_multd_L_summul_n257) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U73 ( .A1(SBOX_Inst_f4_multd_L_sB[5]), 
        .A2(SBOX_Inst_f4_multd_L_sB[1]), .B1(SBOX_Inst_f4_multd_L_summul_n287), 
        .B2(SBOX_Inst_f4_multd_L_summul_n255), .ZN(
        SBOX_Inst_f4_multd_L_summul_n256) );
  OAI221_X1 SBOX_Inst_f4_multd_L_summul_U72 ( .B1(SBOX_Inst_f4_multd_L_sB[5]), 
        .B2(SBOX_Inst_f4_multd_L_sB[4]), .C1(SBOX_Inst_f4_multd_L_summul_n255), 
        .C2(SBOX_Inst_f4_multd_L_summul_n254), .A(SBOX_Inst_f4_multd_L_sA[1]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n258) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U71 ( .A1(SBOX_Inst_f4_multd_L_sA[1]), 
        .A2(SBOX_Inst_f4_multd_L_sB[0]), .B1(SBOX_Inst_f4_multd_L_summul_n288), 
        .B2(SBOX_Inst_f4_multd_L_summul_n286), .ZN(
        SBOX_Inst_f4_multd_L_summul_n260) );
  XOR2_X1 SBOX_Inst_f4_multd_L_summul_U70 ( .A(
        SBOX_Inst_f4_multd_L_summul_n253), .B(SBOX_Inst_f4_multd_L_summul_n252), .Z(SBOX_Inst_f4_multd_L_summul_n265) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U69 ( .A1(SBOX_Inst_f4_multd_L_sB[1]), 
        .A2(SBOX_Inst_f4_multd_L_sA[4]), .ZN(SBOX_Inst_f4_multd_L_summul_n252)
         );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U68 ( .A1(SBOX_Inst_f4_multd_L_sB[0]), 
        .A2(SBOX_Inst_f4_multd_L_sA[5]), .ZN(SBOX_Inst_f4_multd_L_summul_n253)
         );
  XOR2_X1 SBOX_Inst_f4_multd_L_summul_U67 ( .A(
        SBOX_Inst_f4_multd_L_summul_n251), .B(SBOX_Inst_f4_multd_L_summul_n250), .Z(SBOX_Inst_f4_multd_L_summul_n273) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U66 ( .A1(SBOX_Inst_f4_multd_L_sA[1]), 
        .A2(SBOX_Inst_f4_multd_L_sB[0]), .ZN(SBOX_Inst_f4_multd_L_summul_n251)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U65 ( .A(
        SBOX_Inst_f4_multd_L_summul_n249), .B(SBOX_Inst_f4_multd_L_summul_n248), .ZN(SBOX_Inst_f4_multd_L_Orig_p[1]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U64 ( .A(
        SBOX_Inst_f4_multd_L_summul_n247), .B(SBOX_Inst_f4_multd_L_summul_n246), .ZN(SBOX_Inst_f4_multd_L_summul_n248) );
  OAI221_X1 SBOX_Inst_f4_multd_L_summul_U63 ( .B1(SBOX_Inst_f4_multd_L_sA[4]), 
        .B2(SBOX_Inst_f4_multd_L_sA[3]), .C1(SBOX_Inst_f4_multd_L_summul_n245), 
        .C2(SBOX_Inst_f4_multd_L_summul_n282), .A(SBOX_Inst_f4_multd_L_sB[4]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n246) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U62 ( .A(
        SBOX_Inst_f4_multd_L_summul_n244), .B(SBOX_Inst_f4_multd_L_summul_n243), .ZN(SBOX_Inst_f4_multd_L_summul_n247) );
  OAI221_X1 SBOX_Inst_f4_multd_L_summul_U61 ( .B1(SBOX_Inst_f4_multd_L_sB[3]), 
        .B2(SBOX_Inst_f4_multd_L_sB[2]), .C1(SBOX_Inst_f4_multd_L_summul_n283), 
        .C2(SBOX_Inst_f4_multd_L_summul_n290), .A(SBOX_Inst_f4_multd_L_sA[3]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n243) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U60 ( .A(
        SBOX_Inst_f4_multd_L_summul_n242), .B(SBOX_Inst_f4_multd_L_sA[4]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n244) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U59 ( .A(
        SBOX_Inst_f4_multd_L_summul_n241), .B(SBOX_Inst_f4_multd_L_summul_n240), .ZN(SBOX_Inst_f4_multd_L_summul_n242) );
  OAI221_X1 SBOX_Inst_f4_multd_L_summul_U58 ( .B1(SBOX_Inst_f4_multd_L_sB[4]), 
        .B2(SBOX_Inst_f4_multd_L_summul_n239), .C1(
        SBOX_Inst_f4_multd_L_summul_n254), .C2(
        SBOX_Inst_f4_multd_L_summul_n238), .A(SBOX_Inst_f4_multd_L_sA[2]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n240) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U57 ( .A1(SBOX_Inst_f4_multd_L_sB[5]), 
        .A2(SBOX_Inst_f4_multd_L_sB[2]), .B1(SBOX_Inst_f4_multd_L_summul_n290), 
        .B2(SBOX_Inst_f4_multd_L_summul_n255), .ZN(
        SBOX_Inst_f4_multd_L_summul_n239) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U56 ( .A1(SBOX_Inst_f4_multd_L_sB[3]), 
        .A2(SBOX_Inst_f4_multd_L_summul_n290), .B1(SBOX_Inst_f4_multd_L_sB[2]), 
        .B2(SBOX_Inst_f4_multd_L_summul_n283), .ZN(
        SBOX_Inst_f4_multd_L_summul_n274) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U55 ( .A(
        SBOX_Inst_f4_multd_L_summul_n237), .B(SBOX_Inst_f4_multd_L_summul_n236), .ZN(SBOX_Inst_f4_multd_L_Orig_p[0]) );
  OAI22_X1 SBOX_Inst_f4_multd_L_summul_U54 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n268), .A2(SBOX_Inst_f4_multd_L_sB[4]), 
        .B1(SBOX_Inst_f4_multd_L_summul_n255), .B2(
        SBOX_Inst_f4_multd_L_summul_n235), .ZN(
        SBOX_Inst_f4_multd_L_summul_n236) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U53 ( .A1(SBOX_Inst_f4_multd_L_sA[4]), 
        .A2(SBOX_Inst_f4_multd_L_sB[4]), .ZN(SBOX_Inst_f4_multd_L_summul_n235)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U52 ( .A(
        SBOX_Inst_f4_multd_L_summul_n234), .B(SBOX_Inst_f4_multd_L_summul_n233), .ZN(SBOX_Inst_f4_multd_L_summul_n237) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U51 ( .A(
        SBOX_Inst_f4_multd_L_summul_n232), .B(SBOX_Inst_f4_multd_L_summul_n231), .ZN(SBOX_Inst_f4_multd_L_summul_n234) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U50 ( .A(
        SBOX_Inst_f4_multd_L_summul_n230), .B(SBOX_Inst_f4_multd_L_summul_n229), .ZN(SBOX_Inst_f4_multd_L_summul_n231) );
  AOI21_X1 SBOX_Inst_f4_multd_L_summul_U49 ( .B1(SBOX_Inst_f4_multd_L_sB[4]), 
        .B2(SBOX_Inst_f4_multd_L_summul_n228), .A(
        SBOX_Inst_f4_multd_L_summul_n227), .ZN(
        SBOX_Inst_f4_multd_L_summul_n229) );
  OAI21_X1 SBOX_Inst_f4_multd_L_summul_U48 ( .B1(SBOX_Inst_f4_multd_L_sB[4]), 
        .B2(SBOX_Inst_f4_multd_L_summul_n228), .A(SBOX_Inst_f4_multd_L_sA[3]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n227) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U47 ( .A1(SBOX_Inst_f4_multd_L_sB[5]), 
        .A2(SBOX_Inst_f4_multd_L_sB[3]), .B1(SBOX_Inst_f4_multd_L_summul_n283), 
        .B2(SBOX_Inst_f4_multd_L_summul_n255), .ZN(
        SBOX_Inst_f4_multd_L_summul_n228) );
  OAI221_X1 SBOX_Inst_f4_multd_L_summul_U46 ( .B1(SBOX_Inst_f4_multd_L_sB[5]), 
        .B2(SBOX_Inst_f4_multd_L_sB[2]), .C1(SBOX_Inst_f4_multd_L_summul_n255), 
        .C2(SBOX_Inst_f4_multd_L_summul_n290), .A(SBOX_Inst_f4_multd_L_sA[2]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n230) );
  OAI221_X1 SBOX_Inst_f4_multd_L_summul_U45 ( .B1(SBOX_Inst_f4_multd_L_sA[3]), 
        .B2(SBOX_Inst_f4_multd_L_sA[5]), .C1(SBOX_Inst_f4_multd_L_summul_n282), 
        .C2(SBOX_Inst_f4_multd_L_summul_n266), .A(SBOX_Inst_f4_multd_L_sB[2]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n232) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U44 ( .A(
        SBOX_Inst_f4_multd_L_summul_n226), .B(SBOX_Inst_f4_multd_L_summul_n225), .ZN(SBOX_Inst_f4_multd_L_Orig_p[3]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U43 ( .A(
        SBOX_Inst_f4_multd_L_summul_n221), .B(SBOX_Inst_f4_multd_L_summul_n223), .ZN(SBOX_Inst_f4_multd_L_summul_n226) );
  OAI221_X1 SBOX_Inst_f4_multd_L_summul_U42 ( .B1(
        SBOX_Inst_f4_multd_L_summul_n215), .B2(SBOX_Inst_f4_multd_L_sA[1]), 
        .C1(SBOX_Inst_f4_multd_L_summul_n224), .C2(
        SBOX_Inst_f4_multd_L_summul_n286), .A(SBOX_Inst_f4_multd_L_sB[4]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n225) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U41 ( .A(SBOX_Inst_f4_multd_L_summul_n215), .ZN(SBOX_Inst_f4_multd_L_summul_n224) );
  OAI21_X1 SBOX_Inst_f4_multd_L_summul_U40 ( .B1(
        SBOX_Inst_f4_multd_L_summul_n268), .B2(
        SBOX_Inst_f4_multd_L_summul_n267), .A(SBOX_Inst_f4_multd_L_summul_n222), .ZN(SBOX_Inst_f4_multd_L_summul_n223) );
  NAND3_X1 SBOX_Inst_f4_multd_L_summul_U39 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n268), .A2(SBOX_Inst_f4_multd_L_sA[4]), 
        .A3(SBOX_Inst_f4_multd_L_summul_n266), .ZN(
        SBOX_Inst_f4_multd_L_summul_n222) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U38 ( .A(
        SBOX_Inst_f4_multd_L_summul_n219), .B(SBOX_Inst_f4_multd_L_summul_n220), .ZN(SBOX_Inst_f4_multd_L_summul_n221) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U37 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n215), .A2(SBOX_Inst_f4_multd_L_sB[5]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n220) );
  XOR2_X1 SBOX_Inst_f4_multd_L_summul_U36 ( .A(
        SBOX_Inst_f4_multd_L_summul_n265), .B(SBOX_Inst_f4_multd_L_summul_n218), .Z(SBOX_Inst_f4_multd_L_summul_n219) );
  XOR2_X1 SBOX_Inst_f4_multd_L_summul_U35 ( .A(
        SBOX_Inst_f4_multd_L_summul_n216), .B(SBOX_Inst_f4_multd_L_summul_n217), .Z(SBOX_Inst_f4_multd_L_summul_n218) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U34 ( .A1(SBOX_Inst_f4_multd_L_sB[0]), 
        .A2(SBOX_Inst_f4_multd_L_sA[4]), .ZN(SBOX_Inst_f4_multd_L_summul_n217)
         );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U33 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n287), .A2(SBOX_Inst_f4_multd_L_sA[1]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n216) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U32 ( .A1(SBOX_Inst_f4_multd_L_sA[5]), 
        .A2(SBOX_Inst_f4_multd_L_sA[0]), .B1(SBOX_Inst_f4_multd_L_summul_n266), 
        .B2(SBOX_Inst_f4_multd_L_summul_n291), .ZN(
        SBOX_Inst_f4_multd_L_summul_n215) );
  AOI221_X1 SBOX_Inst_f4_multd_L_summul_U31 ( .B1(SBOX_Inst_f4_multd_L_sA[2]), 
        .B2(SBOX_Inst_f4_multd_L_sA[0]), .C1(SBOX_Inst_f4_multd_L_summul_n292), 
        .C2(SBOX_Inst_f4_multd_L_summul_n291), .A(
        SBOX_Inst_f4_multd_L_summul_n290), .ZN(
        SBOX_Inst_f4_multd_L_summul_n293) );
  NOR2_X1 SBOX_Inst_f4_multd_L_summul_U30 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n287), .A2(
        SBOX_Inst_f4_multd_L_summul_n286), .ZN(
        SBOX_Inst_f4_multd_L_summul_n296) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U29 ( .A(
        SBOX_Inst_f4_multd_L_summul_n285), .B(SBOX_Inst_f4_multd_L_summul_n284), .ZN(SBOX_Inst_f4_multd_L_summul_n298) );
  NOR2_X1 SBOX_Inst_f4_multd_L_summul_U28 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n292), .A2(
        SBOX_Inst_f4_multd_L_summul_n274), .ZN(
        SBOX_Inst_f4_multd_L_summul_n275) );
  NOR2_X1 SBOX_Inst_f4_multd_L_summul_U27 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n286), .A2(SBOX_Inst_f4_multd_L_sB[3]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n276) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U26 ( .A1(SBOX_Inst_f4_multd_L_sA[3]), 
        .A2(SBOX_Inst_f4_multd_L_sA[1]), .B1(SBOX_Inst_f4_multd_L_summul_n286), 
        .B2(SBOX_Inst_f4_multd_L_summul_n282), .ZN(
        SBOX_Inst_f4_multd_L_summul_n277) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U25 ( .A(
        SBOX_Inst_f4_multd_L_summul_n273), .B(SBOX_Inst_f4_multd_L_summul_n285), .ZN(SBOX_Inst_f4_multd_L_summul_n281) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U24 ( .A1(SBOX_Inst_f4_multd_L_sA[0]), 
        .A2(SBOX_Inst_f4_multd_L_sB[5]), .ZN(SBOX_Inst_f4_multd_L_summul_n261)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_summul_U23 ( .A(
        SBOX_Inst_f4_multd_L_summul_n273), .B(SBOX_Inst_f4_multd_L_summul_n265), .ZN(SBOX_Inst_f4_multd_L_summul_n264) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U22 ( .A(SBOX_Inst_f4_multd_L_summul_n239), .ZN(SBOX_Inst_f4_multd_L_summul_n238) );
  NOR2_X1 SBOX_Inst_f4_multd_L_summul_U21 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n239), .A2(
        SBOX_Inst_f4_multd_L_summul_n266), .ZN(
        SBOX_Inst_f4_multd_L_summul_n241) );
  AOI221_X1 SBOX_Inst_f4_multd_L_summul_U20 ( .B1(SBOX_Inst_f4_multd_L_sA[4]), 
        .B2(SBOX_Inst_f4_multd_L_sA[2]), .C1(SBOX_Inst_f4_multd_L_summul_n245), 
        .C2(SBOX_Inst_f4_multd_L_summul_n292), .A(
        SBOX_Inst_f4_multd_L_summul_n274), .ZN(
        SBOX_Inst_f4_multd_L_summul_n249) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U19 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n267), .A2(SBOX_Inst_f4_multd_L_sB[3]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n233) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U18 ( .A(SBOX_Inst_f4_multd_L_sA[1]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n286) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U17 ( .A(SBOX_Inst_f4_multd_L_sA[2]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n292) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U16 ( .A1(SBOX_Inst_f4_multd_L_sA[0]), 
        .A2(SBOX_Inst_f4_multd_L_sB[3]), .ZN(SBOX_Inst_f4_multd_L_summul_n269)
         );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U15 ( .A1(SBOX_Inst_f4_multd_L_sA[1]), 
        .A2(SBOX_Inst_f4_multd_L_sB[2]), .ZN(SBOX_Inst_f4_multd_L_summul_n270)
         );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U14 ( .A(SBOX_Inst_f4_multd_L_sA[3]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n282) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U13 ( .A(SBOX_Inst_f4_multd_L_sB[0]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n288) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U12 ( .A(SBOX_Inst_f4_multd_L_sB[3]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n283) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U11 ( .A(SBOX_Inst_f4_multd_L_sB[2]), 
        .ZN(SBOX_Inst_f4_multd_L_summul_n290) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U10 ( .A1(SBOX_Inst_f4_multd_L_sA[2]), 
        .A2(SBOX_Inst_f4_multd_L_sA[0]), .B1(SBOX_Inst_f4_multd_L_summul_n291), 
        .B2(SBOX_Inst_f4_multd_L_summul_n292), .ZN(
        SBOX_Inst_f4_multd_L_summul_n289) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U9 ( .A(SBOX_Inst_f4_multd_L_sA[0]), .ZN(
        SBOX_Inst_f4_multd_L_summul_n291) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U8 ( .A(SBOX_Inst_f4_multd_L_sB[1]), .ZN(
        SBOX_Inst_f4_multd_L_summul_n287) );
  NAND2_X1 SBOX_Inst_f4_multd_L_summul_U7 ( .A1(SBOX_Inst_f4_multd_L_sB[1]), 
        .A2(SBOX_Inst_f4_multd_L_sA[0]), .ZN(SBOX_Inst_f4_multd_L_summul_n250)
         );
  NOR2_X1 SBOX_Inst_f4_multd_L_summul_U6 ( .A1(
        SBOX_Inst_f4_multd_L_summul_n245), .A2(
        SBOX_Inst_f4_multd_L_summul_n255), .ZN(
        SBOX_Inst_f4_multd_L_summul_n268) );
  AOI22_X1 SBOX_Inst_f4_multd_L_summul_U5 ( .A1(SBOX_Inst_f4_multd_L_sA[4]), 
        .A2(SBOX_Inst_f4_multd_L_sA[5]), .B1(SBOX_Inst_f4_multd_L_summul_n266), 
        .B2(SBOX_Inst_f4_multd_L_summul_n245), .ZN(
        SBOX_Inst_f4_multd_L_summul_n267) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U4 ( .A(SBOX_Inst_f4_multd_L_sA[5]), .ZN(
        SBOX_Inst_f4_multd_L_summul_n266) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U3 ( .A(SBOX_Inst_f4_multd_L_sB[5]), .ZN(
        SBOX_Inst_f4_multd_L_summul_n255) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U2 ( .A(SBOX_Inst_f4_multd_L_sB[4]), .ZN(
        SBOX_Inst_f4_multd_L_summul_n254) );
  INV_X1 SBOX_Inst_f4_multd_L_summul_U1 ( .A(SBOX_Inst_f4_multd_L_sA[4]), .ZN(
        SBOX_Inst_f4_multd_L_summul_n245) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U8 ( .A(PRNGQ[45]), .B(
        SBOX_Inst_f4_multd_L_Orig_p[5]), .ZN(
        SBOX_Inst_f4_multd_L_AddNewMaskp_n6) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U7 ( .A(PRNGQ[44]), .B(
        SBOX_Inst_f4_multd_L_Orig_p[4]), .ZN(
        SBOX_Inst_f4_multd_L_AddNewMaskp_n5) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U6 ( .A(PRNGQ[46]), .B(
        SBOX_Inst_f4_multd_L_Orig_p[2]), .Z(SBOX_p_L[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U5 ( .A(PRNGQ[45]), .B(
        SBOX_Inst_f4_multd_L_Orig_p[1]), .Z(SBOX_p_L[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U4 ( .A(PRNGQ[44]), .B(
        SBOX_Inst_f4_multd_L_Orig_p[0]), .Z(SBOX_p_L[0]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U3 ( .A(PRNGQ[47]), .B(
        SBOX_Inst_f4_multd_L_Orig_p[3]), .Z(SBOX_p_L[3]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U2 ( .A(
        SBOX_Inst_f4_multd_L_AddNewMaskp_n6), .B(PRNGQ[47]), .ZN(SBOX_p_L[5])
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskp_U1 ( .A(
        SBOX_Inst_f4_multd_L_AddNewMaskp_n5), .B(PRNGQ[46]), .ZN(SBOX_p_L[4])
         );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U93 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n294), .B(SBOX_Inst_f4_multd_L_lowmul_n293), .ZN(SBOX_Inst_f4_multd_L_lowmul_n302) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U92 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n292), .B(SBOX_Inst_f4_multd_L_lowmul_n291), .ZN(SBOX_Inst_f4_multd_L_lowmul_n293) );
  AOI221_X1 SBOX_Inst_f4_multd_L_lowmul_U91 ( .B1(SBOX_FF3_out[1]), .B2(
        SBOX_FF3_out[5]), .C1(SBOX_Inst_f4_multd_L_lowmul_n290), .C2(
        SBOX_Inst_f4_multd_L_lowmul_n289), .A(SBOX_Inst_f4_multd_L_lowmul_n299), .ZN(SBOX_Inst_f4_multd_L_lowmul_n294) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U90 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n285), .B(SBOX_Inst_f4_multd_L_lowmul_n284), .ZN(SBOX_Inst_f4_multd_L_Orig_pl[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U89 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n282), .B(SBOX_Inst_f4_multd_L_lowmul_n281), .Z(SBOX_Inst_f4_multd_L_lowmul_n295) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U88 ( .A1(SBOX_FF3_out[1]), .A2(
        SBOX_FF3_out[24]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n281) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U87 ( .A1(SBOX_FF3_out[0]), .A2(
        SBOX_FF3_out[25]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n282) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U86 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n280), .B(SBOX_Inst_f4_multd_L_lowmul_n279), .ZN(SBOX_Inst_f4_multd_L_lowmul_n283) );
  AOI22_X1 SBOX_Inst_f4_multd_L_lowmul_U85 ( .A1(SBOX_FF3_out[0]), .A2(
        SBOX_FF3_out[25]), .B1(SBOX_Inst_f4_multd_L_lowmul_n297), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n278), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n279) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U84 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n276), .B(SBOX_Inst_f4_multd_L_lowmul_n275), .ZN(SBOX_Inst_f4_multd_L_lowmul_n277) );
  AOI21_X1 SBOX_Inst_f4_multd_L_lowmul_U83 ( .B1(
        SBOX_Inst_f4_multd_L_lowmul_n274), .B2(SBOX_FF3_out[8]), .A(
        SBOX_Inst_f4_multd_L_lowmul_n273), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n275) );
  OAI21_X1 SBOX_Inst_f4_multd_L_lowmul_U82 ( .B1(
        SBOX_Inst_f4_multd_L_lowmul_n274), .B2(SBOX_FF3_out[8]), .A(
        SBOX_FF3_out[33]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n273) );
  AOI22_X1 SBOX_Inst_f4_multd_L_lowmul_U81 ( .A1(SBOX_FF3_out[1]), .A2(
        SBOX_FF3_out[9]), .B1(SBOX_Inst_f4_multd_L_lowmul_n288), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n290), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n274) );
  AOI22_X1 SBOX_Inst_f4_multd_L_lowmul_U80 ( .A1(SBOX_FF3_out[25]), .A2(
        SBOX_FF3_out[9]), .B1(SBOX_FF3_out[8]), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n297), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n276) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U79 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n272), .B(SBOX_Inst_f4_multd_L_lowmul_n271), .ZN(SBOX_Inst_f4_multd_L_Orig_pl[1]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U78 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n270), .B(SBOX_Inst_f4_multd_L_lowmul_n269), .ZN(SBOX_Inst_f4_multd_L_lowmul_n271) );
  OAI221_X1 SBOX_Inst_f4_multd_L_lowmul_U77 ( .B1(SBOX_FF3_out[5]), .B2(
        SBOX_FF3_out[4]), .C1(SBOX_Inst_f4_multd_L_lowmul_n289), .C2(
        SBOX_Inst_f4_multd_L_lowmul_n268), .A(SBOX_FF3_out[29]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n269) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U76 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n267), .B(SBOX_Inst_f4_multd_L_lowmul_n266), .ZN(SBOX_Inst_f4_multd_L_lowmul_n270) );
  OAI221_X1 SBOX_Inst_f4_multd_L_lowmul_U75 ( .B1(SBOX_FF3_out[28]), .B2(
        SBOX_FF3_out[29]), .C1(SBOX_Inst_f4_multd_L_lowmul_n300), .C2(
        SBOX_Inst_f4_multd_L_lowmul_n298), .A(SBOX_FF3_out[8]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n266) );
  OAI221_X1 SBOX_Inst_f4_multd_L_lowmul_U74 ( .B1(SBOX_FF3_out[32]), .B2(
        SBOX_FF3_out[28]), .C1(SBOX_Inst_f4_multd_L_lowmul_n265), .C2(
        SBOX_Inst_f4_multd_L_lowmul_n300), .A(SBOX_Inst_f4_multd_L_lowmul_n296), .ZN(SBOX_Inst_f4_multd_L_lowmul_n267) );
  AOI22_X1 SBOX_Inst_f4_multd_L_lowmul_U73 ( .A1(SBOX_FF3_out[5]), .A2(
        SBOX_FF3_out[4]), .B1(SBOX_Inst_f4_multd_L_lowmul_n268), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n289), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n296) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U72 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n264), .B(SBOX_Inst_f4_multd_L_lowmul_n263), .ZN(SBOX_Inst_f4_multd_L_lowmul_n272) );
  AOI221_X1 SBOX_Inst_f4_multd_L_lowmul_U71 ( .B1(SBOX_FF3_out[33]), .B2(
        SBOX_FF3_out[28]), .C1(SBOX_FF3_out[4]), .C2(SBOX_FF3_out[9]), .A(
        SBOX_Inst_f4_multd_L_lowmul_n258), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n264) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U70 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n257), .B(SBOX_Inst_f4_multd_L_lowmul_n256), .ZN(SBOX_Inst_f4_multd_L_Orig_pl[0]) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U69 ( .A1(SBOX_FF3_out[5]), .A2(
        SBOX_Inst_f4_multd_L_lowmul_n260), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n256) );
  OAI21_X1 SBOX_Inst_f4_multd_L_lowmul_U68 ( .B1(SBOX_FF3_out[32]), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n287), .A(SBOX_Inst_f4_multd_L_lowmul_n261), .ZN(SBOX_Inst_f4_multd_L_lowmul_n260) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U67 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n255), .B(SBOX_Inst_f4_multd_L_lowmul_n254), .Z(SBOX_Inst_f4_multd_L_lowmul_n257) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U66 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n253), .B(SBOX_Inst_f4_multd_L_lowmul_n252), .ZN(SBOX_Inst_f4_multd_L_lowmul_n254) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U65 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n250), .B(SBOX_Inst_f4_multd_L_lowmul_n249), .ZN(SBOX_Inst_f4_multd_L_lowmul_n251) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U64 ( .A(SBOX_FF3_out[9]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n288) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U63 ( .A1(
        SBOX_Inst_f4_multd_L_lowmul_n298), .A2(SBOX_FF3_out[8]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n250) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U62 ( .A(SBOX_FF3_out[4]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n268) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U61 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n248), .B(SBOX_Inst_f4_multd_L_lowmul_n247), .ZN(SBOX_Inst_f4_multd_L_Orig_pl[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U60 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n295), .B(SBOX_Inst_f4_multd_L_lowmul_n244), .ZN(SBOX_Inst_f4_multd_L_lowmul_n248) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U59 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n245), .B(SBOX_Inst_f4_multd_L_lowmul_n246), .Z(SBOX_Inst_f4_multd_L_lowmul_n247) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U58 ( .A1(
        SBOX_Inst_f4_multd_L_lowmul_n296), .A2(SBOX_FF3_out[28]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n246) );
  NOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U57 ( .A1(SBOX_FF3_out[5]), .A2(
        SBOX_Inst_f4_multd_L_lowmul_n297), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n245) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U56 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n302), .B(SBOX_Inst_f4_multd_L_lowmul_n243), .ZN(SBOX_Inst_f4_multd_L_lowmul_n244) );
  MUX2_X1 SBOX_Inst_f4_multd_L_lowmul_U55 ( .A(SBOX_FF3_out[0]), .B(
        SBOX_FF3_out[1]), .S(SBOX_Inst_f4_multd_L_lowmul_n242), .Z(
        SBOX_Inst_f4_multd_L_lowmul_n243) );
  AOI22_X1 SBOX_Inst_f4_multd_L_lowmul_U54 ( .A1(SBOX_FF3_out[29]), .A2(
        SBOX_FF3_out[25]), .B1(SBOX_Inst_f4_multd_L_lowmul_n297), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n298), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n242) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U53 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n302), .B(SBOX_Inst_f4_multd_L_lowmul_n241), .ZN(SBOX_Inst_f4_multd_L_Orig_pl[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U52 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n234), .B(SBOX_Inst_f4_multd_L_lowmul_n240), .ZN(SBOX_Inst_f4_multd_L_lowmul_n241) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U51 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n239), .B(SBOX_Inst_f4_multd_L_lowmul_n238), .ZN(SBOX_Inst_f4_multd_L_lowmul_n240) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U50 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n237), .B(SBOX_Inst_f4_multd_L_lowmul_n301), .ZN(SBOX_Inst_f4_multd_L_lowmul_n239) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U49 ( .A1(SBOX_FF3_out[0]), .A2(
        SBOX_FF3_out[29]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n238) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U48 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n235), .B(SBOX_Inst_f4_multd_L_lowmul_n236), .Z(SBOX_Inst_f4_multd_L_lowmul_n237) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U47 ( .A1(SBOX_FF3_out[4]), .A2(
        SBOX_FF3_out[24]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n236) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U46 ( .A1(SBOX_FF3_out[1]), .A2(
        SBOX_FF3_out[25]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n235) );
  AOI22_X1 SBOX_Inst_f4_multd_L_lowmul_U45 ( .A1(SBOX_FF3_out[0]), .A2(
        SBOX_Inst_f4_multd_L_lowmul_n232), .B1(SBOX_FF3_out[25]), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n233), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n234) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U44 ( .A(SBOX_FF3_out[0]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n233) );
  OAI22_X1 SBOX_Inst_f4_multd_L_lowmul_U43 ( .A1(SBOX_FF3_out[24]), .A2(
        SBOX_Inst_f4_multd_L_lowmul_n300), .B1(SBOX_FF3_out[28]), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n299), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n232) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U42 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n230), .B(SBOX_Inst_f4_multd_L_lowmul_n231), .ZN(SBOX_Inst_f4_multd_L_lowmul_n301) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U41 ( .A1(SBOX_FF3_out[28]), .A2(
        SBOX_FF3_out[4]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n231) );
  NOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U40 ( .A1(
        SBOX_Inst_f4_multd_L_lowmul_n289), .A2(
        SBOX_Inst_f4_multd_L_lowmul_n298), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n230) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U39 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n228), .B(SBOX_Inst_f4_multd_L_lowmul_n229), .Z(SBOX_Inst_f4_multd_L_lowmul_n286) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U38 ( .A1(SBOX_FF3_out[0]), .A2(
        SBOX_FF3_out[33]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n229) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U37 ( .A1(SBOX_FF3_out[32]), .A2(
        SBOX_FF3_out[1]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n228) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U36 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n226), .B(SBOX_Inst_f4_multd_L_lowmul_n227), .Z(SBOX_Inst_f4_multd_L_Orig_pl[3]) );
  OAI221_X1 SBOX_Inst_f4_multd_L_lowmul_U35 ( .B1(
        SBOX_Inst_f4_multd_L_lowmul_n217), .B2(SBOX_FF3_out[25]), .C1(
        SBOX_Inst_f4_multd_L_lowmul_n216), .C2(
        SBOX_Inst_f4_multd_L_lowmul_n297), .A(SBOX_FF3_out[8]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n227) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U34 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n224), .B(SBOX_Inst_f4_multd_L_lowmul_n225), .ZN(SBOX_Inst_f4_multd_L_lowmul_n226) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U33 ( .A1(
        SBOX_Inst_f4_multd_L_lowmul_n288), .A2(SBOX_FF3_out[32]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n225) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U32 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n223), .B(SBOX_Inst_f4_multd_L_lowmul_n287), .Z(SBOX_Inst_f4_multd_L_lowmul_n224) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U31 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n221), .B(SBOX_Inst_f4_multd_L_lowmul_n222), .ZN(SBOX_Inst_f4_multd_L_lowmul_n223) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U30 ( .A1(
        SBOX_Inst_f4_multd_L_lowmul_n217), .A2(SBOX_FF3_out[9]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n222) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U29 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n220), .B(SBOX_Inst_f4_multd_L_lowmul_n286), .Z(SBOX_Inst_f4_multd_L_lowmul_n221) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U28 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n218), .B(SBOX_Inst_f4_multd_L_lowmul_n219), .Z(SBOX_Inst_f4_multd_L_lowmul_n220) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U27 ( .A1(
        SBOX_Inst_f4_multd_L_lowmul_n290), .A2(SBOX_FF3_out[25]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n219) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U26 ( .A1(SBOX_FF3_out[32]), .A2(
        SBOX_FF3_out[0]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n218) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U25 ( .A(SBOX_Inst_f4_multd_L_lowmul_n216), .ZN(SBOX_Inst_f4_multd_L_lowmul_n217) );
  OAI22_X1 SBOX_Inst_f4_multd_L_lowmul_U24 ( .A1(SBOX_FF3_out[24]), .A2(
        SBOX_FF3_out[33]), .B1(SBOX_Inst_f4_multd_L_lowmul_n287), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n299), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n216) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U23 ( .A(SBOX_FF3_out[0]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n278) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U22 ( .A1(SBOX_FF3_out[24]), .A2(
        SBOX_FF3_out[9]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n280) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U21 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n277), .B(SBOX_Inst_f4_multd_L_lowmul_n286), .Z(SBOX_Inst_f4_multd_L_lowmul_n285) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U20 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n283), .B(SBOX_Inst_f4_multd_L_lowmul_n295), .ZN(SBOX_Inst_f4_multd_L_lowmul_n284) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U19 ( .A1(SBOX_FF3_out[32]), .A2(
        SBOX_FF3_out[8]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n259) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U18 ( .A(SBOX_Inst_f4_multd_L_lowmul_n259), .ZN(SBOX_Inst_f4_multd_L_lowmul_n262) );
  OAI22_X1 SBOX_Inst_f4_multd_L_lowmul_U17 ( .A1(SBOX_FF3_out[33]), .A2(
        SBOX_FF3_out[28]), .B1(SBOX_FF3_out[9]), .B2(SBOX_FF3_out[4]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n258) );
  AOI22_X1 SBOX_Inst_f4_multd_L_lowmul_U16 ( .A1(
        SBOX_Inst_f4_multd_L_lowmul_n262), .A2(
        SBOX_Inst_f4_multd_L_lowmul_n261), .B1(
        SBOX_Inst_f4_multd_L_lowmul_n260), .B2(
        SBOX_Inst_f4_multd_L_lowmul_n259), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n263) );
  AOI221_X1 SBOX_Inst_f4_multd_L_lowmul_U15 ( .B1(SBOX_FF3_out[32]), .B2(
        SBOX_FF3_out[28]), .C1(SBOX_Inst_f4_multd_L_lowmul_n265), .C2(
        SBOX_Inst_f4_multd_L_lowmul_n300), .A(SBOX_Inst_f4_multd_L_lowmul_n288), .ZN(SBOX_Inst_f4_multd_L_lowmul_n249) );
  XOR2_X1 SBOX_Inst_f4_multd_L_lowmul_U14 ( .A(
        SBOX_Inst_f4_multd_L_lowmul_n301), .B(SBOX_Inst_f4_multd_L_lowmul_n251), .Z(SBOX_Inst_f4_multd_L_lowmul_n253) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U13 ( .A1(SBOX_FF3_out[29]), .A2(
        SBOX_FF3_out[9]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n252) );
  AOI221_X1 SBOX_Inst_f4_multd_L_lowmul_U12 ( .B1(SBOX_FF3_out[33]), .B2(
        SBOX_FF3_out[29]), .C1(SBOX_Inst_f4_multd_L_lowmul_n287), .C2(
        SBOX_Inst_f4_multd_L_lowmul_n298), .A(SBOX_Inst_f4_multd_L_lowmul_n268), .ZN(SBOX_Inst_f4_multd_L_lowmul_n255) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U11 ( .A1(SBOX_FF3_out[4]), .A2(
        SBOX_FF3_out[25]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n292) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U10 ( .A1(SBOX_FF3_out[28]), .A2(
        SBOX_FF3_out[1]), .ZN(SBOX_Inst_f4_multd_L_lowmul_n291) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U9 ( .A(SBOX_FF3_out[28]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n300) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U8 ( .A(SBOX_FF3_out[24]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n299) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U7 ( .A(SBOX_FF3_out[25]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n297) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U6 ( .A(SBOX_FF3_out[29]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n298) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U5 ( .A(SBOX_FF3_out[33]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n287) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U4 ( .A(SBOX_FF3_out[1]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n290) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U3 ( .A(SBOX_FF3_out[5]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n289) );
  NAND2_X1 SBOX_Inst_f4_multd_L_lowmul_U2 ( .A1(SBOX_FF3_out[32]), .A2(
        SBOX_Inst_f4_multd_L_lowmul_n287), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n261) );
  INV_X1 SBOX_Inst_f4_multd_L_lowmul_U1 ( .A(SBOX_FF3_out[32]), .ZN(
        SBOX_Inst_f4_multd_L_lowmul_n265) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U8 ( .A(PRNGQ[50]), .B(
        SBOX_Inst_f4_multd_L_Orig_pl[2]), .Z(SBOX_pl_L[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U7 ( .A(PRNGQ[49]), .B(
        SBOX_Inst_f4_multd_L_Orig_pl[1]), .Z(SBOX_pl_L[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U6 ( .A(PRNGQ[48]), .B(
        SBOX_Inst_f4_multd_L_Orig_pl[0]), .Z(SBOX_pl_L[0]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U5 ( .A(
        SBOX_Inst_f4_multd_L_AddNewMaskpl_n6), .B(PRNGQ[50]), .ZN(SBOX_pl_L[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U4 ( .A(PRNGQ[48]), .B(
        SBOX_Inst_f4_multd_L_Orig_pl[4]), .ZN(
        SBOX_Inst_f4_multd_L_AddNewMaskpl_n6) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U3 ( .A(
        SBOX_Inst_f4_multd_L_AddNewMaskpl_n5), .B(PRNGQ[51]), .ZN(SBOX_pl_L[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U2 ( .A(PRNGQ[49]), .B(
        SBOX_Inst_f4_multd_L_Orig_pl[5]), .ZN(
        SBOX_Inst_f4_multd_L_AddNewMaskpl_n5) );
  XOR2_X1 SBOX_Inst_f4_multd_L_AddNewMaskpl_U1 ( .A(PRNGQ[51]), .B(
        SBOX_Inst_f4_multd_L_Orig_pl[3]), .Z(SBOX_pl_L[3]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_U12 ( .A(SBOX_FF3_out[11]), .B(SBOX_FF3_out[9]), 
        .Z(SBOX_Inst_f4_multd_H_sA[5]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_U11 ( .A(SBOX_FF3_out[4]), .B(SBOX_FF3_out[6]), 
        .Z(SBOX_Inst_f4_multd_H_sA[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_U10 ( .A(SBOX_FF3_out[1]), .B(SBOX_FF3_out[3]), 
        .Z(SBOX_Inst_f4_multd_H_sA[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_U9 ( .A(SBOX_FF3_out[0]), .B(SBOX_FF3_out[2]), 
        .Z(SBOX_Inst_f4_multd_H_sA[0]) );
  XOR2_X2 SBOX_Inst_f4_multd_H_U8 ( .A(SBOX_FF3_out[10]), .B(SBOX_FF3_out[8]), 
        .Z(SBOX_Inst_f4_multd_H_sA[4]) );
  XOR2_X2 SBOX_Inst_f4_multd_H_U7 ( .A(SBOX_FF3_out[12]), .B(SBOX_FF3_out[14]), 
        .Z(SBOX_Inst_f4_multd_H_sB[0]) );
  XOR2_X2 SBOX_Inst_f4_multd_H_U6 ( .A(SBOX_FF3_out[17]), .B(SBOX_FF3_out[19]), 
        .Z(SBOX_Inst_f4_multd_H_sB[3]) );
  XOR2_X2 SBOX_Inst_f4_multd_H_U5 ( .A(SBOX_FF3_out[22]), .B(SBOX_FF3_out[20]), 
        .Z(SBOX_Inst_f4_multd_H_sB[4]) );
  XOR2_X2 SBOX_Inst_f4_multd_H_U4 ( .A(SBOX_FF3_out[23]), .B(SBOX_FF3_out[21]), 
        .Z(SBOX_Inst_f4_multd_H_sB[5]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_U3 ( .A(SBOX_FF3_out[13]), .B(SBOX_FF3_out[15]), 
        .Z(SBOX_Inst_f4_multd_H_sB[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_U2 ( .A(SBOX_FF3_out[5]), .B(SBOX_FF3_out[7]), 
        .Z(SBOX_Inst_f4_multd_H_sA[3]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_U1 ( .A(SBOX_FF3_out[16]), .B(SBOX_FF3_out[18]), 
        .Z(SBOX_Inst_f4_multd_H_sB[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U100 ( .A(
        SBOX_Inst_f4_multd_H_himul_n296), .B(SBOX_Inst_f4_multd_H_himul_n295), 
        .ZN(SBOX_Inst_f4_multd_H_himul_n301) );
  XOR2_X1 SBOX_Inst_f4_multd_H_himul_U99 ( .A(SBOX_Inst_f4_multd_H_himul_n294), 
        .B(SBOX_Inst_f4_multd_H_himul_n293), .Z(
        SBOX_Inst_f4_multd_H_himul_n295) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U98 ( .A1(SBOX_FF3_out[6]), .A2(
        SBOX_FF3_out[2]), .B1(SBOX_Inst_f4_multd_H_himul_n307), .B2(
        SBOX_Inst_f4_multd_H_himul_n308), .ZN(SBOX_Inst_f4_multd_H_himul_n305)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U97 ( .A(SBOX_Inst_f4_multd_H_himul_n288), .B(SBOX_Inst_f4_multd_H_himul_n287), .ZN(SBOX_Inst_f4_multd_H_Orig_ph[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U96 ( .A(SBOX_Inst_f4_multd_H_himul_n286), .B(SBOX_Inst_f4_multd_H_himul_n285), .ZN(SBOX_Inst_f4_multd_H_himul_n287) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U95 ( .A1(SBOX_FF3_out[2]), .A2(
        SBOX_FF3_out[23]), .ZN(SBOX_Inst_f4_multd_H_himul_n285) );
  XOR2_X1 SBOX_Inst_f4_multd_H_himul_U94 ( .A(SBOX_Inst_f4_multd_H_himul_n284), 
        .B(SBOX_Inst_f4_multd_H_himul_n283), .Z(
        SBOX_Inst_f4_multd_H_himul_n286) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U93 ( .A(SBOX_Inst_f4_multd_H_himul_n282), .B(SBOX_Inst_f4_multd_H_himul_n281), .ZN(SBOX_Inst_f4_multd_H_himul_n283) );
  MUX2_X1 SBOX_Inst_f4_multd_H_himul_U92 ( .A(SBOX_FF3_out[22]), .B(
        SBOX_Inst_f4_multd_H_himul_n280), .S(SBOX_FF3_out[11]), .Z(
        SBOX_Inst_f4_multd_H_himul_n281) );
  OAI221_X1 SBOX_Inst_f4_multd_H_himul_U91 ( .B1(SBOX_FF3_out[23]), .B2(
        SBOX_FF3_out[22]), .C1(SBOX_Inst_f4_multd_H_himul_n279), .C2(
        SBOX_Inst_f4_multd_H_himul_n278), .A(SBOX_FF3_out[3]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n282) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U90 ( .A1(SBOX_FF3_out[3]), .A2(
        SBOX_FF3_out[14]), .B1(SBOX_Inst_f4_multd_H_himul_n304), .B2(
        SBOX_Inst_f4_multd_H_himul_n302), .ZN(SBOX_Inst_f4_multd_H_himul_n284)
         );
  XOR2_X1 SBOX_Inst_f4_multd_H_himul_U89 ( .A(SBOX_Inst_f4_multd_H_himul_n277), 
        .B(SBOX_Inst_f4_multd_H_himul_n276), .Z(
        SBOX_Inst_f4_multd_H_himul_n289) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U88 ( .A1(SBOX_FF3_out[15]), .A2(
        SBOX_FF3_out[10]), .ZN(SBOX_Inst_f4_multd_H_himul_n276) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U87 ( .A1(SBOX_FF3_out[14]), .A2(
        SBOX_FF3_out[11]), .ZN(SBOX_Inst_f4_multd_H_himul_n277) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U86 ( .A1(SBOX_FF3_out[10]), .A2(
        SBOX_FF3_out[11]), .B1(SBOX_Inst_f4_multd_H_himul_n290), .B2(
        SBOX_Inst_f4_multd_H_himul_n275), .ZN(SBOX_Inst_f4_multd_H_himul_n291)
         );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U85 ( .A(SBOX_FF3_out[11]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n290) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U84 ( .A(SBOX_Inst_f4_multd_H_himul_n272), .B(SBOX_Inst_f4_multd_H_himul_n274), .ZN(SBOX_Inst_f4_multd_H_Orig_ph[1]) );
  AOI211_X1 SBOX_Inst_f4_multd_H_himul_U83 ( .C1(SBOX_FF3_out[10]), .C2(
        SBOX_FF3_out[6]), .A(SBOX_Inst_f4_multd_H_himul_n298), .B(
        SBOX_Inst_f4_multd_H_himul_n273), .ZN(SBOX_Inst_f4_multd_H_himul_n274)
         );
  AND2_X1 SBOX_Inst_f4_multd_H_himul_U82 ( .A1(SBOX_Inst_f4_multd_H_himul_n275), .A2(SBOX_Inst_f4_multd_H_himul_n308), .ZN(SBOX_Inst_f4_multd_H_himul_n273)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U81 ( .A(SBOX_Inst_f4_multd_H_himul_n271), .B(SBOX_Inst_f4_multd_H_himul_n268), .ZN(SBOX_Inst_f4_multd_H_himul_n272) );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U80 ( .A1(SBOX_Inst_f4_multd_H_himul_n270), .A2(SBOX_Inst_f4_multd_H_himul_n269), .ZN(SBOX_Inst_f4_multd_H_himul_n271)
         );
  OAI22_X1 SBOX_Inst_f4_multd_H_himul_U79 ( .A1(SBOX_FF3_out[7]), .A2(
        SBOX_FF3_out[10]), .B1(SBOX_Inst_f4_multd_H_himul_n275), .B2(
        SBOX_Inst_f4_multd_H_himul_n299), .ZN(SBOX_Inst_f4_multd_H_himul_n270)
         );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U78 ( .A(SBOX_FF3_out[22]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n269) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U77 ( .A(SBOX_Inst_f4_multd_H_himul_n266), .B(SBOX_Inst_f4_multd_H_himul_n267), .ZN(SBOX_Inst_f4_multd_H_himul_n268) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U76 ( .A(SBOX_FF3_out[10]), .B(
        SBOX_Inst_f4_multd_H_himul_n264), .ZN(SBOX_Inst_f4_multd_H_himul_n267)
         );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U75 ( .A1(SBOX_Inst_f4_multd_H_himul_n259), .A2(SBOX_Inst_f4_multd_H_himul_n265), .ZN(SBOX_Inst_f4_multd_H_himul_n266)
         );
  OAI22_X1 SBOX_Inst_f4_multd_H_himul_U74 ( .A1(SBOX_FF3_out[18]), .A2(
        SBOX_FF3_out[19]), .B1(SBOX_Inst_f4_multd_H_himul_n306), .B2(
        SBOX_Inst_f4_multd_H_himul_n300), .ZN(SBOX_Inst_f4_multd_H_himul_n265)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U73 ( .A(SBOX_Inst_f4_multd_H_himul_n263), .B(SBOX_Inst_f4_multd_H_himul_n262), .ZN(SBOX_Inst_f4_multd_H_himul_n264) );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U72 ( .A1(SBOX_Inst_f4_multd_H_himul_n260), .A2(SBOX_Inst_f4_multd_H_himul_n290), .ZN(SBOX_Inst_f4_multd_H_himul_n263)
         );
  OAI221_X1 SBOX_Inst_f4_multd_H_himul_U71 ( .B1(
        SBOX_Inst_f4_multd_H_himul_n260), .B2(SBOX_FF3_out[22]), .C1(
        SBOX_Inst_f4_multd_H_himul_n261), .C2(SBOX_Inst_f4_multd_H_himul_n278), 
        .A(SBOX_FF3_out[6]), .ZN(SBOX_Inst_f4_multd_H_himul_n262) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U70 ( .A(SBOX_Inst_f4_multd_H_himul_n260), 
        .ZN(SBOX_Inst_f4_multd_H_himul_n261) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U69 ( .A1(SBOX_FF3_out[23]), .A2(
        SBOX_FF3_out[18]), .B1(SBOX_Inst_f4_multd_H_himul_n306), .B2(
        SBOX_Inst_f4_multd_H_himul_n279), .ZN(SBOX_Inst_f4_multd_H_himul_n260)
         );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U68 ( .A(SBOX_FF3_out[7]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n259) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U67 ( .A(SBOX_Inst_f4_multd_H_himul_n257), .B(SBOX_Inst_f4_multd_H_himul_n258), .ZN(SBOX_Inst_f4_multd_H_Orig_ph[5]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_himul_U66 ( .A(SBOX_Inst_f4_multd_H_himul_n253), 
        .B(SBOX_Inst_f4_multd_H_himul_n255), .Z(
        SBOX_Inst_f4_multd_H_himul_n258) );
  AOI211_X1 SBOX_Inst_f4_multd_H_himul_U65 ( .C1(SBOX_FF3_out[14]), .C2(
        SBOX_FF3_out[19]), .A(SBOX_Inst_f4_multd_H_himul_n256), .B(
        SBOX_Inst_f4_multd_H_himul_n299), .ZN(SBOX_Inst_f4_multd_H_himul_n257)
         );
  AND2_X1 SBOX_Inst_f4_multd_H_himul_U64 ( .A1(SBOX_Inst_f4_multd_H_himul_n304), .A2(SBOX_Inst_f4_multd_H_himul_n300), .ZN(SBOX_Inst_f4_multd_H_himul_n256)
         );
  AOI211_X1 SBOX_Inst_f4_multd_H_himul_U63 ( .C1(SBOX_FF3_out[2]), .C2(
        SBOX_FF3_out[6]), .A(SBOX_Inst_f4_multd_H_himul_n306), .B(
        SBOX_Inst_f4_multd_H_himul_n254), .ZN(SBOX_Inst_f4_multd_H_himul_n255)
         );
  AND2_X1 SBOX_Inst_f4_multd_H_himul_U62 ( .A1(SBOX_Inst_f4_multd_H_himul_n307), .A2(SBOX_Inst_f4_multd_H_himul_n308), .ZN(SBOX_Inst_f4_multd_H_himul_n254)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U61 ( .A(SBOX_Inst_f4_multd_H_himul_n251), .B(SBOX_Inst_f4_multd_H_himul_n252), .ZN(SBOX_Inst_f4_multd_H_himul_n253) );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U60 ( .A1(SBOX_Inst_f4_multd_H_himul_n303), .A2(SBOX_Inst_f4_multd_H_himul_n302), .ZN(SBOX_Inst_f4_multd_H_himul_n252)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U59 ( .A(SBOX_Inst_f4_multd_H_himul_n301), .B(SBOX_Inst_f4_multd_H_himul_n250), .ZN(SBOX_Inst_f4_multd_H_himul_n251) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U58 ( .A1(SBOX_FF3_out[3]), .A2(
        SBOX_Inst_f4_multd_H_himul_n304), .B1(SBOX_FF3_out[14]), .B2(
        SBOX_Inst_f4_multd_H_himul_n305), .ZN(SBOX_Inst_f4_multd_H_himul_n250)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U57 ( .A(SBOX_Inst_f4_multd_H_himul_n249), .B(SBOX_Inst_f4_multd_H_himul_n248), .ZN(SBOX_Inst_f4_multd_H_Orig_ph[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U56 ( .A(SBOX_Inst_f4_multd_H_himul_n297), .B(SBOX_Inst_f4_multd_H_himul_n245), .ZN(SBOX_Inst_f4_multd_H_himul_n249) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U55 ( .A(SBOX_Inst_f4_multd_H_himul_n246), .B(SBOX_Inst_f4_multd_H_himul_n247), .ZN(SBOX_Inst_f4_multd_H_himul_n248) );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U54 ( .A1(SBOX_FF3_out[19]), .A2(
        SBOX_Inst_f4_multd_H_himul_n302), .ZN(SBOX_Inst_f4_multd_H_himul_n247)
         );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U53 ( .A1(SBOX_Inst_f4_multd_H_himul_n308), .A2(SBOX_Inst_f4_multd_H_himul_n298), .ZN(SBOX_Inst_f4_multd_H_himul_n246)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U52 ( .A(SBOX_Inst_f4_multd_H_himul_n301), .B(SBOX_Inst_f4_multd_H_himul_n244), .ZN(SBOX_Inst_f4_multd_H_himul_n245) );
  MUX2_X1 SBOX_Inst_f4_multd_H_himul_U51 ( .A(SBOX_FF3_out[14]), .B(
        SBOX_FF3_out[15]), .S(SBOX_Inst_f4_multd_H_himul_n243), .Z(
        SBOX_Inst_f4_multd_H_himul_n244) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U50 ( .A1(SBOX_FF3_out[7]), .A2(
        SBOX_FF3_out[3]), .B1(SBOX_Inst_f4_multd_H_himul_n302), .B2(
        SBOX_Inst_f4_multd_H_himul_n299), .ZN(SBOX_Inst_f4_multd_H_himul_n243)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U49 ( .A(SBOX_Inst_f4_multd_H_himul_n242), .B(SBOX_Inst_f4_multd_H_himul_n241), .ZN(SBOX_Inst_f4_multd_H_Orig_ph[3]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U48 ( .A(SBOX_Inst_f4_multd_H_himul_n237), .B(SBOX_Inst_f4_multd_H_himul_n239), .ZN(SBOX_Inst_f4_multd_H_himul_n242) );
  OAI221_X1 SBOX_Inst_f4_multd_H_himul_U47 ( .B1(
        SBOX_Inst_f4_multd_H_himul_n231), .B2(SBOX_FF3_out[3]), .C1(
        SBOX_Inst_f4_multd_H_himul_n240), .C2(SBOX_Inst_f4_multd_H_himul_n302), 
        .A(SBOX_FF3_out[22]), .ZN(SBOX_Inst_f4_multd_H_himul_n241) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U46 ( .A(SBOX_Inst_f4_multd_H_himul_n231), 
        .ZN(SBOX_Inst_f4_multd_H_himul_n240) );
  OAI21_X1 SBOX_Inst_f4_multd_H_himul_U45 ( .B1(
        SBOX_Inst_f4_multd_H_himul_n292), .B2(SBOX_Inst_f4_multd_H_himul_n291), 
        .A(SBOX_Inst_f4_multd_H_himul_n238), .ZN(
        SBOX_Inst_f4_multd_H_himul_n239) );
  NAND3_X1 SBOX_Inst_f4_multd_H_himul_U44 ( .A1(
        SBOX_Inst_f4_multd_H_himul_n292), .A2(SBOX_FF3_out[10]), .A3(
        SBOX_Inst_f4_multd_H_himul_n290), .ZN(SBOX_Inst_f4_multd_H_himul_n238)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U43 ( .A(SBOX_Inst_f4_multd_H_himul_n235), .B(SBOX_Inst_f4_multd_H_himul_n236), .ZN(SBOX_Inst_f4_multd_H_himul_n237) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U42 ( .A1(
        SBOX_Inst_f4_multd_H_himul_n231), .A2(SBOX_FF3_out[23]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n236) );
  XOR2_X1 SBOX_Inst_f4_multd_H_himul_U41 ( .A(SBOX_Inst_f4_multd_H_himul_n289), 
        .B(SBOX_Inst_f4_multd_H_himul_n234), .Z(
        SBOX_Inst_f4_multd_H_himul_n235) );
  XOR2_X1 SBOX_Inst_f4_multd_H_himul_U40 ( .A(SBOX_Inst_f4_multd_H_himul_n232), 
        .B(SBOX_Inst_f4_multd_H_himul_n233), .Z(
        SBOX_Inst_f4_multd_H_himul_n234) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U39 ( .A1(SBOX_FF3_out[14]), .A2(
        SBOX_FF3_out[10]), .ZN(SBOX_Inst_f4_multd_H_himul_n233) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U38 ( .A1(
        SBOX_Inst_f4_multd_H_himul_n303), .A2(SBOX_FF3_out[3]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n232) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U37 ( .A1(SBOX_FF3_out[11]), .A2(
        SBOX_FF3_out[2]), .B1(SBOX_Inst_f4_multd_H_himul_n290), .B2(
        SBOX_Inst_f4_multd_H_himul_n307), .ZN(SBOX_Inst_f4_multd_H_himul_n231)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U36 ( .A(SBOX_Inst_f4_multd_H_himul_n228), .B(SBOX_Inst_f4_multd_H_himul_n230), .ZN(SBOX_Inst_f4_multd_H_Orig_ph[0]) );
  OAI22_X1 SBOX_Inst_f4_multd_H_himul_U35 ( .A1(
        SBOX_Inst_f4_multd_H_himul_n279), .A2(SBOX_Inst_f4_multd_H_himul_n229), 
        .B1(SBOX_Inst_f4_multd_H_himul_n292), .B2(SBOX_FF3_out[22]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n230) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U34 ( .A1(SBOX_FF3_out[22]), .A2(
        SBOX_FF3_out[10]), .ZN(SBOX_Inst_f4_multd_H_himul_n229) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U33 ( .A(SBOX_Inst_f4_multd_H_himul_n227), .B(SBOX_Inst_f4_multd_H_himul_n226), .ZN(SBOX_Inst_f4_multd_H_himul_n228) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U32 ( .A1(
        SBOX_Inst_f4_multd_H_himul_n291), .A2(SBOX_FF3_out[19]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n227) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U31 ( .A(SBOX_Inst_f4_multd_H_himul_n225), .B(SBOX_Inst_f4_multd_H_himul_n219), .ZN(SBOX_Inst_f4_multd_H_himul_n226) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U30 ( .A(SBOX_Inst_f4_multd_H_himul_n224), .B(SBOX_Inst_f4_multd_H_himul_n221), .ZN(SBOX_Inst_f4_multd_H_himul_n225) );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U29 ( .A1(SBOX_Inst_f4_multd_H_himul_n223), .A2(SBOX_Inst_f4_multd_H_himul_n222), .ZN(SBOX_Inst_f4_multd_H_himul_n224)
         );
  OAI22_X1 SBOX_Inst_f4_multd_H_himul_U28 ( .A1(SBOX_FF3_out[11]), .A2(
        SBOX_FF3_out[7]), .B1(SBOX_Inst_f4_multd_H_himul_n290), .B2(
        SBOX_Inst_f4_multd_H_himul_n299), .ZN(SBOX_Inst_f4_multd_H_himul_n223)
         );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U27 ( .A(SBOX_FF3_out[18]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n222) );
  OAI211_X1 SBOX_Inst_f4_multd_H_himul_U26 ( .C1(SBOX_FF3_out[18]), .C2(
        SBOX_FF3_out[23]), .A(SBOX_FF3_out[6]), .B(
        SBOX_Inst_f4_multd_H_himul_n220), .ZN(SBOX_Inst_f4_multd_H_himul_n221)
         );
  OR2_X1 SBOX_Inst_f4_multd_H_himul_U25 ( .A1(SBOX_Inst_f4_multd_H_himul_n279), 
        .A2(SBOX_Inst_f4_multd_H_himul_n306), .ZN(
        SBOX_Inst_f4_multd_H_himul_n220) );
  OAI211_X1 SBOX_Inst_f4_multd_H_himul_U24 ( .C1(
        SBOX_Inst_f4_multd_H_himul_n217), .C2(SBOX_FF3_out[22]), .A(
        SBOX_FF3_out[7]), .B(SBOX_Inst_f4_multd_H_himul_n218), .ZN(
        SBOX_Inst_f4_multd_H_himul_n219) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U23 ( .A1(
        SBOX_Inst_f4_multd_H_himul_n217), .A2(SBOX_FF3_out[22]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n218) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U22 ( .A1(SBOX_FF3_out[19]), .A2(
        SBOX_FF3_out[23]), .B1(SBOX_Inst_f4_multd_H_himul_n279), .B2(
        SBOX_Inst_f4_multd_H_himul_n300), .ZN(SBOX_Inst_f4_multd_H_himul_n217)
         );
  XOR2_X1 SBOX_Inst_f4_multd_H_himul_U21 ( .A(SBOX_Inst_f4_multd_H_himul_n215), 
        .B(SBOX_Inst_f4_multd_H_himul_n216), .Z(
        SBOX_Inst_f4_multd_H_himul_n297) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U20 ( .A1(SBOX_FF3_out[15]), .A2(
        SBOX_FF3_out[2]), .ZN(SBOX_Inst_f4_multd_H_himul_n216) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U19 ( .A1(SBOX_FF3_out[3]), .A2(
        SBOX_FF3_out[14]), .ZN(SBOX_Inst_f4_multd_H_himul_n215) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U18 ( .A1(SBOX_FF3_out[23]), .A2(
        SBOX_FF3_out[15]), .B1(SBOX_Inst_f4_multd_H_himul_n303), .B2(
        SBOX_Inst_f4_multd_H_himul_n279), .ZN(SBOX_Inst_f4_multd_H_himul_n280)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_himul_U17 ( .A(SBOX_Inst_f4_multd_H_himul_n297), .B(SBOX_Inst_f4_multd_H_himul_n289), .ZN(SBOX_Inst_f4_multd_H_himul_n288) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U16 ( .A(SBOX_FF3_out[3]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n302) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U15 ( .A(SBOX_FF3_out[6]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n308) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U14 ( .A1(SBOX_FF3_out[2]), .A2(
        SBOX_FF3_out[19]), .ZN(SBOX_Inst_f4_multd_H_himul_n293) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U13 ( .A1(SBOX_FF3_out[3]), .A2(
        SBOX_FF3_out[18]), .ZN(SBOX_Inst_f4_multd_H_himul_n294) );
  NAND2_X1 SBOX_Inst_f4_multd_H_himul_U12 ( .A1(
        SBOX_Inst_f4_multd_H_himul_n305), .A2(SBOX_FF3_out[15]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n296) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U11 ( .A(SBOX_FF3_out[7]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n299) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U10 ( .A(SBOX_FF3_out[14]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n304) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U9 ( .A(SBOX_FF3_out[19]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n300) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U8 ( .A(SBOX_FF3_out[18]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n306) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U7 ( .A(SBOX_FF3_out[2]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n307) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U6 ( .A(SBOX_FF3_out[15]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n303) );
  AOI22_X1 SBOX_Inst_f4_multd_H_himul_U5 ( .A1(SBOX_FF3_out[19]), .A2(
        SBOX_Inst_f4_multd_H_himul_n306), .B1(SBOX_FF3_out[18]), .B2(
        SBOX_Inst_f4_multd_H_himul_n300), .ZN(SBOX_Inst_f4_multd_H_himul_n298)
         );
  NOR2_X1 SBOX_Inst_f4_multd_H_himul_U4 ( .A1(SBOX_Inst_f4_multd_H_himul_n275), 
        .A2(SBOX_Inst_f4_multd_H_himul_n279), .ZN(
        SBOX_Inst_f4_multd_H_himul_n292) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U3 ( .A(SBOX_FF3_out[23]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n279) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U2 ( .A(SBOX_FF3_out[22]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n278) );
  INV_X1 SBOX_Inst_f4_multd_H_himul_U1 ( .A(SBOX_FF3_out[10]), .ZN(
        SBOX_Inst_f4_multd_H_himul_n275) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U8 ( .A(PRNGQ[30]), .B(
        SBOX_Inst_f4_multd_H_Orig_ph[2]), .Z(SBOX_ph_H[2]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U7 ( .A(PRNGQ[29]), .B(
        SBOX_Inst_f4_multd_H_Orig_ph[1]), .Z(SBOX_ph_H[1]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U6 ( .A(
        SBOX_Inst_f4_multd_H_AddNewMaskph_n6), .B(PRNGQ[31]), .ZN(SBOX_ph_H[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U5 ( .A(PRNGQ[29]), .B(
        SBOX_Inst_f4_multd_H_Orig_ph[5]), .ZN(
        SBOX_Inst_f4_multd_H_AddNewMaskph_n6) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U4 ( .A(
        SBOX_Inst_f4_multd_H_AddNewMaskph_n5), .B(PRNGQ[30]), .ZN(SBOX_ph_H[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U3 ( .A(PRNGQ[28]), .B(
        SBOX_Inst_f4_multd_H_Orig_ph[4]), .ZN(
        SBOX_Inst_f4_multd_H_AddNewMaskph_n5) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U2 ( .A(PRNGQ[31]), .B(
        SBOX_Inst_f4_multd_H_Orig_ph[3]), .Z(SBOX_ph_H[3]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskph_U1 ( .A(PRNGQ[28]), .B(
        SBOX_Inst_f4_multd_H_Orig_ph[0]), .Z(SBOX_ph_H[0]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U100 ( .A(
        SBOX_Inst_f4_multd_H_summul_n296), .B(SBOX_Inst_f4_multd_H_summul_n295), .ZN(SBOX_Inst_f4_multd_H_summul_n301) );
  XOR2_X1 SBOX_Inst_f4_multd_H_summul_U99 ( .A(
        SBOX_Inst_f4_multd_H_summul_n294), .B(SBOX_Inst_f4_multd_H_summul_n293), .Z(SBOX_Inst_f4_multd_H_summul_n295) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U98 ( .A1(SBOX_Inst_f4_multd_H_sA[0]), 
        .A2(SBOX_Inst_f4_multd_H_sB[3]), .ZN(SBOX_Inst_f4_multd_H_summul_n293)
         );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U97 ( .A1(SBOX_Inst_f4_multd_H_sA[1]), 
        .A2(SBOX_Inst_f4_multd_H_sB[2]), .ZN(SBOX_Inst_f4_multd_H_summul_n294)
         );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U96 ( .A1(SBOX_Inst_f4_multd_H_sA[2]), 
        .A2(SBOX_Inst_f4_multd_H_sA[0]), .B1(SBOX_Inst_f4_multd_H_summul_n307), 
        .B2(SBOX_Inst_f4_multd_H_summul_n308), .ZN(
        SBOX_Inst_f4_multd_H_summul_n305) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U95 ( .A(
        SBOX_Inst_f4_multd_H_summul_n288), .B(SBOX_Inst_f4_multd_H_summul_n287), .ZN(SBOX_Inst_f4_multd_H_Orig_p[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U94 ( .A(
        SBOX_Inst_f4_multd_H_summul_n286), .B(SBOX_Inst_f4_multd_H_summul_n285), .ZN(SBOX_Inst_f4_multd_H_summul_n287) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U93 ( .A1(SBOX_Inst_f4_multd_H_sA[0]), 
        .A2(SBOX_Inst_f4_multd_H_sB[5]), .ZN(SBOX_Inst_f4_multd_H_summul_n285)
         );
  XOR2_X1 SBOX_Inst_f4_multd_H_summul_U92 ( .A(
        SBOX_Inst_f4_multd_H_summul_n284), .B(SBOX_Inst_f4_multd_H_summul_n283), .Z(SBOX_Inst_f4_multd_H_summul_n286) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U91 ( .A(
        SBOX_Inst_f4_multd_H_summul_n282), .B(SBOX_Inst_f4_multd_H_summul_n281), .ZN(SBOX_Inst_f4_multd_H_summul_n283) );
  MUX2_X1 SBOX_Inst_f4_multd_H_summul_U90 ( .A(SBOX_Inst_f4_multd_H_sB[4]), 
        .B(SBOX_Inst_f4_multd_H_summul_n280), .S(SBOX_Inst_f4_multd_H_sA[5]), 
        .Z(SBOX_Inst_f4_multd_H_summul_n281) );
  OAI221_X1 SBOX_Inst_f4_multd_H_summul_U89 ( .B1(SBOX_Inst_f4_multd_H_sB[5]), 
        .B2(SBOX_Inst_f4_multd_H_sB[4]), .C1(SBOX_Inst_f4_multd_H_summul_n279), 
        .C2(SBOX_Inst_f4_multd_H_summul_n278), .A(SBOX_Inst_f4_multd_H_sA[1]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n282) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U88 ( .A1(SBOX_Inst_f4_multd_H_sA[1]), 
        .A2(SBOX_Inst_f4_multd_H_sB[0]), .B1(SBOX_Inst_f4_multd_H_summul_n304), 
        .B2(SBOX_Inst_f4_multd_H_summul_n302), .ZN(
        SBOX_Inst_f4_multd_H_summul_n284) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U87 ( .A(SBOX_Inst_f4_multd_H_sA[1]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n302) );
  XOR2_X1 SBOX_Inst_f4_multd_H_summul_U86 ( .A(
        SBOX_Inst_f4_multd_H_summul_n277), .B(SBOX_Inst_f4_multd_H_summul_n276), .Z(SBOX_Inst_f4_multd_H_summul_n289) );
  XOR2_X1 SBOX_Inst_f4_multd_H_summul_U85 ( .A(
        SBOX_Inst_f4_multd_H_summul_n275), .B(SBOX_Inst_f4_multd_H_summul_n274), .Z(SBOX_Inst_f4_multd_H_summul_n297) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U84 ( .A1(SBOX_Inst_f4_multd_H_sA[4]), 
        .A2(SBOX_Inst_f4_multd_H_sA[5]), .B1(SBOX_Inst_f4_multd_H_summul_n290), 
        .B2(SBOX_Inst_f4_multd_H_summul_n273), .ZN(
        SBOX_Inst_f4_multd_H_summul_n291) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U83 ( .A(
        SBOX_Inst_f4_multd_H_summul_n271), .B(SBOX_Inst_f4_multd_H_summul_n272), .ZN(SBOX_Inst_f4_multd_H_Orig_p[5]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_summul_U82 ( .A(
        SBOX_Inst_f4_multd_H_summul_n267), .B(SBOX_Inst_f4_multd_H_summul_n269), .Z(SBOX_Inst_f4_multd_H_summul_n272) );
  AOI211_X1 SBOX_Inst_f4_multd_H_summul_U81 ( .C1(SBOX_Inst_f4_multd_H_sB[0]), 
        .C2(SBOX_Inst_f4_multd_H_sB[3]), .A(SBOX_Inst_f4_multd_H_summul_n270), 
        .B(SBOX_Inst_f4_multd_H_summul_n299), .ZN(
        SBOX_Inst_f4_multd_H_summul_n271) );
  AND2_X1 SBOX_Inst_f4_multd_H_summul_U80 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n304), .A2(
        SBOX_Inst_f4_multd_H_summul_n300), .ZN(
        SBOX_Inst_f4_multd_H_summul_n270) );
  AOI211_X1 SBOX_Inst_f4_multd_H_summul_U79 ( .C1(SBOX_Inst_f4_multd_H_sA[0]), 
        .C2(SBOX_Inst_f4_multd_H_sA[2]), .A(SBOX_Inst_f4_multd_H_summul_n306), 
        .B(SBOX_Inst_f4_multd_H_summul_n268), .ZN(
        SBOX_Inst_f4_multd_H_summul_n269) );
  AND2_X1 SBOX_Inst_f4_multd_H_summul_U78 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n307), .A2(
        SBOX_Inst_f4_multd_H_summul_n308), .ZN(
        SBOX_Inst_f4_multd_H_summul_n268) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U77 ( .A(
        SBOX_Inst_f4_multd_H_summul_n265), .B(SBOX_Inst_f4_multd_H_summul_n266), .ZN(SBOX_Inst_f4_multd_H_summul_n267) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U76 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n303), .A2(
        SBOX_Inst_f4_multd_H_summul_n302), .ZN(
        SBOX_Inst_f4_multd_H_summul_n266) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U75 ( .A(
        SBOX_Inst_f4_multd_H_summul_n301), .B(SBOX_Inst_f4_multd_H_summul_n264), .ZN(SBOX_Inst_f4_multd_H_summul_n265) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U74 ( .A1(SBOX_Inst_f4_multd_H_sA[1]), 
        .A2(SBOX_Inst_f4_multd_H_summul_n304), .B1(SBOX_Inst_f4_multd_H_sB[0]), 
        .B2(SBOX_Inst_f4_multd_H_summul_n305), .ZN(
        SBOX_Inst_f4_multd_H_summul_n264) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U73 ( .A(
        SBOX_Inst_f4_multd_H_summul_n263), .B(SBOX_Inst_f4_multd_H_summul_n262), .ZN(SBOX_Inst_f4_multd_H_Orig_p[3]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U72 ( .A(
        SBOX_Inst_f4_multd_H_summul_n258), .B(SBOX_Inst_f4_multd_H_summul_n260), .ZN(SBOX_Inst_f4_multd_H_summul_n263) );
  OAI221_X1 SBOX_Inst_f4_multd_H_summul_U71 ( .B1(
        SBOX_Inst_f4_multd_H_summul_n252), .B2(SBOX_Inst_f4_multd_H_sA[1]), 
        .C1(SBOX_Inst_f4_multd_H_summul_n261), .C2(
        SBOX_Inst_f4_multd_H_summul_n302), .A(SBOX_Inst_f4_multd_H_sB[4]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n262) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U70 ( .A(SBOX_Inst_f4_multd_H_summul_n252), .ZN(SBOX_Inst_f4_multd_H_summul_n261) );
  OAI21_X1 SBOX_Inst_f4_multd_H_summul_U69 ( .B1(
        SBOX_Inst_f4_multd_H_summul_n292), .B2(
        SBOX_Inst_f4_multd_H_summul_n291), .A(SBOX_Inst_f4_multd_H_summul_n259), .ZN(SBOX_Inst_f4_multd_H_summul_n260) );
  NAND3_X1 SBOX_Inst_f4_multd_H_summul_U68 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n292), .A2(SBOX_Inst_f4_multd_H_sA[4]), 
        .A3(SBOX_Inst_f4_multd_H_summul_n290), .ZN(
        SBOX_Inst_f4_multd_H_summul_n259) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U67 ( .A(
        SBOX_Inst_f4_multd_H_summul_n256), .B(SBOX_Inst_f4_multd_H_summul_n257), .ZN(SBOX_Inst_f4_multd_H_summul_n258) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U66 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n252), .A2(SBOX_Inst_f4_multd_H_sB[5]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n257) );
  XOR2_X1 SBOX_Inst_f4_multd_H_summul_U65 ( .A(
        SBOX_Inst_f4_multd_H_summul_n289), .B(SBOX_Inst_f4_multd_H_summul_n255), .Z(SBOX_Inst_f4_multd_H_summul_n256) );
  XOR2_X1 SBOX_Inst_f4_multd_H_summul_U64 ( .A(
        SBOX_Inst_f4_multd_H_summul_n253), .B(SBOX_Inst_f4_multd_H_summul_n254), .Z(SBOX_Inst_f4_multd_H_summul_n255) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U63 ( .A1(SBOX_Inst_f4_multd_H_sB[0]), 
        .A2(SBOX_Inst_f4_multd_H_sA[4]), .ZN(SBOX_Inst_f4_multd_H_summul_n254)
         );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U62 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n303), .A2(SBOX_Inst_f4_multd_H_sA[1]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n253) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U61 ( .A1(SBOX_Inst_f4_multd_H_sA[5]), 
        .A2(SBOX_Inst_f4_multd_H_sA[0]), .B1(SBOX_Inst_f4_multd_H_summul_n290), 
        .B2(SBOX_Inst_f4_multd_H_summul_n307), .ZN(
        SBOX_Inst_f4_multd_H_summul_n252) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U60 ( .A(
        SBOX_Inst_f4_multd_H_summul_n251), .B(SBOX_Inst_f4_multd_H_summul_n250), .ZN(SBOX_Inst_f4_multd_H_Orig_p[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U59 ( .A(
        SBOX_Inst_f4_multd_H_summul_n297), .B(SBOX_Inst_f4_multd_H_summul_n247), .ZN(SBOX_Inst_f4_multd_H_summul_n251) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U58 ( .A(
        SBOX_Inst_f4_multd_H_summul_n248), .B(SBOX_Inst_f4_multd_H_summul_n249), .ZN(SBOX_Inst_f4_multd_H_summul_n250) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U57 ( .A1(SBOX_Inst_f4_multd_H_sB[3]), 
        .A2(SBOX_Inst_f4_multd_H_summul_n302), .ZN(
        SBOX_Inst_f4_multd_H_summul_n249) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U56 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n308), .A2(
        SBOX_Inst_f4_multd_H_summul_n298), .ZN(
        SBOX_Inst_f4_multd_H_summul_n248) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U55 ( .A(
        SBOX_Inst_f4_multd_H_summul_n301), .B(SBOX_Inst_f4_multd_H_summul_n246), .ZN(SBOX_Inst_f4_multd_H_summul_n247) );
  MUX2_X1 SBOX_Inst_f4_multd_H_summul_U54 ( .A(SBOX_Inst_f4_multd_H_sB[0]), 
        .B(SBOX_Inst_f4_multd_H_sB[1]), .S(SBOX_Inst_f4_multd_H_summul_n245), 
        .Z(SBOX_Inst_f4_multd_H_summul_n246) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U53 ( .A1(SBOX_Inst_f4_multd_H_sA[3]), 
        .A2(SBOX_Inst_f4_multd_H_sA[1]), .B1(SBOX_Inst_f4_multd_H_summul_n302), 
        .B2(SBOX_Inst_f4_multd_H_summul_n299), .ZN(
        SBOX_Inst_f4_multd_H_summul_n245) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U52 ( .A(
        SBOX_Inst_f4_multd_H_summul_n242), .B(SBOX_Inst_f4_multd_H_summul_n244), .ZN(SBOX_Inst_f4_multd_H_Orig_p[1]) );
  AOI211_X1 SBOX_Inst_f4_multd_H_summul_U51 ( .C1(SBOX_Inst_f4_multd_H_sA[4]), 
        .C2(SBOX_Inst_f4_multd_H_sA[2]), .A(SBOX_Inst_f4_multd_H_summul_n298), 
        .B(SBOX_Inst_f4_multd_H_summul_n243), .ZN(
        SBOX_Inst_f4_multd_H_summul_n244) );
  AND2_X1 SBOX_Inst_f4_multd_H_summul_U50 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n273), .A2(
        SBOX_Inst_f4_multd_H_summul_n308), .ZN(
        SBOX_Inst_f4_multd_H_summul_n243) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U49 ( .A(
        SBOX_Inst_f4_multd_H_summul_n241), .B(SBOX_Inst_f4_multd_H_summul_n238), .ZN(SBOX_Inst_f4_multd_H_summul_n242) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U48 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n240), .A2(
        SBOX_Inst_f4_multd_H_summul_n239), .ZN(
        SBOX_Inst_f4_multd_H_summul_n241) );
  OAI22_X1 SBOX_Inst_f4_multd_H_summul_U47 ( .A1(SBOX_Inst_f4_multd_H_sA[3]), 
        .A2(SBOX_Inst_f4_multd_H_sA[4]), .B1(SBOX_Inst_f4_multd_H_summul_n273), 
        .B2(SBOX_Inst_f4_multd_H_summul_n299), .ZN(
        SBOX_Inst_f4_multd_H_summul_n240) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U46 ( .A(SBOX_Inst_f4_multd_H_sB[4]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n239) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U45 ( .A(
        SBOX_Inst_f4_multd_H_summul_n236), .B(SBOX_Inst_f4_multd_H_summul_n237), .ZN(SBOX_Inst_f4_multd_H_summul_n238) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U44 ( .A(SBOX_Inst_f4_multd_H_sA[4]), 
        .B(SBOX_Inst_f4_multd_H_summul_n234), .ZN(
        SBOX_Inst_f4_multd_H_summul_n237) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U43 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n229), .A2(
        SBOX_Inst_f4_multd_H_summul_n235), .ZN(
        SBOX_Inst_f4_multd_H_summul_n236) );
  OAI22_X1 SBOX_Inst_f4_multd_H_summul_U42 ( .A1(SBOX_Inst_f4_multd_H_sB[2]), 
        .A2(SBOX_Inst_f4_multd_H_sB[3]), .B1(SBOX_Inst_f4_multd_H_summul_n306), 
        .B2(SBOX_Inst_f4_multd_H_summul_n300), .ZN(
        SBOX_Inst_f4_multd_H_summul_n235) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U41 ( .A(
        SBOX_Inst_f4_multd_H_summul_n233), .B(SBOX_Inst_f4_multd_H_summul_n232), .ZN(SBOX_Inst_f4_multd_H_summul_n234) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U40 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n230), .A2(
        SBOX_Inst_f4_multd_H_summul_n290), .ZN(
        SBOX_Inst_f4_multd_H_summul_n233) );
  OAI221_X1 SBOX_Inst_f4_multd_H_summul_U39 ( .B1(
        SBOX_Inst_f4_multd_H_summul_n230), .B2(SBOX_Inst_f4_multd_H_sB[4]), 
        .C1(SBOX_Inst_f4_multd_H_summul_n231), .C2(
        SBOX_Inst_f4_multd_H_summul_n278), .A(SBOX_Inst_f4_multd_H_sA[2]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n232) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U38 ( .A(SBOX_Inst_f4_multd_H_summul_n230), .ZN(SBOX_Inst_f4_multd_H_summul_n231) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U37 ( .A1(SBOX_Inst_f4_multd_H_sB[5]), 
        .A2(SBOX_Inst_f4_multd_H_sB[2]), .B1(SBOX_Inst_f4_multd_H_summul_n306), 
        .B2(SBOX_Inst_f4_multd_H_summul_n279), .ZN(
        SBOX_Inst_f4_multd_H_summul_n230) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U36 ( .A(SBOX_Inst_f4_multd_H_sA[3]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n229) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U35 ( .A(
        SBOX_Inst_f4_multd_H_summul_n226), .B(SBOX_Inst_f4_multd_H_summul_n228), .ZN(SBOX_Inst_f4_multd_H_Orig_p[0]) );
  OAI22_X1 SBOX_Inst_f4_multd_H_summul_U34 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n279), .A2(
        SBOX_Inst_f4_multd_H_summul_n227), .B1(
        SBOX_Inst_f4_multd_H_summul_n292), .B2(SBOX_Inst_f4_multd_H_sB[4]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n228) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U33 ( .A1(SBOX_Inst_f4_multd_H_sB[4]), 
        .A2(SBOX_Inst_f4_multd_H_sA[4]), .ZN(SBOX_Inst_f4_multd_H_summul_n227)
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U32 ( .A(
        SBOX_Inst_f4_multd_H_summul_n225), .B(SBOX_Inst_f4_multd_H_summul_n224), .ZN(SBOX_Inst_f4_multd_H_summul_n226) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U31 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n291), .A2(SBOX_Inst_f4_multd_H_sB[3]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n225) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U30 ( .A(
        SBOX_Inst_f4_multd_H_summul_n223), .B(SBOX_Inst_f4_multd_H_summul_n217), .ZN(SBOX_Inst_f4_multd_H_summul_n224) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U29 ( .A(
        SBOX_Inst_f4_multd_H_summul_n222), .B(SBOX_Inst_f4_multd_H_summul_n219), .ZN(SBOX_Inst_f4_multd_H_summul_n223) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U28 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n221), .A2(
        SBOX_Inst_f4_multd_H_summul_n220), .ZN(
        SBOX_Inst_f4_multd_H_summul_n222) );
  OAI22_X1 SBOX_Inst_f4_multd_H_summul_U27 ( .A1(SBOX_Inst_f4_multd_H_sA[5]), 
        .A2(SBOX_Inst_f4_multd_H_sA[3]), .B1(SBOX_Inst_f4_multd_H_summul_n290), 
        .B2(SBOX_Inst_f4_multd_H_summul_n299), .ZN(
        SBOX_Inst_f4_multd_H_summul_n221) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U26 ( .A(SBOX_Inst_f4_multd_H_sB[2]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n220) );
  OAI211_X1 SBOX_Inst_f4_multd_H_summul_U25 ( .C1(SBOX_Inst_f4_multd_H_sB[2]), 
        .C2(SBOX_Inst_f4_multd_H_sB[5]), .A(SBOX_Inst_f4_multd_H_sA[2]), .B(
        SBOX_Inst_f4_multd_H_summul_n218), .ZN(
        SBOX_Inst_f4_multd_H_summul_n219) );
  OR2_X1 SBOX_Inst_f4_multd_H_summul_U24 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n279), .A2(
        SBOX_Inst_f4_multd_H_summul_n306), .ZN(
        SBOX_Inst_f4_multd_H_summul_n218) );
  OAI211_X1 SBOX_Inst_f4_multd_H_summul_U23 ( .C1(
        SBOX_Inst_f4_multd_H_summul_n215), .C2(SBOX_Inst_f4_multd_H_sB[4]), 
        .A(SBOX_Inst_f4_multd_H_sA[3]), .B(SBOX_Inst_f4_multd_H_summul_n216), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n217) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U22 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n215), .A2(SBOX_Inst_f4_multd_H_sB[4]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n216) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U21 ( .A1(SBOX_Inst_f4_multd_H_sB[3]), 
        .A2(SBOX_Inst_f4_multd_H_sB[5]), .B1(SBOX_Inst_f4_multd_H_summul_n279), 
        .B2(SBOX_Inst_f4_multd_H_summul_n300), .ZN(
        SBOX_Inst_f4_multd_H_summul_n215) );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U20 ( .A1(SBOX_Inst_f4_multd_H_sB[5]), 
        .A2(SBOX_Inst_f4_multd_H_sB[1]), .B1(SBOX_Inst_f4_multd_H_summul_n303), 
        .B2(SBOX_Inst_f4_multd_H_summul_n279), .ZN(
        SBOX_Inst_f4_multd_H_summul_n280) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_summul_U19 ( .A(
        SBOX_Inst_f4_multd_H_summul_n297), .B(SBOX_Inst_f4_multd_H_summul_n289), .ZN(SBOX_Inst_f4_multd_H_summul_n288) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U18 ( .A(SBOX_Inst_f4_multd_H_sA[2]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n308) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U17 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n305), .A2(SBOX_Inst_f4_multd_H_sB[1]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n296) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U16 ( .A(SBOX_Inst_f4_multd_H_sA[3]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n299) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U15 ( .A(SBOX_Inst_f4_multd_H_sB[0]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n304) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U14 ( .A(SBOX_Inst_f4_multd_H_sB[3]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n300) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U13 ( .A(SBOX_Inst_f4_multd_H_sB[2]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n306) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U12 ( .A(SBOX_Inst_f4_multd_H_sA[0]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n307) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U11 ( .A(SBOX_Inst_f4_multd_H_sB[1]), 
        .ZN(SBOX_Inst_f4_multd_H_summul_n303) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U10 ( .A1(SBOX_Inst_f4_multd_H_sB[1]), 
        .A2(SBOX_Inst_f4_multd_H_sA[0]), .ZN(SBOX_Inst_f4_multd_H_summul_n274)
         );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U9 ( .A1(SBOX_Inst_f4_multd_H_sA[1]), 
        .A2(SBOX_Inst_f4_multd_H_sB[0]), .ZN(SBOX_Inst_f4_multd_H_summul_n275)
         );
  AOI22_X1 SBOX_Inst_f4_multd_H_summul_U8 ( .A1(SBOX_Inst_f4_multd_H_sB[3]), 
        .A2(SBOX_Inst_f4_multd_H_summul_n306), .B1(SBOX_Inst_f4_multd_H_sB[2]), 
        .B2(SBOX_Inst_f4_multd_H_summul_n300), .ZN(
        SBOX_Inst_f4_multd_H_summul_n298) );
  NOR2_X1 SBOX_Inst_f4_multd_H_summul_U7 ( .A1(
        SBOX_Inst_f4_multd_H_summul_n273), .A2(
        SBOX_Inst_f4_multd_H_summul_n279), .ZN(
        SBOX_Inst_f4_multd_H_summul_n292) );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U6 ( .A1(SBOX_Inst_f4_multd_H_sB[1]), 
        .A2(SBOX_Inst_f4_multd_H_sA[4]), .ZN(SBOX_Inst_f4_multd_H_summul_n276)
         );
  NAND2_X1 SBOX_Inst_f4_multd_H_summul_U5 ( .A1(SBOX_Inst_f4_multd_H_sB[0]), 
        .A2(SBOX_Inst_f4_multd_H_sA[5]), .ZN(SBOX_Inst_f4_multd_H_summul_n277)
         );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U4 ( .A(SBOX_Inst_f4_multd_H_sA[5]), .ZN(
        SBOX_Inst_f4_multd_H_summul_n290) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U3 ( .A(SBOX_Inst_f4_multd_H_sB[5]), .ZN(
        SBOX_Inst_f4_multd_H_summul_n279) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U2 ( .A(SBOX_Inst_f4_multd_H_sB[4]), .ZN(
        SBOX_Inst_f4_multd_H_summul_n278) );
  INV_X1 SBOX_Inst_f4_multd_H_summul_U1 ( .A(SBOX_Inst_f4_multd_H_sA[4]), .ZN(
        SBOX_Inst_f4_multd_H_summul_n273) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U8 ( .A(PRNGQ[34]), .B(
        SBOX_Inst_f4_multd_H_Orig_p[2]), .Z(SBOX_p_H[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U7 ( .A(
        SBOX_Inst_f4_multd_H_AddNewMaskp_n6), .B(PRNGQ[35]), .ZN(SBOX_p_H[5])
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U6 ( .A(PRNGQ[33]), .B(
        SBOX_Inst_f4_multd_H_Orig_p[5]), .ZN(
        SBOX_Inst_f4_multd_H_AddNewMaskp_n6) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U5 ( .A(PRNGQ[35]), .B(
        SBOX_Inst_f4_multd_H_Orig_p[3]), .Z(SBOX_p_H[3]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U4 ( .A(
        SBOX_Inst_f4_multd_H_AddNewMaskp_n5), .B(PRNGQ[34]), .ZN(SBOX_p_H[4])
         );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U3 ( .A(PRNGQ[32]), .B(
        SBOX_Inst_f4_multd_H_Orig_p[4]), .ZN(
        SBOX_Inst_f4_multd_H_AddNewMaskp_n5) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U2 ( .A(PRNGQ[33]), .B(
        SBOX_Inst_f4_multd_H_Orig_p[1]), .Z(SBOX_p_H[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskp_U1 ( .A(PRNGQ[32]), .B(
        SBOX_Inst_f4_multd_H_Orig_p[0]), .Z(SBOX_p_H[0]) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U100 ( .A1(SBOX_FF3_out[4]), .A2(
        SBOX_FF3_out[0]), .B1(SBOX_Inst_f4_multd_H_lowmul_n307), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n308), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n305) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U99 ( .A(SBOX_FF3_out[0]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n307) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U98 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n292), .B(SBOX_Inst_f4_multd_H_lowmul_n291), .ZN(SBOX_Inst_f4_multd_H_Orig_pl[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U97 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n290), .B(SBOX_Inst_f4_multd_H_lowmul_n289), .ZN(SBOX_Inst_f4_multd_H_lowmul_n291) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U96 ( .A1(SBOX_FF3_out[0]), .A2(
        SBOX_FF3_out[21]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n289) );
  XOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U95 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n288), .B(SBOX_Inst_f4_multd_H_lowmul_n287), .Z(SBOX_Inst_f4_multd_H_lowmul_n290) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U94 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n286), .B(SBOX_Inst_f4_multd_H_lowmul_n285), .ZN(SBOX_Inst_f4_multd_H_lowmul_n287) );
  MUX2_X1 SBOX_Inst_f4_multd_H_lowmul_U93 ( .A(SBOX_FF3_out[20]), .B(
        SBOX_Inst_f4_multd_H_lowmul_n284), .S(SBOX_FF3_out[9]), .Z(
        SBOX_Inst_f4_multd_H_lowmul_n285) );
  OAI221_X1 SBOX_Inst_f4_multd_H_lowmul_U92 ( .B1(SBOX_FF3_out[21]), .B2(
        SBOX_FF3_out[20]), .C1(SBOX_Inst_f4_multd_H_lowmul_n283), .C2(
        SBOX_Inst_f4_multd_H_lowmul_n282), .A(SBOX_FF3_out[1]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n286) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U91 ( .A1(SBOX_FF3_out[1]), .A2(
        SBOX_FF3_out[12]), .B1(SBOX_Inst_f4_multd_H_lowmul_n304), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n302), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n288) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U90 ( .A(SBOX_FF3_out[1]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n302) );
  XOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U89 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n281), .B(SBOX_Inst_f4_multd_H_lowmul_n280), .Z(SBOX_Inst_f4_multd_H_lowmul_n297) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U88 ( .A1(SBOX_FF3_out[13]), .A2(
        SBOX_FF3_out[0]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n280) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U87 ( .A1(SBOX_FF3_out[1]), .A2(
        SBOX_FF3_out[12]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n281) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U86 ( .A(SBOX_FF3_out[4]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n308) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U85 ( .A1(SBOX_FF3_out[8]), .A2(
        SBOX_FF3_out[9]), .B1(SBOX_Inst_f4_multd_H_lowmul_n294), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n279), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n295) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U84 ( .A(SBOX_FF3_out[8]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n279) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U83 ( .A(SBOX_FF3_out[9]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n294) );
  XOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U82 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n277), .B(SBOX_Inst_f4_multd_H_lowmul_n278), .Z(SBOX_Inst_f4_multd_H_lowmul_n293) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U81 ( .A1(SBOX_FF3_out[13]), .A2(
        SBOX_FF3_out[8]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n278) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U80 ( .A1(SBOX_FF3_out[12]), .A2(
        SBOX_FF3_out[9]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n277) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U79 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n275), .B(SBOX_Inst_f4_multd_H_lowmul_n276), .ZN(SBOX_Inst_f4_multd_H_Orig_pl[5]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U78 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n271), .B(SBOX_Inst_f4_multd_H_lowmul_n273), .Z(SBOX_Inst_f4_multd_H_lowmul_n276) );
  AOI211_X1 SBOX_Inst_f4_multd_H_lowmul_U77 ( .C1(SBOX_FF3_out[12]), .C2(
        SBOX_FF3_out[17]), .A(SBOX_Inst_f4_multd_H_lowmul_n274), .B(
        SBOX_Inst_f4_multd_H_lowmul_n299), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n275) );
  AND2_X1 SBOX_Inst_f4_multd_H_lowmul_U76 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n304), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n300), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n274) );
  AOI211_X1 SBOX_Inst_f4_multd_H_lowmul_U75 ( .C1(SBOX_FF3_out[0]), .C2(
        SBOX_FF3_out[4]), .A(SBOX_Inst_f4_multd_H_lowmul_n306), .B(
        SBOX_Inst_f4_multd_H_lowmul_n272), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n273) );
  AND2_X1 SBOX_Inst_f4_multd_H_lowmul_U74 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n307), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n308), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n272) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U73 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n269), .B(SBOX_Inst_f4_multd_H_lowmul_n270), .ZN(SBOX_Inst_f4_multd_H_lowmul_n271) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U72 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n303), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n302), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n270) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U71 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n301), .B(SBOX_Inst_f4_multd_H_lowmul_n268), .ZN(SBOX_Inst_f4_multd_H_lowmul_n269) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U70 ( .A1(SBOX_FF3_out[1]), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n304), .B1(SBOX_FF3_out[12]), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n305), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n268) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U69 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n267), .B(SBOX_Inst_f4_multd_H_lowmul_n266), .ZN(SBOX_Inst_f4_multd_H_Orig_pl[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U68 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n297), .B(SBOX_Inst_f4_multd_H_lowmul_n263), .ZN(SBOX_Inst_f4_multd_H_lowmul_n267) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U67 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n264), .B(SBOX_Inst_f4_multd_H_lowmul_n265), .ZN(SBOX_Inst_f4_multd_H_lowmul_n266) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U66 ( .A1(SBOX_FF3_out[17]), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n302), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n265) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U65 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n308), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n298), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n264) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U64 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n301), .B(SBOX_Inst_f4_multd_H_lowmul_n262), .ZN(SBOX_Inst_f4_multd_H_lowmul_n263) );
  MUX2_X1 SBOX_Inst_f4_multd_H_lowmul_U63 ( .A(SBOX_FF3_out[12]), .B(
        SBOX_FF3_out[13]), .S(SBOX_Inst_f4_multd_H_lowmul_n261), .Z(
        SBOX_Inst_f4_multd_H_lowmul_n262) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U62 ( .A1(SBOX_FF3_out[5]), .A2(
        SBOX_FF3_out[1]), .B1(SBOX_Inst_f4_multd_H_lowmul_n302), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n299), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n261) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U61 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n260), .B(SBOX_Inst_f4_multd_H_lowmul_n259), .ZN(SBOX_Inst_f4_multd_H_lowmul_n301) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U60 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n305), .A2(SBOX_FF3_out[13]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n260) );
  XOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U59 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n257), .B(SBOX_Inst_f4_multd_H_lowmul_n258), .Z(SBOX_Inst_f4_multd_H_lowmul_n259) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U58 ( .A1(SBOX_FF3_out[17]), .A2(
        SBOX_FF3_out[0]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n258) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U57 ( .A1(SBOX_FF3_out[1]), .A2(
        SBOX_FF3_out[16]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n257) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U56 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n256), .B(SBOX_Inst_f4_multd_H_lowmul_n255), .ZN(SBOX_Inst_f4_multd_H_Orig_pl[3]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U55 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n251), .B(SBOX_Inst_f4_multd_H_lowmul_n253), .ZN(SBOX_Inst_f4_multd_H_lowmul_n256) );
  OAI221_X1 SBOX_Inst_f4_multd_H_lowmul_U54 ( .B1(
        SBOX_Inst_f4_multd_H_lowmul_n245), .B2(SBOX_FF3_out[1]), .C1(
        SBOX_Inst_f4_multd_H_lowmul_n254), .C2(
        SBOX_Inst_f4_multd_H_lowmul_n302), .A(SBOX_FF3_out[20]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n255) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U53 ( .A(SBOX_Inst_f4_multd_H_lowmul_n245), .ZN(SBOX_Inst_f4_multd_H_lowmul_n254) );
  OAI21_X1 SBOX_Inst_f4_multd_H_lowmul_U52 ( .B1(
        SBOX_Inst_f4_multd_H_lowmul_n296), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n295), .A(SBOX_Inst_f4_multd_H_lowmul_n252), .ZN(SBOX_Inst_f4_multd_H_lowmul_n253) );
  NAND3_X1 SBOX_Inst_f4_multd_H_lowmul_U51 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n296), .A2(SBOX_FF3_out[8]), .A3(
        SBOX_Inst_f4_multd_H_lowmul_n294), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n252) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U50 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n249), .B(SBOX_Inst_f4_multd_H_lowmul_n250), .ZN(SBOX_Inst_f4_multd_H_lowmul_n251) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U49 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n245), .A2(SBOX_FF3_out[21]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n250) );
  XOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U48 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n293), .B(SBOX_Inst_f4_multd_H_lowmul_n248), .Z(SBOX_Inst_f4_multd_H_lowmul_n249) );
  XOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U47 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n246), .B(SBOX_Inst_f4_multd_H_lowmul_n247), .Z(SBOX_Inst_f4_multd_H_lowmul_n248) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U46 ( .A1(SBOX_FF3_out[12]), .A2(
        SBOX_FF3_out[8]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n247) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U45 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n303), .A2(SBOX_FF3_out[1]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n246) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U44 ( .A1(SBOX_FF3_out[9]), .A2(
        SBOX_FF3_out[0]), .B1(SBOX_Inst_f4_multd_H_lowmul_n294), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n307), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n245) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U43 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n242), .B(SBOX_Inst_f4_multd_H_lowmul_n244), .ZN(SBOX_Inst_f4_multd_H_Orig_pl[1]) );
  AOI211_X1 SBOX_Inst_f4_multd_H_lowmul_U42 ( .C1(SBOX_FF3_out[8]), .C2(
        SBOX_FF3_out[4]), .A(SBOX_Inst_f4_multd_H_lowmul_n298), .B(
        SBOX_Inst_f4_multd_H_lowmul_n243), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n244) );
  AND2_X1 SBOX_Inst_f4_multd_H_lowmul_U41 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n279), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n308), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n243) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U40 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n241), .B(SBOX_Inst_f4_multd_H_lowmul_n238), .ZN(SBOX_Inst_f4_multd_H_lowmul_n242) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U39 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n240), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n239), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n241) );
  OAI22_X1 SBOX_Inst_f4_multd_H_lowmul_U38 ( .A1(SBOX_FF3_out[5]), .A2(
        SBOX_FF3_out[8]), .B1(SBOX_Inst_f4_multd_H_lowmul_n279), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n299), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n240) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U37 ( .A(SBOX_FF3_out[20]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n239) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U36 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n236), .B(SBOX_Inst_f4_multd_H_lowmul_n237), .ZN(SBOX_Inst_f4_multd_H_lowmul_n238) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U35 ( .A(SBOX_FF3_out[8]), .B(
        SBOX_Inst_f4_multd_H_lowmul_n234), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n237) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U34 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n229), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n235), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n236) );
  OAI22_X1 SBOX_Inst_f4_multd_H_lowmul_U33 ( .A1(SBOX_FF3_out[16]), .A2(
        SBOX_FF3_out[17]), .B1(SBOX_Inst_f4_multd_H_lowmul_n306), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n300), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n235) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U32 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n233), .B(SBOX_Inst_f4_multd_H_lowmul_n232), .ZN(SBOX_Inst_f4_multd_H_lowmul_n234) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U31 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n230), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n294), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n233) );
  OAI221_X1 SBOX_Inst_f4_multd_H_lowmul_U30 ( .B1(
        SBOX_Inst_f4_multd_H_lowmul_n230), .B2(SBOX_FF3_out[20]), .C1(
        SBOX_Inst_f4_multd_H_lowmul_n231), .C2(
        SBOX_Inst_f4_multd_H_lowmul_n282), .A(SBOX_FF3_out[4]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n232) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U29 ( .A(SBOX_Inst_f4_multd_H_lowmul_n230), .ZN(SBOX_Inst_f4_multd_H_lowmul_n231) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U28 ( .A1(SBOX_FF3_out[21]), .A2(
        SBOX_FF3_out[16]), .B1(SBOX_Inst_f4_multd_H_lowmul_n306), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n283), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n230) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U27 ( .A(SBOX_FF3_out[5]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n229) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U26 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n226), .B(SBOX_Inst_f4_multd_H_lowmul_n228), .ZN(SBOX_Inst_f4_multd_H_Orig_pl[0]) );
  OAI22_X1 SBOX_Inst_f4_multd_H_lowmul_U25 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n283), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n227), .B1(
        SBOX_Inst_f4_multd_H_lowmul_n296), .B2(SBOX_FF3_out[20]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n228) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U24 ( .A1(SBOX_FF3_out[20]), .A2(
        SBOX_FF3_out[8]), .ZN(SBOX_Inst_f4_multd_H_lowmul_n227) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U23 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n225), .B(SBOX_Inst_f4_multd_H_lowmul_n224), .ZN(SBOX_Inst_f4_multd_H_lowmul_n226) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U22 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n295), .A2(SBOX_FF3_out[17]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n225) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U21 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n223), .B(SBOX_Inst_f4_multd_H_lowmul_n217), .ZN(SBOX_Inst_f4_multd_H_lowmul_n224) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U20 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n222), .B(SBOX_Inst_f4_multd_H_lowmul_n219), .ZN(SBOX_Inst_f4_multd_H_lowmul_n223) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U19 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n221), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n220), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n222) );
  OAI22_X1 SBOX_Inst_f4_multd_H_lowmul_U18 ( .A1(SBOX_FF3_out[9]), .A2(
        SBOX_FF3_out[5]), .B1(SBOX_Inst_f4_multd_H_lowmul_n294), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n299), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n221) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U17 ( .A(SBOX_FF3_out[16]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n220) );
  OAI211_X1 SBOX_Inst_f4_multd_H_lowmul_U16 ( .C1(SBOX_FF3_out[16]), .C2(
        SBOX_FF3_out[21]), .A(SBOX_FF3_out[4]), .B(
        SBOX_Inst_f4_multd_H_lowmul_n218), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n219) );
  OR2_X1 SBOX_Inst_f4_multd_H_lowmul_U15 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n283), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n306), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n218) );
  OAI211_X1 SBOX_Inst_f4_multd_H_lowmul_U14 ( .C1(
        SBOX_Inst_f4_multd_H_lowmul_n215), .C2(SBOX_FF3_out[20]), .A(
        SBOX_FF3_out[5]), .B(SBOX_Inst_f4_multd_H_lowmul_n216), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n217) );
  NAND2_X1 SBOX_Inst_f4_multd_H_lowmul_U13 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n215), .A2(SBOX_FF3_out[20]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n216) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U12 ( .A1(SBOX_FF3_out[17]), .A2(
        SBOX_FF3_out[21]), .B1(SBOX_Inst_f4_multd_H_lowmul_n283), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n300), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n215) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U11 ( .A1(SBOX_FF3_out[21]), .A2(
        SBOX_FF3_out[13]), .B1(SBOX_Inst_f4_multd_H_lowmul_n303), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n283), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n284) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U10 ( .A(
        SBOX_Inst_f4_multd_H_lowmul_n297), .B(SBOX_Inst_f4_multd_H_lowmul_n293), .ZN(SBOX_Inst_f4_multd_H_lowmul_n292) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U9 ( .A(SBOX_FF3_out[5]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n299) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U8 ( .A(SBOX_FF3_out[12]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n304) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U7 ( .A(SBOX_FF3_out[17]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n300) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U6 ( .A(SBOX_FF3_out[16]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n306) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U5 ( .A(SBOX_FF3_out[13]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n303) );
  AOI22_X1 SBOX_Inst_f4_multd_H_lowmul_U4 ( .A1(SBOX_FF3_out[17]), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n306), .B1(SBOX_FF3_out[16]), .B2(
        SBOX_Inst_f4_multd_H_lowmul_n300), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n298) );
  NOR2_X1 SBOX_Inst_f4_multd_H_lowmul_U3 ( .A1(
        SBOX_Inst_f4_multd_H_lowmul_n279), .A2(
        SBOX_Inst_f4_multd_H_lowmul_n283), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n296) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U2 ( .A(SBOX_FF3_out[21]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n283) );
  INV_X1 SBOX_Inst_f4_multd_H_lowmul_U1 ( .A(SBOX_FF3_out[20]), .ZN(
        SBOX_Inst_f4_multd_H_lowmul_n282) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U8 ( .A(PRNGQ[38]), .B(
        SBOX_Inst_f4_multd_H_Orig_pl[2]), .Z(SBOX_pl_H[2]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U7 ( .A(
        SBOX_Inst_f4_multd_H_AddNewMaskpl_n6), .B(PRNGQ[39]), .ZN(SBOX_pl_H[5]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U6 ( .A(PRNGQ[37]), .B(
        SBOX_Inst_f4_multd_H_Orig_pl[5]), .ZN(
        SBOX_Inst_f4_multd_H_AddNewMaskpl_n6) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U5 ( .A(
        SBOX_Inst_f4_multd_H_AddNewMaskpl_n5), .B(PRNGQ[38]), .ZN(SBOX_pl_H[4]) );
  XNOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U4 ( .A(PRNGQ[36]), .B(
        SBOX_Inst_f4_multd_H_Orig_pl[4]), .ZN(
        SBOX_Inst_f4_multd_H_AddNewMaskpl_n5) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U3 ( .A(PRNGQ[39]), .B(
        SBOX_Inst_f4_multd_H_Orig_pl[3]), .Z(SBOX_pl_H[3]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U2 ( .A(PRNGQ[37]), .B(
        SBOX_Inst_f4_multd_H_Orig_pl[1]), .Z(SBOX_pl_H[1]) );
  XOR2_X1 SBOX_Inst_f4_multd_H_AddNewMaskpl_U1 ( .A(PRNGQ[36]), .B(
        SBOX_Inst_f4_multd_H_Orig_pl[0]), .Z(SBOX_pl_H[0]) );
  OAI21_X1 SBOX_PL_4_U73 ( .B1(1'b1), .B2(SBOX_PL_4_n180), .A(SBOX_PL_4_n252), 
        .ZN(SBOX_PL_4_n144) );
  NAND2_X1 SBOX_PL_4_U72 ( .A1(1'b1), .A2(SBOX_pl_L[0]), .ZN(SBOX_PL_4_n252)
         );
  OAI21_X1 SBOX_PL_4_U71 ( .B1(1'b1), .B2(SBOX_PL_4_n179), .A(SBOX_PL_4_n251), 
        .ZN(SBOX_PL_4_n143) );
  NAND2_X1 SBOX_PL_4_U70 ( .A1(1'b1), .A2(SBOX_pl_L[1]), .ZN(SBOX_PL_4_n251)
         );
  OAI21_X1 SBOX_PL_4_U69 ( .B1(1'b1), .B2(SBOX_PL_4_n178), .A(SBOX_PL_4_n250), 
        .ZN(SBOX_PL_4_n142) );
  NAND2_X1 SBOX_PL_4_U68 ( .A1(1'b1), .A2(SBOX_pl_L[2]), .ZN(SBOX_PL_4_n250)
         );
  OAI21_X1 SBOX_PL_4_U67 ( .B1(1'b1), .B2(SBOX_PL_4_n174), .A(SBOX_PL_4_n249), 
        .ZN(SBOX_PL_4_n138) );
  NAND2_X1 SBOX_PL_4_U66 ( .A1(1'b1), .A2(SBOX_p_L[0]), .ZN(SBOX_PL_4_n249) );
  OAI21_X1 SBOX_PL_4_U65 ( .B1(1'b1), .B2(SBOX_PL_4_n173), .A(SBOX_PL_4_n248), 
        .ZN(SBOX_PL_4_n137) );
  NAND2_X1 SBOX_PL_4_U64 ( .A1(1'b1), .A2(SBOX_p_L[1]), .ZN(SBOX_PL_4_n248) );
  OAI21_X1 SBOX_PL_4_U63 ( .B1(1'b1), .B2(SBOX_PL_4_n172), .A(SBOX_PL_4_n247), 
        .ZN(SBOX_PL_4_n136) );
  NAND2_X1 SBOX_PL_4_U62 ( .A1(1'b1), .A2(SBOX_p_L[2]), .ZN(SBOX_PL_4_n247) );
  OAI21_X1 SBOX_PL_4_U61 ( .B1(1'b1), .B2(SBOX_PL_4_n170), .A(SBOX_PL_4_n246), 
        .ZN(SBOX_PL_4_n134) );
  NAND2_X1 SBOX_PL_4_U60 ( .A1(1'b1), .A2(SBOX_p_L[4]), .ZN(SBOX_PL_4_n246) );
  OAI21_X1 SBOX_PL_4_U59 ( .B1(1'b1), .B2(SBOX_PL_4_n169), .A(SBOX_PL_4_n245), 
        .ZN(SBOX_PL_4_n133) );
  NAND2_X1 SBOX_PL_4_U58 ( .A1(1'b1), .A2(SBOX_p_L[5]), .ZN(SBOX_PL_4_n245) );
  OAI21_X1 SBOX_PL_4_U57 ( .B1(1'b1), .B2(SBOX_PL_4_n168), .A(SBOX_PL_4_n244), 
        .ZN(SBOX_PL_4_n132) );
  NAND2_X1 SBOX_PL_4_U56 ( .A1(1'b1), .A2(SBOX_ph_L[0]), .ZN(SBOX_PL_4_n244)
         );
  OAI21_X1 SBOX_PL_4_U55 ( .B1(1'b1), .B2(SBOX_PL_4_n167), .A(SBOX_PL_4_n243), 
        .ZN(SBOX_PL_4_n131) );
  NAND2_X1 SBOX_PL_4_U54 ( .A1(1'b1), .A2(SBOX_ph_L[1]), .ZN(SBOX_PL_4_n243)
         );
  OAI21_X1 SBOX_PL_4_U53 ( .B1(1'b1), .B2(SBOX_PL_4_n160), .A(SBOX_PL_4_n242), 
        .ZN(SBOX_PL_4_n124) );
  NAND2_X1 SBOX_PL_4_U52 ( .A1(1'b1), .A2(SBOX_pl_H[2]), .ZN(SBOX_PL_4_n242)
         );
  OAI21_X1 SBOX_PL_4_U51 ( .B1(1'b1), .B2(SBOX_PL_4_n154), .A(SBOX_PL_4_n241), 
        .ZN(SBOX_PL_4_n118) );
  NAND2_X1 SBOX_PL_4_U50 ( .A1(1'b1), .A2(SBOX_p_H[2]), .ZN(SBOX_PL_4_n241) );
  OAI21_X1 SBOX_PL_4_U49 ( .B1(1'b1), .B2(SBOX_PL_4_n148), .A(SBOX_PL_4_n240), 
        .ZN(SBOX_PL_4_n112) );
  NAND2_X1 SBOX_PL_4_U48 ( .A1(1'b1), .A2(SBOX_ph_H[2]), .ZN(SBOX_PL_4_n240)
         );
  OAI21_X1 SBOX_PL_4_U47 ( .B1(1'b1), .B2(SBOX_PL_4_n149), .A(SBOX_PL_4_n239), 
        .ZN(SBOX_PL_4_n113) );
  NAND2_X1 SBOX_PL_4_U46 ( .A1(1'b1), .A2(SBOX_ph_H[1]), .ZN(SBOX_PL_4_n239)
         );
  OAI21_X1 SBOX_PL_4_U45 ( .B1(1'b1), .B2(SBOX_PL_4_n176), .A(SBOX_PL_4_n238), 
        .ZN(SBOX_PL_4_n140) );
  NAND2_X1 SBOX_PL_4_U44 ( .A1(1'b1), .A2(SBOX_pl_L[4]), .ZN(SBOX_PL_4_n238)
         );
  OAI21_X1 SBOX_PL_4_U43 ( .B1(1'b1), .B2(SBOX_PL_4_n145), .A(SBOX_PL_4_n237), 
        .ZN(SBOX_PL_4_n109) );
  NAND2_X1 SBOX_PL_4_U42 ( .A1(1'b1), .A2(SBOX_ph_H[5]), .ZN(SBOX_PL_4_n237)
         );
  OAI21_X1 SBOX_PL_4_U41 ( .B1(1'b1), .B2(SBOX_PL_4_n157), .A(SBOX_PL_4_n236), 
        .ZN(SBOX_PL_4_n121) );
  NAND2_X1 SBOX_PL_4_U40 ( .A1(1'b1), .A2(SBOX_pl_H[5]), .ZN(SBOX_PL_4_n236)
         );
  OAI21_X1 SBOX_PL_4_U39 ( .B1(1'b1), .B2(SBOX_PL_4_n146), .A(SBOX_PL_4_n235), 
        .ZN(SBOX_PL_4_n110) );
  NAND2_X1 SBOX_PL_4_U38 ( .A1(1'b1), .A2(SBOX_ph_H[4]), .ZN(SBOX_PL_4_n235)
         );
  OAI21_X1 SBOX_PL_4_U37 ( .B1(1'b1), .B2(SBOX_PL_4_n158), .A(SBOX_PL_4_n234), 
        .ZN(SBOX_PL_4_n122) );
  NAND2_X1 SBOX_PL_4_U36 ( .A1(1'b1), .A2(SBOX_pl_H[4]), .ZN(SBOX_PL_4_n234)
         );
  OAI21_X1 SBOX_PL_4_U35 ( .B1(1'b1), .B2(SBOX_PL_4_n147), .A(SBOX_PL_4_n233), 
        .ZN(SBOX_PL_4_n111) );
  NAND2_X1 SBOX_PL_4_U34 ( .A1(1'b1), .A2(SBOX_ph_H[3]), .ZN(SBOX_PL_4_n233)
         );
  OAI21_X1 SBOX_PL_4_U33 ( .B1(1'b1), .B2(SBOX_PL_4_n175), .A(SBOX_PL_4_n232), 
        .ZN(SBOX_PL_4_n139) );
  NAND2_X1 SBOX_PL_4_U32 ( .A1(1'b1), .A2(SBOX_pl_L[5]), .ZN(SBOX_PL_4_n232)
         );
  OAI21_X1 SBOX_PL_4_U31 ( .B1(1'b1), .B2(SBOX_PL_4_n150), .A(SBOX_PL_4_n231), 
        .ZN(SBOX_PL_4_n114) );
  NAND2_X1 SBOX_PL_4_U30 ( .A1(1'b1), .A2(SBOX_ph_H[0]), .ZN(SBOX_PL_4_n231)
         );
  OAI21_X1 SBOX_PL_4_U29 ( .B1(1'b1), .B2(SBOX_PL_4_n151), .A(SBOX_PL_4_n230), 
        .ZN(SBOX_PL_4_n115) );
  NAND2_X1 SBOX_PL_4_U28 ( .A1(1'b1), .A2(SBOX_p_H[5]), .ZN(SBOX_PL_4_n230) );
  OAI21_X1 SBOX_PL_4_U27 ( .B1(1'b1), .B2(SBOX_PL_4_n153), .A(SBOX_PL_4_n229), 
        .ZN(SBOX_PL_4_n117) );
  NAND2_X1 SBOX_PL_4_U26 ( .A1(1'b1), .A2(SBOX_p_H[3]), .ZN(SBOX_PL_4_n229) );
  OAI21_X1 SBOX_PL_4_U25 ( .B1(1'b1), .B2(SBOX_PL_4_n159), .A(SBOX_PL_4_n228), 
        .ZN(SBOX_PL_4_n123) );
  NAND2_X1 SBOX_PL_4_U24 ( .A1(1'b1), .A2(SBOX_pl_H[3]), .ZN(SBOX_PL_4_n228)
         );
  OAI21_X1 SBOX_PL_4_U23 ( .B1(1'b1), .B2(SBOX_PL_4_n163), .A(SBOX_PL_4_n227), 
        .ZN(SBOX_PL_4_n127) );
  NAND2_X1 SBOX_PL_4_U22 ( .A1(1'b1), .A2(SBOX_ph_L[5]), .ZN(SBOX_PL_4_n227)
         );
  OAI21_X1 SBOX_PL_4_U21 ( .B1(1'b1), .B2(SBOX_PL_4_n152), .A(SBOX_PL_4_n226), 
        .ZN(SBOX_PL_4_n116) );
  NAND2_X1 SBOX_PL_4_U20 ( .A1(1'b1), .A2(SBOX_p_H[4]), .ZN(SBOX_PL_4_n226) );
  OAI21_X1 SBOX_PL_4_U19 ( .B1(1'b1), .B2(SBOX_PL_4_n171), .A(SBOX_PL_4_n225), 
        .ZN(SBOX_PL_4_n135) );
  NAND2_X1 SBOX_PL_4_U18 ( .A1(1'b1), .A2(SBOX_p_L[3]), .ZN(SBOX_PL_4_n225) );
  OAI21_X1 SBOX_PL_4_U17 ( .B1(1'b1), .B2(SBOX_PL_4_n155), .A(SBOX_PL_4_n224), 
        .ZN(SBOX_PL_4_n119) );
  NAND2_X1 SBOX_PL_4_U16 ( .A1(1'b1), .A2(SBOX_p_H[1]), .ZN(SBOX_PL_4_n224) );
  OAI21_X1 SBOX_PL_4_U15 ( .B1(1'b1), .B2(SBOX_PL_4_n156), .A(SBOX_PL_4_n223), 
        .ZN(SBOX_PL_4_n120) );
  NAND2_X1 SBOX_PL_4_U14 ( .A1(1'b1), .A2(SBOX_p_H[0]), .ZN(SBOX_PL_4_n223) );
  OAI21_X1 SBOX_PL_4_U13 ( .B1(1'b1), .B2(SBOX_PL_4_n161), .A(SBOX_PL_4_n222), 
        .ZN(SBOX_PL_4_n125) );
  NAND2_X1 SBOX_PL_4_U12 ( .A1(1'b1), .A2(SBOX_pl_H[1]), .ZN(SBOX_PL_4_n222)
         );
  OAI21_X1 SBOX_PL_4_U11 ( .B1(1'b1), .B2(SBOX_PL_4_n164), .A(SBOX_PL_4_n221), 
        .ZN(SBOX_PL_4_n128) );
  NAND2_X1 SBOX_PL_4_U10 ( .A1(1'b1), .A2(SBOX_ph_L[4]), .ZN(SBOX_PL_4_n221)
         );
  OAI21_X1 SBOX_PL_4_U9 ( .B1(1'b1), .B2(SBOX_PL_4_n162), .A(SBOX_PL_4_n220), 
        .ZN(SBOX_PL_4_n126) );
  NAND2_X1 SBOX_PL_4_U8 ( .A1(1'b1), .A2(SBOX_pl_H[0]), .ZN(SBOX_PL_4_n220) );
  OAI21_X1 SBOX_PL_4_U7 ( .B1(1'b1), .B2(SBOX_PL_4_n165), .A(SBOX_PL_4_n219), 
        .ZN(SBOX_PL_4_n129) );
  NAND2_X1 SBOX_PL_4_U6 ( .A1(1'b1), .A2(SBOX_ph_L[3]), .ZN(SBOX_PL_4_n219) );
  OAI21_X1 SBOX_PL_4_U5 ( .B1(1'b1), .B2(SBOX_PL_4_n166), .A(SBOX_PL_4_n218), 
        .ZN(SBOX_PL_4_n130) );
  NAND2_X1 SBOX_PL_4_U4 ( .A1(1'b1), .A2(SBOX_ph_L[2]), .ZN(SBOX_PL_4_n218) );
  OAI21_X1 SBOX_PL_4_U3 ( .B1(1'b1), .B2(SBOX_PL_4_n177), .A(SBOX_PL_4_n217), 
        .ZN(SBOX_PL_4_n141) );
  NAND2_X1 SBOX_PL_4_U2 ( .A1(1'b1), .A2(SBOX_pl_L[3]), .ZN(SBOX_PL_4_n217) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_0_ ( .D(SBOX_PL_4_n144), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[0]), .QN(SBOX_PL_4_n180) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_1_ ( .D(SBOX_PL_4_n143), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[1]), .QN(SBOX_PL_4_n179) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_2_ ( .D(SBOX_PL_4_n142), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[2]), .QN(SBOX_PL_4_n178) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_3_ ( .D(SBOX_PL_4_n141), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[3]), .QN(SBOX_PL_4_n177) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_4_ ( .D(SBOX_PL_4_n140), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[4]), .QN(SBOX_PL_4_n176) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_5_ ( .D(SBOX_PL_4_n139), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[5]), .QN(SBOX_PL_4_n175) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_6_ ( .D(SBOX_PL_4_n138), .CK(ClkxCI), 
        .Q(SBOX_Inst_f5_plwillwin_pw2_1_), .QN(SBOX_PL_4_n174) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_7_ ( .D(SBOX_PL_4_n137), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[7]), .QN(SBOX_PL_4_n173) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_8_ ( .D(SBOX_PL_4_n136), .CK(ClkxCI), 
        .Q(SBOX_Inst_f5_plwillwin_pw2_3_), .QN(SBOX_PL_4_n172) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_9_ ( .D(SBOX_PL_4_n135), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[9]), .QN(SBOX_PL_4_n171) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_10_ ( .D(SBOX_PL_4_n134), .CK(ClkxCI), 
        .Q(SBOX_Inst_f5_plwillwin_pw2_5_), .QN(SBOX_PL_4_n170) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_11_ ( .D(SBOX_PL_4_n133), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[11]), .QN(SBOX_PL_4_n169) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_12_ ( .D(SBOX_PL_4_n132), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[12]), .QN(SBOX_PL_4_n168) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_13_ ( .D(SBOX_PL_4_n131), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[13]), .QN(SBOX_PL_4_n167) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_14_ ( .D(SBOX_PL_4_n130), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[14]), .QN(SBOX_PL_4_n166) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_15_ ( .D(SBOX_PL_4_n129), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[15]), .QN(SBOX_PL_4_n165) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_16_ ( .D(SBOX_PL_4_n128), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[16]), .QN(SBOX_PL_4_n164) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_17_ ( .D(SBOX_PL_4_n127), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[17]), .QN(SBOX_PL_4_n163) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_18_ ( .D(SBOX_PL_4_n126), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[18]), .QN(SBOX_PL_4_n162) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_19_ ( .D(SBOX_PL_4_n125), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[19]), .QN(SBOX_PL_4_n161) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_20_ ( .D(SBOX_PL_4_n124), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[20]), .QN(SBOX_PL_4_n160) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_21_ ( .D(SBOX_PL_4_n123), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[21]), .QN(SBOX_PL_4_n159) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_22_ ( .D(SBOX_PL_4_n122), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[22]), .QN(SBOX_PL_4_n158) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_23_ ( .D(SBOX_PL_4_n121), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[23]), .QN(SBOX_PL_4_n157) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_24_ ( .D(SBOX_PL_4_n120), .CK(ClkxCI), 
        .Q(SBOX_Inst_f5_phwillwin_pw2_1_), .QN(SBOX_PL_4_n156) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_25_ ( .D(SBOX_PL_4_n119), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[25]), .QN(SBOX_PL_4_n155) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_26_ ( .D(SBOX_PL_4_n118), .CK(ClkxCI), 
        .Q(SBOX_Inst_f5_phwillwin_pw2_3_), .QN(SBOX_PL_4_n154) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_27_ ( .D(SBOX_PL_4_n117), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[27]), .QN(SBOX_PL_4_n153) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_28_ ( .D(SBOX_PL_4_n116), .CK(ClkxCI), 
        .Q(SBOX_Inst_f5_phwillwin_pw2_5_), .QN(SBOX_PL_4_n152) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_29_ ( .D(SBOX_PL_4_n115), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[29]), .QN(SBOX_PL_4_n151) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_30_ ( .D(SBOX_PL_4_n114), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[30]), .QN(SBOX_PL_4_n150) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_31_ ( .D(SBOX_PL_4_n113), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[31]), .QN(SBOX_PL_4_n149) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_32_ ( .D(SBOX_PL_4_n112), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[32]), .QN(SBOX_PL_4_n148) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_33_ ( .D(SBOX_PL_4_n111), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[33]), .QN(SBOX_PL_4_n147) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_34_ ( .D(SBOX_PL_4_n110), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[34]), .QN(SBOX_PL_4_n146) );
  DFF_X1 SBOX_PL_4_s_current_state_reg_35_ ( .D(SBOX_PL_4_n109), .CK(ClkxCI), 
        .Q(SBOX_FF4_out[35]), .QN(SBOX_PL_4_n145) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U12 ( .A(SBOX_Inst_f5_phwillwin_pw2_5_), .B(
        SBOX_FF4_out[35]), .Z(SBOX_Inst_f5_ph[11]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U11 ( .A(SBOX_Inst_f5_phwillwin_pw2_1_), .B(
        SBOX_FF4_out[31]), .Z(SBOX_Inst_f5_ph[3]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U10 ( .A(SBOX_Inst_f5_phwillwin_pw2_3_), .B(
        SBOX_FF4_out[33]), .Z(SBOX_Inst_f5_ph[7]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U9 ( .A(SBOX_Inst_f5_phwillwin_pw2_5_), .B(
        SBOX_FF4_out[23]), .Z(SBOX_Inst_f5_ph[9]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U8 ( .A(SBOX_Inst_f5_phwillwin_pw2_4_), .B(
        SBOX_FF4_out[22]), .Z(SBOX_Inst_f5_ph[8]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U7 ( .A(SBOX_Inst_f5_phwillwin_pw2_3_), .B(
        SBOX_FF4_out[21]), .Z(SBOX_Inst_f5_ph[5]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U6 ( .A(SBOX_Inst_f5_phwillwin_pw2_2_), .B(
        SBOX_FF4_out[20]), .Z(SBOX_Inst_f5_ph[4]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U5 ( .A(SBOX_Inst_f5_phwillwin_pw2_1_), .B(
        SBOX_FF4_out[19]), .Z(SBOX_Inst_f5_ph[1]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U4 ( .A(SBOX_Inst_f5_phwillwin_pw2_0_), .B(
        SBOX_FF4_out[18]), .Z(SBOX_Inst_f5_ph[0]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U3 ( .A(SBOX_Inst_f5_phwillwin_pw2_4_), .B(
        SBOX_FF4_out[34]), .Z(SBOX_Inst_f5_ph[10]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U2 ( .A(SBOX_Inst_f5_phwillwin_pw2_2_), .B(
        SBOX_FF4_out[32]), .Z(SBOX_Inst_f5_ph[6]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_U1 ( .A(SBOX_Inst_f5_phwillwin_pw2_0_), .B(
        SBOX_FF4_out[30]), .Z(SBOX_Inst_f5_ph[2]) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_NxGAMMA_U3 ( .A(SBOX_Inst_f5_phwillwin_pw2_5_), .B(SBOX_FF4_out[29]), .Z(SBOX_Inst_f5_phwillwin_pw2_4_) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_NxGAMMA_U2 ( .A(SBOX_Inst_f5_phwillwin_pw2_3_), .B(SBOX_FF4_out[27]), .Z(SBOX_Inst_f5_phwillwin_pw2_2_) );
  XOR2_X1 SBOX_Inst_f5_phwillwin_NxGAMMA_U1 ( .A(SBOX_Inst_f5_phwillwin_pw2_1_), .B(SBOX_FF4_out[25]), .Z(SBOX_Inst_f5_phwillwin_pw2_0_) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U12 ( .A(SBOX_Inst_f5_plwillwin_pw2_4_), .B(
        SBOX_FF4_out[16]), .Z(SBOX_Inst_f5_pl[10]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U11 ( .A(SBOX_Inst_f5_plwillwin_pw2_2_), .B(
        SBOX_FF4_out[14]), .Z(SBOX_Inst_f5_pl[6]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U10 ( .A(SBOX_Inst_f5_plwillwin_pw2_0_), .B(
        SBOX_FF4_out[12]), .Z(SBOX_Inst_f5_pl[2]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U9 ( .A(SBOX_Inst_f5_plwillwin_pw2_2_), .B(
        SBOX_FF4_out[2]), .Z(SBOX_Inst_f5_pl[4]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U8 ( .A(SBOX_Inst_f5_plwillwin_pw2_4_), .B(
        SBOX_FF4_out[4]), .Z(SBOX_Inst_f5_pl[8]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U7 ( .A(SBOX_Inst_f5_plwillwin_pw2_0_), .B(
        SBOX_FF4_out[0]), .Z(SBOX_Inst_f5_pl[0]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U6 ( .A(SBOX_Inst_f5_plwillwin_pw2_5_), .B(
        SBOX_FF4_out[5]), .Z(SBOX_Inst_f5_pl[9]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U5 ( .A(SBOX_Inst_f5_plwillwin_pw2_3_), .B(
        SBOX_FF4_out[3]), .Z(SBOX_Inst_f5_pl[5]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U4 ( .A(SBOX_Inst_f5_plwillwin_pw2_1_), .B(
        SBOX_FF4_out[1]), .Z(SBOX_Inst_f5_pl[1]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U3 ( .A(SBOX_Inst_f5_plwillwin_pw2_5_), .B(
        SBOX_FF4_out[17]), .Z(SBOX_Inst_f5_pl[11]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U2 ( .A(SBOX_Inst_f5_plwillwin_pw2_3_), .B(
        SBOX_FF4_out[15]), .Z(SBOX_Inst_f5_pl[7]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_U1 ( .A(SBOX_Inst_f5_plwillwin_pw2_1_), .B(
        SBOX_FF4_out[13]), .Z(SBOX_Inst_f5_pl[3]) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_NxGAMMA_U3 ( .A(SBOX_Inst_f5_plwillwin_pw2_5_), .B(SBOX_FF4_out[11]), .Z(SBOX_Inst_f5_plwillwin_pw2_4_) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_NxGAMMA_U2 ( .A(SBOX_Inst_f5_plwillwin_pw2_3_), .B(SBOX_FF4_out[9]), .Z(SBOX_Inst_f5_plwillwin_pw2_2_) );
  XOR2_X1 SBOX_Inst_f5_plwillwin_NxGAMMA_U1 ( .A(SBOX_Inst_f5_plwillwin_pw2_1_), .B(SBOX_FF4_out[7]), .Z(SBOX_Inst_f5_plwillwin_pw2_0_) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U33 ( .A(SBOX_Inst_f5_ph[8]), .B(
        SBOX_Inst_f5_invlinearMapping_n6), .ZN(SBOX_Qoutput[17]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U32 ( .A(SBOX_Inst_f5_pl[9]), .B(
        SBOX_Inst_f5_ph[9]), .Z(SBOX_Inst_f5_invlinearMapping_n6) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U31 ( .A(SBOX_Inst_f5_ph[4]), .B(
        SBOX_Inst_f5_invlinearMapping_n5), .ZN(SBOX_Qoutput[9]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U30 ( .A(SBOX_Inst_f5_pl[5]), .B(
        SBOX_Inst_f5_ph[5]), .Z(SBOX_Inst_f5_invlinearMapping_n5) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U29 ( .A(SBOX_Inst_f5_ph[0]), .B(
        SBOX_Inst_f5_invlinearMapping_n4), .ZN(SBOX_Qoutput[1]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U28 ( .A(SBOX_Inst_f5_pl[1]), .B(
        SBOX_Inst_f5_ph[1]), .Z(SBOX_Inst_f5_invlinearMapping_n4) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U27 ( .A(SBOX_Inst_f5_pl[9]), .B(
        SBOX_Inst_f5_invlinearMapping_n7), .Z(SBOX_Qoutput[16]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U26 ( .A(SBOX_Inst_f5_pl[5]), .B(
        SBOX_Inst_f5_invlinearMapping_n9), .Z(SBOX_Qoutput[8]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U25 ( .A(SBOX_Inst_f5_pl[1]), .B(
        SBOX_Inst_f5_invlinearMapping_n8), .Z(SBOX_Qoutput[0]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U24 ( .A(SBOX_Qoutput[20]), .B(
        SBOX_Inst_f5_invlinearMapping_n7), .ZN(SBOX_Qoutput[19]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U23 ( .A(SBOX_Qoutput[12]), .B(
        SBOX_Inst_f5_invlinearMapping_n9), .ZN(SBOX_Qoutput[11]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U22 ( .A(SBOX_Qoutput[4]), .B(
        SBOX_Inst_f5_invlinearMapping_n8), .ZN(SBOX_Qoutput[3]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U21 ( .A(SBOX_Inst_f5_pl[10]), .B(
        SBOX_Inst_f5_invlinearMapping_n3), .ZN(SBOX_Qoutput[18]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U20 ( .A(SBOX_Qoutput[21]), .B(
        SBOX_Qoutput[23]), .Z(SBOX_Inst_f5_invlinearMapping_n3) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U19 ( .A(SBOX_Inst_f5_pl[6]), .B(
        SBOX_Inst_f5_invlinearMapping_n2), .ZN(SBOX_Qoutput[10]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U18 ( .A(SBOX_Qoutput[13]), .B(
        SBOX_Qoutput[15]), .Z(SBOX_Inst_f5_invlinearMapping_n2) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U17 ( .A(SBOX_Inst_f5_pl[2]), .B(
        SBOX_Inst_f5_invlinearMapping_n1), .ZN(SBOX_Qoutput[2]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U16 ( .A(SBOX_Qoutput[5]), .B(
        SBOX_Qoutput[7]), .Z(SBOX_Inst_f5_invlinearMapping_n1) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U15 ( .A(SBOX_Inst_f5_pl[11]), .B(
        SBOX_Inst_f5_ph[11]), .ZN(SBOX_Qoutput[22]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U14 ( .A(SBOX_Inst_f5_ph[6]), .B(
        SBOX_Inst_f5_pl[4]), .ZN(SBOX_Qoutput[13]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U13 ( .A(SBOX_Inst_f5_pl[3]), .B(
        SBOX_Inst_f5_ph[3]), .ZN(SBOX_Qoutput[6]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U12 ( .A(SBOX_Inst_f5_ph[10]), .B(
        SBOX_Inst_f5_pl[8]), .ZN(SBOX_Qoutput[21]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U11 ( .A(SBOX_Inst_f5_pl[7]), .B(
        SBOX_Inst_f5_ph[7]), .ZN(SBOX_Qoutput[14]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U10 ( .A(SBOX_Inst_f5_ph[2]), .B(
        SBOX_Inst_f5_pl[0]), .ZN(SBOX_Qoutput[5]) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U9 ( .A(SBOX_Inst_f5_ph[9]), .B(
        SBOX_Inst_f5_pl[11]), .Z(SBOX_Qoutput[23]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U8 ( .A(SBOX_Inst_f5_ph[9]), .B(
        SBOX_Qoutput[22]), .ZN(SBOX_Qoutput[20]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U7 ( .A(SBOX_Inst_f5_ph[10]), .B(
        SBOX_Inst_f5_ph[8]), .ZN(SBOX_Inst_f5_invlinearMapping_n7) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U6 ( .A(SBOX_Inst_f5_ph[5]), .B(
        SBOX_Inst_f5_pl[7]), .Z(SBOX_Qoutput[15]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U5 ( .A(SBOX_Inst_f5_ph[5]), .B(
        SBOX_Qoutput[14]), .ZN(SBOX_Qoutput[12]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U4 ( .A(SBOX_Inst_f5_ph[6]), .B(
        SBOX_Inst_f5_ph[4]), .ZN(SBOX_Inst_f5_invlinearMapping_n9) );
  XOR2_X1 SBOX_Inst_f5_invlinearMapping_U3 ( .A(SBOX_Inst_f5_ph[1]), .B(
        SBOX_Inst_f5_pl[3]), .Z(SBOX_Qoutput[7]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U2 ( .A(SBOX_Inst_f5_ph[1]), .B(
        SBOX_Qoutput[6]), .ZN(SBOX_Qoutput[4]) );
  XNOR2_X1 SBOX_Inst_f5_invlinearMapping_U1 ( .A(SBOX_Inst_f5_ph[2]), .B(
        SBOX_Inst_f5_ph[0]), .ZN(SBOX_Inst_f5_invlinearMapping_n8) );
  OAI21_X1 SBOX_PL_5_U49 ( .B1(1'b1), .B2(SBOX_PL_5_n97), .A(SBOX_PL_5_n168), 
        .ZN(SBOX_PL_5_n73) );
  NAND2_X1 SBOX_PL_5_U48 ( .A1(1'b1), .A2(SBOX_Qoutput[23]), .ZN(
        SBOX_PL_5_n168) );
  OAI21_X1 SBOX_PL_5_U47 ( .B1(1'b1), .B2(SBOX_PL_5_n99), .A(SBOX_PL_5_n167), 
        .ZN(SBOX_PL_5_n75) );
  NAND2_X1 SBOX_PL_5_U46 ( .A1(1'b1), .A2(SBOX_Qoutput[21]), .ZN(
        SBOX_PL_5_n167) );
  OAI21_X1 SBOX_PL_5_U45 ( .B1(1'b1), .B2(SBOX_PL_5_n105), .A(SBOX_PL_5_n166), 
        .ZN(SBOX_PL_5_n81) );
  NAND2_X1 SBOX_PL_5_U44 ( .A1(1'b1), .A2(SBOX_Qoutput[15]), .ZN(
        SBOX_PL_5_n166) );
  OAI21_X1 SBOX_PL_5_U43 ( .B1(1'b1), .B2(SBOX_PL_5_n107), .A(SBOX_PL_5_n165), 
        .ZN(SBOX_PL_5_n83) );
  NAND2_X1 SBOX_PL_5_U42 ( .A1(1'b1), .A2(SBOX_Qoutput[13]), .ZN(
        SBOX_PL_5_n165) );
  OAI21_X1 SBOX_PL_5_U41 ( .B1(1'b1), .B2(SBOX_PL_5_n113), .A(SBOX_PL_5_n164), 
        .ZN(SBOX_PL_5_n89) );
  NAND2_X1 SBOX_PL_5_U40 ( .A1(1'b1), .A2(SBOX_Qoutput[7]), .ZN(SBOX_PL_5_n164) );
  OAI21_X1 SBOX_PL_5_U39 ( .B1(1'b1), .B2(SBOX_PL_5_n115), .A(SBOX_PL_5_n163), 
        .ZN(SBOX_PL_5_n91) );
  NAND2_X1 SBOX_PL_5_U38 ( .A1(1'b1), .A2(SBOX_Qoutput[5]), .ZN(SBOX_PL_5_n163) );
  OAI21_X1 SBOX_PL_5_U37 ( .B1(1'b1), .B2(SBOX_PL_5_n98), .A(SBOX_PL_5_n162), 
        .ZN(SBOX_PL_5_n74) );
  NAND2_X1 SBOX_PL_5_U36 ( .A1(1'b1), .A2(SBOX_Qoutput[22]), .ZN(
        SBOX_PL_5_n162) );
  OAI21_X1 SBOX_PL_5_U35 ( .B1(1'b1), .B2(SBOX_PL_5_n103), .A(SBOX_PL_5_n161), 
        .ZN(SBOX_PL_5_n79) );
  NAND2_X1 SBOX_PL_5_U34 ( .A1(1'b1), .A2(SBOX_Qoutput[17]), .ZN(
        SBOX_PL_5_n161) );
  OAI21_X1 SBOX_PL_5_U33 ( .B1(1'b1), .B2(SBOX_PL_5_n106), .A(SBOX_PL_5_n160), 
        .ZN(SBOX_PL_5_n82) );
  NAND2_X1 SBOX_PL_5_U32 ( .A1(1'b1), .A2(SBOX_Qoutput[14]), .ZN(
        SBOX_PL_5_n160) );
  OAI21_X1 SBOX_PL_5_U31 ( .B1(1'b1), .B2(SBOX_PL_5_n111), .A(SBOX_PL_5_n159), 
        .ZN(SBOX_PL_5_n87) );
  NAND2_X1 SBOX_PL_5_U30 ( .A1(1'b1), .A2(SBOX_Qoutput[9]), .ZN(SBOX_PL_5_n159) );
  OAI21_X1 SBOX_PL_5_U29 ( .B1(1'b1), .B2(SBOX_PL_5_n114), .A(SBOX_PL_5_n158), 
        .ZN(SBOX_PL_5_n90) );
  NAND2_X1 SBOX_PL_5_U28 ( .A1(1'b1), .A2(SBOX_Qoutput[6]), .ZN(SBOX_PL_5_n158) );
  OAI21_X1 SBOX_PL_5_U27 ( .B1(1'b1), .B2(SBOX_PL_5_n119), .A(SBOX_PL_5_n157), 
        .ZN(SBOX_PL_5_n95) );
  NAND2_X1 SBOX_PL_5_U26 ( .A1(1'b1), .A2(SBOX_Qoutput[1]), .ZN(SBOX_PL_5_n157) );
  OAI21_X1 SBOX_PL_5_U25 ( .B1(1'b1), .B2(SBOX_PL_5_n100), .A(SBOX_PL_5_n156), 
        .ZN(SBOX_PL_5_n76) );
  NAND2_X1 SBOX_PL_5_U24 ( .A1(1'b1), .A2(SBOX_Qoutput[20]), .ZN(
        SBOX_PL_5_n156) );
  OAI21_X1 SBOX_PL_5_U23 ( .B1(1'b1), .B2(SBOX_PL_5_n104), .A(SBOX_PL_5_n155), 
        .ZN(SBOX_PL_5_n80) );
  NAND2_X1 SBOX_PL_5_U22 ( .A1(1'b1), .A2(SBOX_Qoutput[16]), .ZN(
        SBOX_PL_5_n155) );
  OAI21_X1 SBOX_PL_5_U21 ( .B1(1'b1), .B2(SBOX_PL_5_n108), .A(SBOX_PL_5_n154), 
        .ZN(SBOX_PL_5_n84) );
  NAND2_X1 SBOX_PL_5_U20 ( .A1(1'b1), .A2(SBOX_Qoutput[12]), .ZN(
        SBOX_PL_5_n154) );
  OAI21_X1 SBOX_PL_5_U19 ( .B1(1'b1), .B2(SBOX_PL_5_n112), .A(SBOX_PL_5_n153), 
        .ZN(SBOX_PL_5_n88) );
  NAND2_X1 SBOX_PL_5_U18 ( .A1(1'b1), .A2(SBOX_Qoutput[8]), .ZN(SBOX_PL_5_n153) );
  OAI21_X1 SBOX_PL_5_U17 ( .B1(1'b1), .B2(SBOX_PL_5_n116), .A(SBOX_PL_5_n152), 
        .ZN(SBOX_PL_5_n92) );
  NAND2_X1 SBOX_PL_5_U16 ( .A1(1'b1), .A2(SBOX_Qoutput[4]), .ZN(SBOX_PL_5_n152) );
  OAI21_X1 SBOX_PL_5_U15 ( .B1(1'b1), .B2(SBOX_PL_5_n120), .A(SBOX_PL_5_n151), 
        .ZN(SBOX_PL_5_n96) );
  NAND2_X1 SBOX_PL_5_U14 ( .A1(1'b1), .A2(SBOX_Qoutput[0]), .ZN(SBOX_PL_5_n151) );
  OAI21_X1 SBOX_PL_5_U13 ( .B1(1'b1), .B2(SBOX_PL_5_n101), .A(SBOX_PL_5_n150), 
        .ZN(SBOX_PL_5_n77) );
  NAND2_X1 SBOX_PL_5_U12 ( .A1(1'b1), .A2(SBOX_Qoutput[19]), .ZN(
        SBOX_PL_5_n150) );
  OAI21_X1 SBOX_PL_5_U11 ( .B1(1'b1), .B2(SBOX_PL_5_n109), .A(SBOX_PL_5_n149), 
        .ZN(SBOX_PL_5_n85) );
  NAND2_X1 SBOX_PL_5_U10 ( .A1(1'b1), .A2(SBOX_Qoutput[11]), .ZN(
        SBOX_PL_5_n149) );
  OAI21_X1 SBOX_PL_5_U9 ( .B1(1'b1), .B2(SBOX_PL_5_n117), .A(SBOX_PL_5_n148), 
        .ZN(SBOX_PL_5_n93) );
  NAND2_X1 SBOX_PL_5_U8 ( .A1(1'b1), .A2(SBOX_Qoutput[3]), .ZN(SBOX_PL_5_n148)
         );
  OAI21_X1 SBOX_PL_5_U7 ( .B1(1'b1), .B2(SBOX_PL_5_n102), .A(SBOX_PL_5_n147), 
        .ZN(SBOX_PL_5_n78) );
  NAND2_X1 SBOX_PL_5_U6 ( .A1(1'b1), .A2(SBOX_Qoutput[18]), .ZN(SBOX_PL_5_n147) );
  OAI21_X1 SBOX_PL_5_U5 ( .B1(1'b1), .B2(SBOX_PL_5_n110), .A(SBOX_PL_5_n146), 
        .ZN(SBOX_PL_5_n86) );
  NAND2_X1 SBOX_PL_5_U4 ( .A1(1'b1), .A2(SBOX_Qoutput[10]), .ZN(SBOX_PL_5_n146) );
  OAI21_X1 SBOX_PL_5_U3 ( .B1(1'b1), .B2(SBOX_PL_5_n118), .A(SBOX_PL_5_n145), 
        .ZN(SBOX_PL_5_n94) );
  NAND2_X1 SBOX_PL_5_U2 ( .A1(1'b1), .A2(SBOX_Qoutput[2]), .ZN(SBOX_PL_5_n145)
         );
  DFF_X1 SBOX_PL_5_s_current_state_reg_0_ ( .D(SBOX_PL_5_n96), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[0]), .QN(SBOX_PL_5_n120) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_1_ ( .D(SBOX_PL_5_n95), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[1]), .QN(SBOX_PL_5_n119) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_2_ ( .D(SBOX_PL_5_n94), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[2]), .QN(SBOX_PL_5_n118) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_3_ ( .D(SBOX_PL_5_n93), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[3]), .QN(SBOX_PL_5_n117) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_4_ ( .D(SBOX_PL_5_n92), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[4]), .QN(SBOX_PL_5_n116) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_5_ ( .D(SBOX_PL_5_n91), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[5]), .QN(SBOX_PL_5_n115) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_6_ ( .D(SBOX_PL_5_n90), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[6]), .QN(SBOX_PL_5_n114) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_7_ ( .D(SBOX_PL_5_n89), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[7]), .QN(SBOX_PL_5_n113) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_8_ ( .D(SBOX_PL_5_n88), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[8]), .QN(SBOX_PL_5_n112) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_9_ ( .D(SBOX_PL_5_n87), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[9]), .QN(SBOX_PL_5_n111) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_10_ ( .D(SBOX_PL_5_n86), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[10]), .QN(SBOX_PL_5_n110) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_11_ ( .D(SBOX_PL_5_n85), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[11]), .QN(SBOX_PL_5_n109) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_12_ ( .D(SBOX_PL_5_n84), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[12]), .QN(SBOX_PL_5_n108) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_13_ ( .D(SBOX_PL_5_n83), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[13]), .QN(SBOX_PL_5_n107) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_14_ ( .D(SBOX_PL_5_n82), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[14]), .QN(SBOX_PL_5_n106) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_15_ ( .D(SBOX_PL_5_n81), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[15]), .QN(SBOX_PL_5_n105) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_16_ ( .D(SBOX_PL_5_n80), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[16]), .QN(SBOX_PL_5_n104) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_17_ ( .D(SBOX_PL_5_n79), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[17]), .QN(SBOX_PL_5_n103) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_18_ ( .D(SBOX_PL_5_n78), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[18]), .QN(SBOX_PL_5_n102) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_19_ ( .D(SBOX_PL_5_n77), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[19]), .QN(SBOX_PL_5_n101) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_20_ ( .D(SBOX_PL_5_n76), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[20]), .QN(SBOX_PL_5_n100) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_21_ ( .D(SBOX_PL_5_n75), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[21]), .QN(SBOX_PL_5_n99) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_22_ ( .D(SBOX_PL_5_n74), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[22]), .QN(SBOX_PL_5_n98) );
  DFF_X1 SBOX_PL_5_s_current_state_reg_23_ ( .D(SBOX_PL_5_n73), .CK(ClkxCI), 
        .Q(SBOX_Qreg5[23]), .QN(SBOX_PL_5_n97) );
  OAI21_X1 SBOX_PL_6_U49 ( .B1(1'b1), .B2(SBOX_PL_6_n120), .A(SBOX_PL_6_n168), 
        .ZN(SBOX_PL_6_n96) );
  NAND2_X1 SBOX_PL_6_U48 ( .A1(1'b1), .A2(SBOX_Qreg5[0]), .ZN(SBOX_PL_6_n168)
         );
  OAI21_X1 SBOX_PL_6_U47 ( .B1(1'b1), .B2(SBOX_PL_6_n119), .A(SBOX_PL_6_n167), 
        .ZN(SBOX_PL_6_n95) );
  NAND2_X1 SBOX_PL_6_U46 ( .A1(1'b1), .A2(SBOX_Qreg5[1]), .ZN(SBOX_PL_6_n167)
         );
  OAI21_X1 SBOX_PL_6_U45 ( .B1(1'b1), .B2(SBOX_PL_6_n118), .A(SBOX_PL_6_n166), 
        .ZN(SBOX_PL_6_n94) );
  NAND2_X1 SBOX_PL_6_U44 ( .A1(1'b1), .A2(SBOX_Qreg5[2]), .ZN(SBOX_PL_6_n166)
         );
  OAI21_X1 SBOX_PL_6_U43 ( .B1(1'b1), .B2(SBOX_PL_6_n117), .A(SBOX_PL_6_n165), 
        .ZN(SBOX_PL_6_n93) );
  NAND2_X1 SBOX_PL_6_U42 ( .A1(1'b1), .A2(SBOX_Qreg5[3]), .ZN(SBOX_PL_6_n165)
         );
  OAI21_X1 SBOX_PL_6_U41 ( .B1(1'b1), .B2(SBOX_PL_6_n116), .A(SBOX_PL_6_n164), 
        .ZN(SBOX_PL_6_n92) );
  NAND2_X1 SBOX_PL_6_U40 ( .A1(1'b1), .A2(SBOX_Qreg5[4]), .ZN(SBOX_PL_6_n164)
         );
  OAI21_X1 SBOX_PL_6_U39 ( .B1(1'b1), .B2(SBOX_PL_6_n115), .A(SBOX_PL_6_n163), 
        .ZN(SBOX_PL_6_n91) );
  NAND2_X1 SBOX_PL_6_U38 ( .A1(1'b1), .A2(SBOX_Qreg5[5]), .ZN(SBOX_PL_6_n163)
         );
  OAI21_X1 SBOX_PL_6_U37 ( .B1(1'b1), .B2(SBOX_PL_6_n114), .A(SBOX_PL_6_n162), 
        .ZN(SBOX_PL_6_n90) );
  NAND2_X1 SBOX_PL_6_U36 ( .A1(1'b1), .A2(SBOX_Qreg5[6]), .ZN(SBOX_PL_6_n162)
         );
  OAI21_X1 SBOX_PL_6_U35 ( .B1(1'b1), .B2(SBOX_PL_6_n113), .A(SBOX_PL_6_n161), 
        .ZN(SBOX_PL_6_n89) );
  NAND2_X1 SBOX_PL_6_U34 ( .A1(1'b1), .A2(SBOX_Qreg5[7]), .ZN(SBOX_PL_6_n161)
         );
  OAI21_X1 SBOX_PL_6_U33 ( .B1(1'b1), .B2(SBOX_PL_6_n112), .A(SBOX_PL_6_n160), 
        .ZN(SBOX_PL_6_n88) );
  NAND2_X1 SBOX_PL_6_U32 ( .A1(1'b1), .A2(SBOX_Qreg5[8]), .ZN(SBOX_PL_6_n160)
         );
  OAI21_X1 SBOX_PL_6_U31 ( .B1(1'b1), .B2(SBOX_PL_6_n111), .A(SBOX_PL_6_n159), 
        .ZN(SBOX_PL_6_n87) );
  NAND2_X1 SBOX_PL_6_U30 ( .A1(1'b1), .A2(SBOX_Qreg5[9]), .ZN(SBOX_PL_6_n159)
         );
  OAI21_X1 SBOX_PL_6_U29 ( .B1(1'b1), .B2(SBOX_PL_6_n110), .A(SBOX_PL_6_n158), 
        .ZN(SBOX_PL_6_n86) );
  NAND2_X1 SBOX_PL_6_U28 ( .A1(1'b1), .A2(SBOX_Qreg5[10]), .ZN(SBOX_PL_6_n158)
         );
  OAI21_X1 SBOX_PL_6_U27 ( .B1(1'b1), .B2(SBOX_PL_6_n109), .A(SBOX_PL_6_n157), 
        .ZN(SBOX_PL_6_n85) );
  NAND2_X1 SBOX_PL_6_U26 ( .A1(1'b1), .A2(SBOX_Qreg5[11]), .ZN(SBOX_PL_6_n157)
         );
  OAI21_X1 SBOX_PL_6_U25 ( .B1(1'b1), .B2(SBOX_PL_6_n108), .A(SBOX_PL_6_n156), 
        .ZN(SBOX_PL_6_n84) );
  NAND2_X1 SBOX_PL_6_U24 ( .A1(1'b1), .A2(SBOX_Qreg5[12]), .ZN(SBOX_PL_6_n156)
         );
  OAI21_X1 SBOX_PL_6_U23 ( .B1(1'b1), .B2(SBOX_PL_6_n107), .A(SBOX_PL_6_n155), 
        .ZN(SBOX_PL_6_n83) );
  NAND2_X1 SBOX_PL_6_U22 ( .A1(1'b1), .A2(SBOX_Qreg5[13]), .ZN(SBOX_PL_6_n155)
         );
  OAI21_X1 SBOX_PL_6_U21 ( .B1(1'b1), .B2(SBOX_PL_6_n106), .A(SBOX_PL_6_n154), 
        .ZN(SBOX_PL_6_n82) );
  NAND2_X1 SBOX_PL_6_U20 ( .A1(1'b1), .A2(SBOX_Qreg5[14]), .ZN(SBOX_PL_6_n154)
         );
  OAI21_X1 SBOX_PL_6_U19 ( .B1(1'b1), .B2(SBOX_PL_6_n105), .A(SBOX_PL_6_n153), 
        .ZN(SBOX_PL_6_n81) );
  NAND2_X1 SBOX_PL_6_U18 ( .A1(1'b1), .A2(SBOX_Qreg5[15]), .ZN(SBOX_PL_6_n153)
         );
  OAI21_X1 SBOX_PL_6_U17 ( .B1(1'b1), .B2(SBOX_PL_6_n104), .A(SBOX_PL_6_n152), 
        .ZN(SBOX_PL_6_n80) );
  NAND2_X1 SBOX_PL_6_U16 ( .A1(1'b1), .A2(SBOX_Qreg5[16]), .ZN(SBOX_PL_6_n152)
         );
  OAI21_X1 SBOX_PL_6_U15 ( .B1(1'b1), .B2(SBOX_PL_6_n103), .A(SBOX_PL_6_n151), 
        .ZN(SBOX_PL_6_n79) );
  NAND2_X1 SBOX_PL_6_U14 ( .A1(1'b1), .A2(SBOX_Qreg5[17]), .ZN(SBOX_PL_6_n151)
         );
  OAI21_X1 SBOX_PL_6_U13 ( .B1(1'b1), .B2(SBOX_PL_6_n102), .A(SBOX_PL_6_n150), 
        .ZN(SBOX_PL_6_n78) );
  NAND2_X1 SBOX_PL_6_U12 ( .A1(1'b1), .A2(SBOX_Qreg5[18]), .ZN(SBOX_PL_6_n150)
         );
  OAI21_X1 SBOX_PL_6_U11 ( .B1(1'b1), .B2(SBOX_PL_6_n101), .A(SBOX_PL_6_n149), 
        .ZN(SBOX_PL_6_n77) );
  NAND2_X1 SBOX_PL_6_U10 ( .A1(1'b1), .A2(SBOX_Qreg5[19]), .ZN(SBOX_PL_6_n149)
         );
  OAI21_X1 SBOX_PL_6_U9 ( .B1(1'b1), .B2(SBOX_PL_6_n100), .A(SBOX_PL_6_n148), 
        .ZN(SBOX_PL_6_n76) );
  NAND2_X1 SBOX_PL_6_U8 ( .A1(1'b1), .A2(SBOX_Qreg5[20]), .ZN(SBOX_PL_6_n148)
         );
  OAI21_X1 SBOX_PL_6_U7 ( .B1(1'b1), .B2(SBOX_PL_6_n99), .A(SBOX_PL_6_n147), 
        .ZN(SBOX_PL_6_n75) );
  NAND2_X1 SBOX_PL_6_U6 ( .A1(1'b1), .A2(SBOX_Qreg5[21]), .ZN(SBOX_PL_6_n147)
         );
  OAI21_X1 SBOX_PL_6_U5 ( .B1(1'b1), .B2(SBOX_PL_6_n98), .A(SBOX_PL_6_n146), 
        .ZN(SBOX_PL_6_n74) );
  NAND2_X1 SBOX_PL_6_U4 ( .A1(1'b1), .A2(SBOX_Qreg5[22]), .ZN(SBOX_PL_6_n146)
         );
  OAI21_X1 SBOX_PL_6_U3 ( .B1(1'b1), .B2(SBOX_PL_6_n97), .A(SBOX_PL_6_n145), 
        .ZN(SBOX_PL_6_n73) );
  NAND2_X1 SBOX_PL_6_U2 ( .A1(1'b1), .A2(SBOX_Qreg5[23]), .ZN(SBOX_PL_6_n145)
         );
  DFF_X1 SBOX_PL_6_s_current_state_reg_0_ ( .D(SBOX_PL_6_n96), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[0]), .QN(SBOX_PL_6_n120) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_1_ ( .D(SBOX_PL_6_n95), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[1]), .QN(SBOX_PL_6_n119) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_2_ ( .D(SBOX_PL_6_n94), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[2]), .QN(SBOX_PL_6_n118) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_3_ ( .D(SBOX_PL_6_n93), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[3]), .QN(SBOX_PL_6_n117) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_4_ ( .D(SBOX_PL_6_n92), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[4]), .QN(SBOX_PL_6_n116) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_5_ ( .D(SBOX_PL_6_n91), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[5]), .QN(SBOX_PL_6_n115) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_6_ ( .D(SBOX_PL_6_n90), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[6]), .QN(SBOX_PL_6_n114) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_7_ ( .D(SBOX_PL_6_n89), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[7]), .QN(SBOX_PL_6_n113) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_8_ ( .D(SBOX_PL_6_n88), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[8]), .QN(SBOX_PL_6_n112) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_9_ ( .D(SBOX_PL_6_n87), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[9]), .QN(SBOX_PL_6_n111) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_10_ ( .D(SBOX_PL_6_n86), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[10]), .QN(SBOX_PL_6_n110) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_11_ ( .D(SBOX_PL_6_n85), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[11]), .QN(SBOX_PL_6_n109) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_12_ ( .D(SBOX_PL_6_n84), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[12]), .QN(SBOX_PL_6_n108) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_13_ ( .D(SBOX_PL_6_n83), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[13]), .QN(SBOX_PL_6_n107) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_14_ ( .D(SBOX_PL_6_n82), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[14]), .QN(SBOX_PL_6_n106) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_15_ ( .D(SBOX_PL_6_n81), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[15]), .QN(SBOX_PL_6_n105) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_16_ ( .D(SBOX_PL_6_n80), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[16]), .QN(SBOX_PL_6_n104) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_17_ ( .D(SBOX_PL_6_n79), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[17]), .QN(SBOX_PL_6_n103) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_18_ ( .D(SBOX_PL_6_n78), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[18]), .QN(SBOX_PL_6_n102) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_19_ ( .D(SBOX_PL_6_n77), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[19]), .QN(SBOX_PL_6_n101) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_20_ ( .D(SBOX_PL_6_n76), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[20]), .QN(SBOX_PL_6_n100) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_21_ ( .D(SBOX_PL_6_n75), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[21]), .QN(SBOX_PL_6_n99) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_22_ ( .D(SBOX_PL_6_n74), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[22]), .QN(SBOX_PL_6_n98) );
  DFF_X1 SBOX_PL_6_s_current_state_reg_23_ ( .D(SBOX_PL_6_n73), .CK(ClkxCI), 
        .Q(SBOX_Qreg6[23]), .QN(SBOX_PL_6_n97) );
  OAI21_X1 SBOX_PL_7_U49 ( .B1(1'b1), .B2(SBOX_PL_7_n120), .A(SBOX_PL_7_n168), 
        .ZN(SBOX_PL_7_n96) );
  NAND2_X1 SBOX_PL_7_U48 ( .A1(1'b1), .A2(SBOX_Qreg6[0]), .ZN(SBOX_PL_7_n168)
         );
  OAI21_X1 SBOX_PL_7_U47 ( .B1(1'b1), .B2(SBOX_PL_7_n119), .A(SBOX_PL_7_n167), 
        .ZN(SBOX_PL_7_n95) );
  NAND2_X1 SBOX_PL_7_U46 ( .A1(1'b1), .A2(SBOX_Qreg6[1]), .ZN(SBOX_PL_7_n167)
         );
  OAI21_X1 SBOX_PL_7_U45 ( .B1(1'b1), .B2(SBOX_PL_7_n118), .A(SBOX_PL_7_n166), 
        .ZN(SBOX_PL_7_n94) );
  NAND2_X1 SBOX_PL_7_U44 ( .A1(1'b1), .A2(SBOX_Qreg6[2]), .ZN(SBOX_PL_7_n166)
         );
  OAI21_X1 SBOX_PL_7_U43 ( .B1(1'b1), .B2(SBOX_PL_7_n117), .A(SBOX_PL_7_n165), 
        .ZN(SBOX_PL_7_n93) );
  NAND2_X1 SBOX_PL_7_U42 ( .A1(1'b1), .A2(SBOX_Qreg6[3]), .ZN(SBOX_PL_7_n165)
         );
  OAI21_X1 SBOX_PL_7_U41 ( .B1(1'b1), .B2(SBOX_PL_7_n116), .A(SBOX_PL_7_n164), 
        .ZN(SBOX_PL_7_n92) );
  NAND2_X1 SBOX_PL_7_U40 ( .A1(1'b1), .A2(SBOX_Qreg6[4]), .ZN(SBOX_PL_7_n164)
         );
  OAI21_X1 SBOX_PL_7_U39 ( .B1(1'b1), .B2(SBOX_PL_7_n115), .A(SBOX_PL_7_n163), 
        .ZN(SBOX_PL_7_n91) );
  NAND2_X1 SBOX_PL_7_U38 ( .A1(1'b1), .A2(SBOX_Qreg6[5]), .ZN(SBOX_PL_7_n163)
         );
  OAI21_X1 SBOX_PL_7_U37 ( .B1(1'b1), .B2(SBOX_PL_7_n114), .A(SBOX_PL_7_n162), 
        .ZN(SBOX_PL_7_n90) );
  NAND2_X1 SBOX_PL_7_U36 ( .A1(1'b1), .A2(SBOX_Qreg6[6]), .ZN(SBOX_PL_7_n162)
         );
  OAI21_X1 SBOX_PL_7_U35 ( .B1(1'b1), .B2(SBOX_PL_7_n113), .A(SBOX_PL_7_n161), 
        .ZN(SBOX_PL_7_n89) );
  NAND2_X1 SBOX_PL_7_U34 ( .A1(1'b1), .A2(SBOX_Qreg6[7]), .ZN(SBOX_PL_7_n161)
         );
  OAI21_X1 SBOX_PL_7_U33 ( .B1(1'b1), .B2(SBOX_PL_7_n112), .A(SBOX_PL_7_n160), 
        .ZN(SBOX_PL_7_n88) );
  NAND2_X1 SBOX_PL_7_U32 ( .A1(1'b1), .A2(SBOX_Qreg6[8]), .ZN(SBOX_PL_7_n160)
         );
  OAI21_X1 SBOX_PL_7_U31 ( .B1(1'b1), .B2(SBOX_PL_7_n111), .A(SBOX_PL_7_n159), 
        .ZN(SBOX_PL_7_n87) );
  NAND2_X1 SBOX_PL_7_U30 ( .A1(1'b1), .A2(SBOX_Qreg6[9]), .ZN(SBOX_PL_7_n159)
         );
  OAI21_X1 SBOX_PL_7_U29 ( .B1(1'b1), .B2(SBOX_PL_7_n110), .A(SBOX_PL_7_n158), 
        .ZN(SBOX_PL_7_n86) );
  NAND2_X1 SBOX_PL_7_U28 ( .A1(1'b1), .A2(SBOX_Qreg6[10]), .ZN(SBOX_PL_7_n158)
         );
  OAI21_X1 SBOX_PL_7_U27 ( .B1(1'b1), .B2(SBOX_PL_7_n109), .A(SBOX_PL_7_n157), 
        .ZN(SBOX_PL_7_n85) );
  NAND2_X1 SBOX_PL_7_U26 ( .A1(1'b1), .A2(SBOX_Qreg6[11]), .ZN(SBOX_PL_7_n157)
         );
  OAI21_X1 SBOX_PL_7_U25 ( .B1(1'b1), .B2(SBOX_PL_7_n108), .A(SBOX_PL_7_n156), 
        .ZN(SBOX_PL_7_n84) );
  NAND2_X1 SBOX_PL_7_U24 ( .A1(1'b1), .A2(SBOX_Qreg6[12]), .ZN(SBOX_PL_7_n156)
         );
  OAI21_X1 SBOX_PL_7_U23 ( .B1(1'b1), .B2(SBOX_PL_7_n107), .A(SBOX_PL_7_n155), 
        .ZN(SBOX_PL_7_n83) );
  NAND2_X1 SBOX_PL_7_U22 ( .A1(1'b1), .A2(SBOX_Qreg6[13]), .ZN(SBOX_PL_7_n155)
         );
  OAI21_X1 SBOX_PL_7_U21 ( .B1(1'b1), .B2(SBOX_PL_7_n106), .A(SBOX_PL_7_n154), 
        .ZN(SBOX_PL_7_n82) );
  NAND2_X1 SBOX_PL_7_U20 ( .A1(1'b1), .A2(SBOX_Qreg6[14]), .ZN(SBOX_PL_7_n154)
         );
  OAI21_X1 SBOX_PL_7_U19 ( .B1(1'b1), .B2(SBOX_PL_7_n105), .A(SBOX_PL_7_n153), 
        .ZN(SBOX_PL_7_n81) );
  NAND2_X1 SBOX_PL_7_U18 ( .A1(1'b1), .A2(SBOX_Qreg6[15]), .ZN(SBOX_PL_7_n153)
         );
  OAI21_X1 SBOX_PL_7_U17 ( .B1(1'b1), .B2(SBOX_PL_7_n104), .A(SBOX_PL_7_n152), 
        .ZN(SBOX_PL_7_n80) );
  NAND2_X1 SBOX_PL_7_U16 ( .A1(1'b1), .A2(SBOX_Qreg6[16]), .ZN(SBOX_PL_7_n152)
         );
  OAI21_X1 SBOX_PL_7_U15 ( .B1(1'b1), .B2(SBOX_PL_7_n103), .A(SBOX_PL_7_n151), 
        .ZN(SBOX_PL_7_n79) );
  NAND2_X1 SBOX_PL_7_U14 ( .A1(1'b1), .A2(SBOX_Qreg6[17]), .ZN(SBOX_PL_7_n151)
         );
  OAI21_X1 SBOX_PL_7_U13 ( .B1(1'b1), .B2(SBOX_PL_7_n102), .A(SBOX_PL_7_n150), 
        .ZN(SBOX_PL_7_n78) );
  NAND2_X1 SBOX_PL_7_U12 ( .A1(1'b1), .A2(SBOX_Qreg6[18]), .ZN(SBOX_PL_7_n150)
         );
  OAI21_X1 SBOX_PL_7_U11 ( .B1(1'b1), .B2(SBOX_PL_7_n101), .A(SBOX_PL_7_n149), 
        .ZN(SBOX_PL_7_n77) );
  NAND2_X1 SBOX_PL_7_U10 ( .A1(1'b1), .A2(SBOX_Qreg6[19]), .ZN(SBOX_PL_7_n149)
         );
  OAI21_X1 SBOX_PL_7_U9 ( .B1(1'b1), .B2(SBOX_PL_7_n100), .A(SBOX_PL_7_n148), 
        .ZN(SBOX_PL_7_n76) );
  NAND2_X1 SBOX_PL_7_U8 ( .A1(1'b1), .A2(SBOX_Qreg6[20]), .ZN(SBOX_PL_7_n148)
         );
  OAI21_X1 SBOX_PL_7_U7 ( .B1(1'b1), .B2(SBOX_PL_7_n99), .A(SBOX_PL_7_n147), 
        .ZN(SBOX_PL_7_n75) );
  NAND2_X1 SBOX_PL_7_U6 ( .A1(1'b1), .A2(SBOX_Qreg6[21]), .ZN(SBOX_PL_7_n147)
         );
  OAI21_X1 SBOX_PL_7_U5 ( .B1(1'b1), .B2(SBOX_PL_7_n98), .A(SBOX_PL_7_n146), 
        .ZN(SBOX_PL_7_n74) );
  NAND2_X1 SBOX_PL_7_U4 ( .A1(1'b1), .A2(SBOX_Qreg6[22]), .ZN(SBOX_PL_7_n146)
         );
  OAI21_X1 SBOX_PL_7_U3 ( .B1(1'b1), .B2(SBOX_PL_7_n97), .A(SBOX_PL_7_n145), 
        .ZN(SBOX_PL_7_n73) );
  NAND2_X1 SBOX_PL_7_U2 ( .A1(1'b1), .A2(SBOX_Qreg6[23]), .ZN(SBOX_PL_7_n145)
         );
  DFF_X1 SBOX_PL_7_s_current_state_reg_0_ ( .D(SBOX_PL_7_n96), .CK(ClkxCI), 
        .Q(StateInxD[0]), .QN(SBOX_PL_7_n120) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_1_ ( .D(SBOX_PL_7_n95), .CK(ClkxCI), 
        .Q(StateInxD[1]), .QN(SBOX_PL_7_n119) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_2_ ( .D(SBOX_PL_7_n94), .CK(ClkxCI), 
        .Q(StateInxD[2]), .QN(SBOX_PL_7_n118) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_3_ ( .D(SBOX_PL_7_n93), .CK(ClkxCI), 
        .Q(StateInxD[3]), .QN(SBOX_PL_7_n117) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_4_ ( .D(SBOX_PL_7_n92), .CK(ClkxCI), 
        .Q(StateInxD[4]), .QN(SBOX_PL_7_n116) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_5_ ( .D(SBOX_PL_7_n91), .CK(ClkxCI), 
        .Q(StateInxD[5]), .QN(SBOX_PL_7_n115) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_6_ ( .D(SBOX_PL_7_n90), .CK(ClkxCI), 
        .Q(StateInxD[6]), .QN(SBOX_PL_7_n114) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_7_ ( .D(SBOX_PL_7_n89), .CK(ClkxCI), 
        .Q(StateInxD[7]), .QN(SBOX_PL_7_n113) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_8_ ( .D(SBOX_PL_7_n88), .CK(ClkxCI), 
        .Q(StateInxD[8]), .QN(SBOX_PL_7_n112) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_9_ ( .D(SBOX_PL_7_n87), .CK(ClkxCI), 
        .Q(StateInxD[9]), .QN(SBOX_PL_7_n111) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_10_ ( .D(SBOX_PL_7_n86), .CK(ClkxCI), 
        .Q(StateInxD[10]), .QN(SBOX_PL_7_n110) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_11_ ( .D(SBOX_PL_7_n85), .CK(ClkxCI), 
        .Q(StateInxD[11]), .QN(SBOX_PL_7_n109) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_12_ ( .D(SBOX_PL_7_n84), .CK(ClkxCI), 
        .Q(StateInxD[12]), .QN(SBOX_PL_7_n108) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_13_ ( .D(SBOX_PL_7_n83), .CK(ClkxCI), 
        .Q(StateInxD[13]), .QN(SBOX_PL_7_n107) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_14_ ( .D(SBOX_PL_7_n82), .CK(ClkxCI), 
        .Q(StateInxD[14]), .QN(SBOX_PL_7_n106) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_15_ ( .D(SBOX_PL_7_n81), .CK(ClkxCI), 
        .Q(StateInxD[15]), .QN(SBOX_PL_7_n105) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_16_ ( .D(SBOX_PL_7_n80), .CK(ClkxCI), 
        .Q(StateInxD[16]), .QN(SBOX_PL_7_n104) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_17_ ( .D(SBOX_PL_7_n79), .CK(ClkxCI), 
        .Q(StateInxD[17]), .QN(SBOX_PL_7_n103) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_18_ ( .D(SBOX_PL_7_n78), .CK(ClkxCI), 
        .Q(StateInxD[18]), .QN(SBOX_PL_7_n102) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_19_ ( .D(SBOX_PL_7_n77), .CK(ClkxCI), 
        .Q(StateInxD[19]), .QN(SBOX_PL_7_n101) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_20_ ( .D(SBOX_PL_7_n76), .CK(ClkxCI), 
        .Q(StateInxD[20]), .QN(SBOX_PL_7_n100) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_21_ ( .D(SBOX_PL_7_n75), .CK(ClkxCI), 
        .Q(StateInxD[21]), .QN(SBOX_PL_7_n99) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_22_ ( .D(SBOX_PL_7_n74), .CK(ClkxCI), 
        .Q(StateInxD[22]), .QN(SBOX_PL_7_n98) );
  DFF_X1 SBOX_PL_7_s_current_state_reg_23_ ( .D(SBOX_PL_7_n73), .CK(ClkxCI), 
        .Q(StateInxD[23]), .QN(SBOX_PL_7_n97) );
  BUF_X1 aes_key_regs_2_U3 ( .A(n170), .Z(aes_key_regs_2_n3) );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_0_ ( .D(aes_key_regs_2_K00xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[16]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_0_ ( .D(aes_key_regs_2_K10xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_0_ ( .D(aes_key_regs_2_K20xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_0_ ( .D(aes_key_regs_2_K01xDP_0_), .SI(
        KeyOutxD[16]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_2_K20xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_0_ ( .D(aes_key_regs_2_K01xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_0_ ( .D(aes_key_regs_2_K11xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_0_ ( .D(aes_key_regs_2_K21xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_0_ ( .D(aes_key_regs_2_K02xDP_0_), .SI(
        aes_key_regs_2_K01xDP_0_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K21xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_0_ ( .D(aes_key_regs_2_K02xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_0_ ( .D(aes_key_regs_2_K12xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_0_ ( .D(aes_key_regs_2_K22xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_0_ ( .D(K03xD[16]), .SI(
        aes_key_regs_2_K02xDP_0_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K22xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_1_ ( .D(aes_key_regs_2_K00xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[17]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_1_ ( .D(aes_key_regs_2_K10xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_1_ ( .D(aes_key_regs_2_K20xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_1_ ( .D(aes_key_regs_2_K01xDP_1_), .SI(
        KeyOutxD[17]), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K20xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_1_ ( .D(aes_key_regs_2_K01xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_1_ ( .D(aes_key_regs_2_K11xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_1_ ( .D(aes_key_regs_2_K21xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_1_ ( .D(aes_key_regs_2_K02xDP_1_), .SI(
        aes_key_regs_2_K01xDP_1_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K21xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_1_ ( .D(aes_key_regs_2_K02xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_1_ ( .D(aes_key_regs_2_K12xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_1_ ( .D(aes_key_regs_2_K22xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_1_ ( .D(K03xD[17]), .SI(
        aes_key_regs_2_K02xDP_1_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K22xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_2_ ( .D(aes_key_regs_2_K00xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[18]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_2_ ( .D(aes_key_regs_2_K10xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_2_ ( .D(aes_key_regs_2_K20xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_2_ ( .D(aes_key_regs_2_K01xDP_2_), .SI(
        KeyOutxD[18]), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K20xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_2_ ( .D(aes_key_regs_2_K01xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_2_ ( .D(aes_key_regs_2_K11xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_2_ ( .D(aes_key_regs_2_K21xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_2_ ( .D(aes_key_regs_2_K02xDP_2_), .SI(
        aes_key_regs_2_K01xDP_2_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K21xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_2_ ( .D(aes_key_regs_2_K02xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_2_ ( .D(aes_key_regs_2_K12xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_2_ ( .D(aes_key_regs_2_K22xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_2_ ( .D(K03xD[18]), .SI(
        aes_key_regs_2_K02xDP_2_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K22xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_3_ ( .D(aes_key_regs_2_K00xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[19]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_3_ ( .D(aes_key_regs_2_K10xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_3_ ( .D(aes_key_regs_2_K20xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_3_ ( .D(aes_key_regs_2_K01xDP_3_), .SI(
        KeyOutxD[19]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_2_K20xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_3_ ( .D(aes_key_regs_2_K01xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_3_ ( .D(aes_key_regs_2_K11xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_3_ ( .D(aes_key_regs_2_K21xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_3_ ( .D(aes_key_regs_2_K02xDP_3_), .SI(
        aes_key_regs_2_K01xDP_3_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K21xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_3_ ( .D(aes_key_regs_2_K02xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_3_ ( .D(aes_key_regs_2_K12xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_3_ ( .D(aes_key_regs_2_K22xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_3_ ( .D(K03xD[19]), .SI(
        aes_key_regs_2_K02xDP_3_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K22xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_4_ ( .D(aes_key_regs_2_K00xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[20]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_4_ ( .D(aes_key_regs_2_K10xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_4_ ( .D(aes_key_regs_2_K20xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_4_ ( .D(aes_key_regs_2_K01xDP_4_), .SI(
        KeyOutxD[20]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_2_K20xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_4_ ( .D(aes_key_regs_2_K01xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_4_ ( .D(aes_key_regs_2_K11xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_4_ ( .D(aes_key_regs_2_K21xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_4_ ( .D(aes_key_regs_2_K02xDP_4_), .SI(
        aes_key_regs_2_K01xDP_4_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K21xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_4_ ( .D(aes_key_regs_2_K02xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_4_ ( .D(aes_key_regs_2_K12xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_4_ ( .D(aes_key_regs_2_K22xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_4_ ( .D(K03xD[20]), .SI(
        aes_key_regs_2_K02xDP_4_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K22xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_5_ ( .D(aes_key_regs_2_K00xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[21]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_5_ ( .D(aes_key_regs_2_K10xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_5_ ( .D(aes_key_regs_2_K20xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_5_ ( .D(aes_key_regs_2_K01xDP_5_), .SI(
        KeyOutxD[21]), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K20xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_5_ ( .D(aes_key_regs_2_K01xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_5_ ( .D(aes_key_regs_2_K11xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_5_ ( .D(aes_key_regs_2_K21xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_5_ ( .D(aes_key_regs_2_K02xDP_5_), .SI(
        aes_key_regs_2_K01xDP_5_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K21xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_5_ ( .D(aes_key_regs_2_K02xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_5_ ( .D(aes_key_regs_2_K12xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_5_ ( .D(aes_key_regs_2_K22xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_5_ ( .D(K03xD[21]), .SI(
        aes_key_regs_2_K02xDP_5_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K22xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_6_ ( .D(aes_key_regs_2_K00xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[22]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_6_ ( .D(aes_key_regs_2_K10xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_6_ ( .D(aes_key_regs_2_K20xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_6_ ( .D(aes_key_regs_2_K01xDP_6_), .SI(
        KeyOutxD[22]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_2_K20xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_6_ ( .D(aes_key_regs_2_K01xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_6_ ( .D(aes_key_regs_2_K11xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_6_ ( .D(aes_key_regs_2_K21xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_6_ ( .D(aes_key_regs_2_K02xDP_6_), .SI(
        aes_key_regs_2_K01xDP_6_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K21xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_6_ ( .D(aes_key_regs_2_K02xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_6_ ( .D(aes_key_regs_2_K12xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_6_ ( .D(aes_key_regs_2_K22xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_6_ ( .D(K03xD[22]), .SI(
        aes_key_regs_2_K02xDP_6_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K22xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_2_K00xDP_reg_7_ ( .D(aes_key_regs_2_K00xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[23]), .QN() );
  DFFR_X1 aes_key_regs_2_K10xDP_reg_7_ ( .D(aes_key_regs_2_K10xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K00xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_2_K20xDP_reg_7_ ( .D(aes_key_regs_2_K20xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K10xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_2_K30xDP_reg_7_ ( .D(aes_key_regs_2_K01xDP_7_), .SI(
        KeyOutxD[23]), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K20xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_2_K01xDP_reg_7_ ( .D(aes_key_regs_2_K01xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_2_K11xDP_reg_7_ ( .D(aes_key_regs_2_K11xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K01xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_2_K21xDP_reg_7_ ( .D(aes_key_regs_2_K21xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K11xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_2_K31xDP_reg_7_ ( .D(aes_key_regs_2_K02xDP_7_), .SI(
        aes_key_regs_2_K01xDP_7_), .SE(aes_key_regs_2_n3), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_2_K21xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_2_K02xDP_reg_7_ ( .D(aes_key_regs_2_K02xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_2_K12xDP_reg_7_ ( .D(aes_key_regs_2_K12xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K02xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_2_K22xDP_reg_7_ ( .D(aes_key_regs_2_K22xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K12xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_2_K32xDP_reg_7_ ( .D(K03xD[23]), .SI(
        aes_key_regs_2_K02xDP_7_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_2_K22xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_0_ ( .D(KeyInxD[16]), .SI(K03xD[16]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[0]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_0_ ( .D(KeyToSboxOutxD[16]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[16]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_0_ ( .D(aes_key_regs_2_K13xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[16]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_0_ ( .D(aes_key_regs_2_K23xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_1_ ( .D(KeyInxD[17]), .SI(K03xD[17]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[1]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_1_ ( .D(KeyToSboxOutxD[17]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[17]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_1_ ( .D(aes_key_regs_2_K13xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[17]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_1_ ( .D(aes_key_regs_2_K23xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_2_ ( .D(KeyInxD[18]), .SI(K03xD[18]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[2]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_2_ ( .D(KeyToSboxOutxD[18]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[18]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_2_ ( .D(aes_key_regs_2_K13xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[18]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_2_ ( .D(aes_key_regs_2_K23xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_3_ ( .D(KeyInxD[19]), .SI(K03xD[19]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[3]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_3_ ( .D(KeyToSboxOutxD[19]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[19]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_3_ ( .D(aes_key_regs_2_K13xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[19]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_3_ ( .D(aes_key_regs_2_K23xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_4_ ( .D(KeyInxD[20]), .SI(K03xD[20]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[4]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_4_ ( .D(KeyToSboxOutxD[20]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[20]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_4_ ( .D(aes_key_regs_2_K13xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[20]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_4_ ( .D(aes_key_regs_2_K23xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_5_ ( .D(KeyInxD[21]), .SI(K03xD[21]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[5]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_5_ ( .D(KeyToSboxOutxD[21]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[21]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_5_ ( .D(aes_key_regs_2_K13xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[21]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_5_ ( .D(aes_key_regs_2_K23xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_6_ ( .D(KeyInxD[22]), .SI(K03xD[22]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[6]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_6_ ( .D(KeyToSboxOutxD[22]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[22]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_6_ ( .D(aes_key_regs_2_K13xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[22]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_6_ ( .D(aes_key_regs_2_K23xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_2_K33xDP_reg_7_ ( .D(KeyInxD[23]), .SI(K03xD[23]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K23xDN[7]), 
        .QN() );
  DFFR_X1 aes_key_regs_2_K03xDP_reg_7_ ( .D(KeyToSboxOutxD[23]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[23]), .QN() );
  DFFR_X1 aes_key_regs_2_K13xDP_reg_7_ ( .D(aes_key_regs_2_K13xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[23]), .QN() );
  DFFR_X1 aes_key_regs_2_K23xDP_reg_7_ ( .D(aes_key_regs_2_K23xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_2_K13xDN[7]), .QN() );
  OAI222_X1 aes_state_regs_2_U60 ( .A1(aes_state_regs_2_n117), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n118), .B2(
        aes_state_regs_2_n98), .C1(aes_state_regs_2_n114), .C2(
        aes_state_regs_2_n47), .ZN(aes_state_regs_2_S10xDN[7]) );
  INV_X1 aes_state_regs_2_U59 ( .A(aes_state_regs_2_MixColumnsS2xD[7]), .ZN(
        aes_state_regs_2_n117) );
  OAI222_X1 aes_state_regs_2_U58 ( .A1(aes_state_regs_2_n116), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n118), .B2(
        aes_state_regs_2_n99), .C1(aes_state_regs_2_n114), .C2(
        aes_state_regs_2_n48), .ZN(aes_state_regs_2_S10xDN[6]) );
  INV_X1 aes_state_regs_2_U57 ( .A(aes_state_regs_2_MixColumnsS2xD[6]), .ZN(
        aes_state_regs_2_n116) );
  OAI222_X1 aes_state_regs_2_U56 ( .A1(aes_state_regs_2_n115), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n118), .B2(
        aes_state_regs_2_n100), .C1(aes_state_regs_2_n114), .C2(
        aes_state_regs_2_n49), .ZN(aes_state_regs_2_S10xDN[5]) );
  INV_X1 aes_state_regs_2_U55 ( .A(aes_state_regs_2_MixColumnsS2xD[5]), .ZN(
        aes_state_regs_2_n115) );
  NAND2_X1 aes_state_regs_2_U54 ( .A1(doMixColumnsxS), .A2(
        aes_state_regs_2_n114), .ZN(aes_state_regs_2_n66) );
  INV_X1 aes_state_regs_2_U53 ( .A(aes_state_regs_2_n114), .ZN(
        aes_state_regs_2_n112) );
  INV_X1 aes_state_regs_2_U52 ( .A(aes_state_regs_2_n114), .ZN(
        aes_state_regs_2_n111) );
  INV_X1 aes_state_regs_2_U51 ( .A(aes_state_regs_2_n114), .ZN(
        aes_state_regs_2_n110) );
  INV_X1 aes_state_regs_2_U50 ( .A(aes_state_regs_2_n114), .ZN(
        aes_state_regs_2_n113) );
  BUF_X2 aes_state_regs_2_U49 ( .A(aes_state_regs_2_n66), .Z(
        aes_state_regs_2_n107) );
  INV_X1 aes_state_regs_2_U48 ( .A(n453), .ZN(aes_state_regs_2_n114) );
  INV_X1 aes_state_regs_2_U47 ( .A(aes_state_regs_2_n107), .ZN(
        aes_state_regs_2_n108) );
  OAI21_X1 aes_state_regs_2_U46 ( .B1(aes_state_regs_2_n91), .B2(
        aes_state_regs_2_n118), .A(aes_state_regs_2_n81), .ZN(
        aes_state_regs_2_S20xDN[6]) );
  AOI22_X1 aes_state_regs_2_U45 ( .A1(aes_state_regs_2_MixColumnsS3xD[6]), 
        .A2(aes_state_regs_2_n109), .B1(aes_state_regs_2_n8), .B2(
        aes_state_regs_2_n113), .ZN(aes_state_regs_2_n81) );
  OAI21_X1 aes_state_regs_2_U44 ( .B1(aes_state_regs_2_n109), .B2(
        aes_state_regs_2_n86), .A(aes_state_regs_2_n80), .ZN(StateOutxD[18])
         );
  NAND2_X1 aes_state_regs_2_U43 ( .A1(aes_state_regs_2_n109), .A2(
        aes_state_regs_2_MixColumnsS0xD[2]), .ZN(aes_state_regs_2_n80) );
  OAI21_X1 aes_state_regs_2_U42 ( .B1(aes_state_regs_2_n108), .B2(
        aes_state_regs_2_n87), .A(aes_state_regs_2_n79), .ZN(StateOutxD[19])
         );
  NAND2_X1 aes_state_regs_2_U41 ( .A1(aes_state_regs_2_MixColumnsS0xD[3]), 
        .A2(aes_state_regs_2_n109), .ZN(aes_state_regs_2_n79) );
  OAI222_X1 aes_state_regs_2_U40 ( .A1(aes_state_regs_2_n78), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n62), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n97), .ZN(aes_state_regs_2_S20xDN[0]) );
  INV_X1 aes_state_regs_2_U39 ( .A(aes_state_regs_2_MixColumnsS3xD[0]), .ZN(
        aes_state_regs_2_n78) );
  OAI21_X1 aes_state_regs_2_U38 ( .B1(aes_state_regs_2_n109), .B2(
        aes_state_regs_2_n83), .A(aes_state_regs_2_n77), .ZN(StateOutxD[22])
         );
  NAND2_X1 aes_state_regs_2_U37 ( .A1(aes_state_regs_2_MixColumnsS0xD[6]), 
        .A2(aes_state_regs_2_n108), .ZN(aes_state_regs_2_n77) );
  OAI222_X1 aes_state_regs_2_U36 ( .A1(aes_state_regs_2_n76), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n54), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n105), .ZN(aes_state_regs_2_S10xDN[0]) );
  INV_X1 aes_state_regs_2_U35 ( .A(aes_state_regs_2_MixColumnsS2xD[0]), .ZN(
        aes_state_regs_2_n76) );
  OAI21_X1 aes_state_regs_2_U34 ( .B1(aes_state_regs_2_n108), .B2(
        aes_state_regs_2_n88), .A(aes_state_regs_2_n75), .ZN(StateOutxD[20])
         );
  NAND2_X1 aes_state_regs_2_U33 ( .A1(aes_state_regs_2_MixColumnsS0xD[4]), 
        .A2(aes_state_regs_2_n109), .ZN(aes_state_regs_2_n75) );
  OAI222_X1 aes_state_regs_2_U32 ( .A1(aes_state_regs_2_n74), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n59), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n94), .ZN(aes_state_regs_2_S20xDN[3]) );
  INV_X1 aes_state_regs_2_U31 ( .A(aes_state_regs_2_MixColumnsS3xD[3]), .ZN(
        aes_state_regs_2_n74) );
  OAI21_X1 aes_state_regs_2_U30 ( .B1(aes_state_regs_2_n108), .B2(
        aes_state_regs_2_n89), .A(aes_state_regs_2_n73), .ZN(StateOutxD[21])
         );
  NAND2_X1 aes_state_regs_2_U29 ( .A1(aes_state_regs_2_n108), .A2(
        aes_state_regs_2_MixColumnsS0xD[5]), .ZN(aes_state_regs_2_n73) );
  OAI222_X1 aes_state_regs_2_U28 ( .A1(aes_state_regs_2_n72), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n61), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n96), .ZN(aes_state_regs_2_S20xDN[1]) );
  INV_X1 aes_state_regs_2_U27 ( .A(aes_state_regs_2_MixColumnsS3xD[1]), .ZN(
        aes_state_regs_2_n72) );
  OAI222_X1 aes_state_regs_2_U26 ( .A1(aes_state_regs_2_n71), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n60), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n95), .ZN(aes_state_regs_2_S20xDN[2]) );
  INV_X1 aes_state_regs_2_U25 ( .A(aes_state_regs_2_MixColumnsS3xD[2]), .ZN(
        aes_state_regs_2_n71) );
  OAI21_X1 aes_state_regs_2_U24 ( .B1(aes_state_regs_2_n109), .B2(
        aes_state_regs_2_n84), .A(aes_state_regs_2_n70), .ZN(StateOutxD[23])
         );
  NAND2_X1 aes_state_regs_2_U23 ( .A1(aes_state_regs_2_n109), .A2(
        aes_state_regs_2_MixColumnsS0xD[7]), .ZN(aes_state_regs_2_n70) );
  OAI222_X1 aes_state_regs_2_U22 ( .A1(aes_state_regs_2_n69), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n58), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n93), .ZN(aes_state_regs_2_S20xDN[4]) );
  INV_X1 aes_state_regs_2_U21 ( .A(aes_state_regs_2_MixColumnsS3xD[4]), .ZN(
        aes_state_regs_2_n69) );
  OAI222_X1 aes_state_regs_2_U20 ( .A1(aes_state_regs_2_n68), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n57), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n92), .ZN(aes_state_regs_2_S20xDN[5]) );
  INV_X1 aes_state_regs_2_U19 ( .A(aes_state_regs_2_MixColumnsS3xD[5]), .ZN(
        aes_state_regs_2_n68) );
  OAI222_X1 aes_state_regs_2_U18 ( .A1(aes_state_regs_2_n67), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n55), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n90), .ZN(aes_state_regs_2_S20xDN[7]) );
  INV_X1 aes_state_regs_2_U17 ( .A(aes_state_regs_2_MixColumnsS3xD[7]), .ZN(
        aes_state_regs_2_n67) );
  OAI222_X1 aes_state_regs_2_U16 ( .A1(aes_state_regs_2_n65), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n53), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n104), .ZN(aes_state_regs_2_S10xDN[1]) );
  INV_X1 aes_state_regs_2_U15 ( .A(aes_state_regs_2_MixColumnsS2xD[1]), .ZN(
        aes_state_regs_2_n65) );
  OAI222_X1 aes_state_regs_2_U14 ( .A1(aes_state_regs_2_n64), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n52), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n103), .ZN(aes_state_regs_2_S10xDN[2]) );
  INV_X1 aes_state_regs_2_U13 ( .A(aes_state_regs_2_MixColumnsS2xD[2]), .ZN(
        aes_state_regs_2_n64) );
  OAI222_X1 aes_state_regs_2_U12 ( .A1(aes_state_regs_2_n63), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n51), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n102), .ZN(aes_state_regs_2_S10xDN[3]) );
  INV_X1 aes_state_regs_2_U11 ( .A(aes_state_regs_2_MixColumnsS2xD[3]), .ZN(
        aes_state_regs_2_n63) );
  OAI21_X1 aes_state_regs_2_U10 ( .B1(aes_state_regs_2_n109), .B2(
        aes_state_regs_2_n85), .A(aes_state_regs_2_n56), .ZN(StateOutxD[17])
         );
  NAND2_X1 aes_state_regs_2_U9 ( .A1(aes_state_regs_2_n109), .A2(
        aes_state_regs_2_MixColumnsS0xD[1]), .ZN(aes_state_regs_2_n56) );
  OAI222_X1 aes_state_regs_2_U8 ( .A1(aes_state_regs_2_n46), .A2(
        aes_state_regs_2_n107), .B1(aes_state_regs_2_n114), .B2(
        aes_state_regs_2_n50), .C1(aes_state_regs_2_n118), .C2(
        aes_state_regs_2_n101), .ZN(aes_state_regs_2_S10xDN[4]) );
  INV_X1 aes_state_regs_2_U7 ( .A(aes_state_regs_2_MixColumnsS2xD[4]), .ZN(
        aes_state_regs_2_n46) );
  OAI21_X1 aes_state_regs_2_U6 ( .B1(aes_state_regs_2_n108), .B2(
        aes_state_regs_2_n82), .A(aes_state_regs_2_n45), .ZN(StateOutxD[16])
         );
  NAND2_X1 aes_state_regs_2_U5 ( .A1(aes_state_regs_2_n108), .A2(
        aes_state_regs_2_MixColumnsS0xD[0]), .ZN(aes_state_regs_2_n45) );
  OR2_X1 aes_state_regs_2_U4 ( .A1(aes_state_regs_2_n113), .A2(doMixColumnsxS), 
        .ZN(aes_state_regs_2_n118) );
  INV_X1 aes_state_regs_2_U3 ( .A(aes_state_regs_2_n107), .ZN(
        aes_state_regs_2_n109) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_7_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[7]), .SI(aes_state_regs_2_S10xDP_7_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[7]), .QN(aes_state_regs_2_n84) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_6_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[6]), .SI(aes_state_regs_2_S10xDP_6_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[6]), .QN(aes_state_regs_2_n83) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_5_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[5]), .SI(aes_state_regs_2_S10xDP_5_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[5]), .QN(aes_state_regs_2_n89) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_4_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[4]), .SI(aes_state_regs_2_S10xDP_4_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[4]), .QN(aes_state_regs_2_n88) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_3_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[3]), .SI(aes_state_regs_2_S10xDP_3_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[3]), .QN(aes_state_regs_2_n87) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_2_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[2]), .SI(aes_state_regs_2_S10xDP_2_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[2]), .QN(aes_state_regs_2_n86) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_1_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[1]), .SI(aes_state_regs_2_S10xDP_1_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[1]), .QN(aes_state_regs_2_n85) );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_7_ ( .D(aes_state_regs_2_S10xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_7_), .QN() );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_6_ ( .D(aes_state_regs_2_S10xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_6_), .QN() );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_5_ ( .D(aes_state_regs_2_S10xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_5_), .QN() );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_4_ ( .D(aes_state_regs_2_S10xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_4_), .QN() );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_3_ ( .D(aes_state_regs_2_S10xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_3_), .QN() );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_2_ ( .D(aes_state_regs_2_S10xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_2_), .QN() );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_1_ ( .D(aes_state_regs_2_S10xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_7_ ( .D(aes_state_regs_2_S01xDO_7_), 
        .SI(StateInxD[23]), .SE(aes_state_regs_2_n111), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_7_), .QN(aes_state_regs_2_n90) );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_7_ ( .D(aes_state_regs_2_n1), .SI(
        aes_state_regs_2_n4), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S21xDP[7]), .QN(aes_state_regs_2_n47) );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_7_ ( .D(aes_state_regs_2_S02xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_7_ ( .D(aes_state_regs_2_n2), .SI(
        aes_state_regs_2_S23xDP_7_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_7_ ( .D(aes_state_regs_2_n4), .SI(
        aes_state_regs_2_n1), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S23xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_7_ ( .D(aes_state_regs_2_S02xDP_7_), 
        .SI(aes_state_regs_2_S01xDO_7_), .SE(aes_state_regs_2_n112), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n1), .QN() );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_7_ ( .D(aes_state_regs_2_S01xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_7_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_7_ ( .D(aes_state_regs_2_S21xDP[7]), 
        .SI(aes_state_regs_2_n2), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_7_ ( .D(aes_state_regs_2_n3), .SI(
        aes_state_regs_2_S30xDP_7_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n2), .QN() );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_7_ ( .D(aes_state_regs_2_n5), .SI(
        aes_state_regs_2_S02xDP_7_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n3), .QN(aes_state_regs_2_n55) );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_7_ ( .D(StateInxD[23]), .SI(
        aes_state_regs_2_n5), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_n4), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_7_ ( .D(aes_state_regs_2_S03xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n5), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_7_ ( .D(aes_state_regs_2_S23xDP_7_), 
        .SI(aes_state_regs_2_S20xDP_7_), .SE(aes_state_regs_2_n110), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[7]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_7_ ( .D(aes_state_regs_2_S20xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_7_), .QN(
        aes_state_regs_2_n98) );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_6_ ( .D(aes_state_regs_2_S01xDO_6_), 
        .SI(StateInxD[22]), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_6_), .QN(aes_state_regs_2_n91) );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_6_ ( .D(aes_state_regs_2_n6), .SI(
        aes_state_regs_2_n9), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S21xDP[6]), .QN(aes_state_regs_2_n48) );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_6_ ( .D(aes_state_regs_2_S02xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_6_ ( .D(aes_state_regs_2_n7), .SI(
        aes_state_regs_2_S23xDP_6_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_6_ ( .D(aes_state_regs_2_n9), .SI(
        aes_state_regs_2_n6), .SE(aes_state_regs_2_n111), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S23xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_6_ ( .D(aes_state_regs_2_S02xDP_6_), 
        .SI(aes_state_regs_2_S01xDO_6_), .SE(aes_state_regs_2_n111), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n6), .QN() );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_6_ ( .D(aes_state_regs_2_S01xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_6_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_6_ ( .D(aes_state_regs_2_S21xDP[6]), 
        .SI(aes_state_regs_2_n7), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_6_ ( .D(aes_state_regs_2_n8), .SI(
        aes_state_regs_2_S30xDP_6_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n7), .QN() );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_6_ ( .D(aes_state_regs_2_n10), .SI(
        aes_state_regs_2_S02xDP_6_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n8), .QN() );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_6_ ( .D(StateInxD[22]), .SI(
        aes_state_regs_2_n10), .SE(aes_state_regs_2_n111), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_n9), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_6_ ( .D(aes_state_regs_2_S03xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n10), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_6_ ( .D(aes_state_regs_2_S23xDP_6_), 
        .SI(aes_state_regs_2_S20xDP_6_), .SE(aes_state_regs_2_n112), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[6]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_6_ ( .D(aes_state_regs_2_S20xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_6_), .QN(
        aes_state_regs_2_n99) );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_5_ ( .D(aes_state_regs_2_S01xDO_5_), 
        .SI(StateInxD[21]), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_5_), .QN(aes_state_regs_2_n92) );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_5_ ( .D(aes_state_regs_2_n11), .SI(
        aes_state_regs_2_n14), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S21xDP[5]), .QN(aes_state_regs_2_n49) );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_5_ ( .D(aes_state_regs_2_S02xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_5_ ( .D(aes_state_regs_2_n12), .SI(
        aes_state_regs_2_S23xDP_5_), .SE(aes_state_regs_2_n112), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_5_ ( .D(aes_state_regs_2_n14), .SI(
        aes_state_regs_2_n11), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S23xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_5_ ( .D(aes_state_regs_2_S02xDP_5_), 
        .SI(aes_state_regs_2_S01xDO_5_), .SE(aes_state_regs_2_n111), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n11), .QN() );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_5_ ( .D(aes_state_regs_2_S01xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_5_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_5_ ( .D(aes_state_regs_2_S21xDP[5]), 
        .SI(aes_state_regs_2_n12), .SE(aes_state_regs_2_n112), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_5_ ( .D(aes_state_regs_2_n13), .SI(
        aes_state_regs_2_S30xDP_5_), .SE(aes_state_regs_2_n112), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n12), .QN() );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_5_ ( .D(aes_state_regs_2_n15), .SI(
        aes_state_regs_2_S02xDP_5_), .SE(aes_state_regs_2_n112), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n13), .QN(aes_state_regs_2_n57) );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_5_ ( .D(StateInxD[21]), .SI(
        aes_state_regs_2_n15), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_n14), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_5_ ( .D(aes_state_regs_2_S03xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n15), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_5_ ( .D(aes_state_regs_2_S23xDP_5_), 
        .SI(aes_state_regs_2_S20xDP_5_), .SE(aes_state_regs_2_n112), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[5]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_5_ ( .D(aes_state_regs_2_S20xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_5_), .QN(
        aes_state_regs_2_n100) );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_4_ ( .D(aes_state_regs_2_S01xDO_4_), 
        .SI(StateInxD[20]), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_4_), .QN(aes_state_regs_2_n93) );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_4_ ( .D(aes_state_regs_2_n16), .SI(
        aes_state_regs_2_n19), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S21xDP[4]), .QN(aes_state_regs_2_n50) );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_4_ ( .D(aes_state_regs_2_S02xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_4_ ( .D(aes_state_regs_2_n17), .SI(
        aes_state_regs_2_S23xDP_4_), .SE(aes_state_regs_2_n112), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_4_ ( .D(aes_state_regs_2_n19), .SI(
        aes_state_regs_2_n16), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S23xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_4_ ( .D(aes_state_regs_2_S02xDP_4_), 
        .SI(aes_state_regs_2_S01xDO_4_), .SE(aes_state_regs_2_n111), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n16), .QN() );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_4_ ( .D(aes_state_regs_2_S01xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_4_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_4_ ( .D(aes_state_regs_2_S21xDP[4]), 
        .SI(aes_state_regs_2_n17), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_4_ ( .D(aes_state_regs_2_n18), .SI(
        aes_state_regs_2_S30xDP_4_), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n17), .QN() );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_4_ ( .D(aes_state_regs_2_n20), .SI(
        aes_state_regs_2_S02xDP_4_), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n18), .QN(aes_state_regs_2_n58) );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_4_ ( .D(StateInxD[20]), .SI(
        aes_state_regs_2_n20), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_n19), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_4_ ( .D(aes_state_regs_2_S03xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n20), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_4_ ( .D(aes_state_regs_2_S23xDP_4_), 
        .SI(aes_state_regs_2_S20xDP_4_), .SE(aes_state_regs_2_n111), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[4]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_4_ ( .D(aes_state_regs_2_S20xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_4_), .QN(
        aes_state_regs_2_n101) );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_3_ ( .D(aes_state_regs_2_S01xDO_3_), 
        .SI(StateInxD[19]), .SE(aes_state_regs_2_n111), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_3_), .QN(aes_state_regs_2_n94) );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_3_ ( .D(aes_state_regs_2_n21), .SI(
        aes_state_regs_2_n24), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S21xDP[3]), .QN(aes_state_regs_2_n51) );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_3_ ( .D(aes_state_regs_2_S02xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_3_ ( .D(aes_state_regs_2_n22), .SI(
        aes_state_regs_2_S23xDP_3_), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_3_ ( .D(aes_state_regs_2_n24), .SI(
        aes_state_regs_2_n21), .SE(aes_state_regs_2_n111), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S23xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_3_ ( .D(aes_state_regs_2_S02xDP_3_), 
        .SI(aes_state_regs_2_S01xDO_3_), .SE(aes_state_regs_2_n111), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n21), .QN() );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_3_ ( .D(aes_state_regs_2_S01xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_3_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_3_ ( .D(aes_state_regs_2_S21xDP[3]), 
        .SI(aes_state_regs_2_n22), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_3_ ( .D(aes_state_regs_2_n23), .SI(
        aes_state_regs_2_S30xDP_3_), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n22), .QN() );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_3_ ( .D(aes_state_regs_2_n25), .SI(
        aes_state_regs_2_S02xDP_3_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n23), .QN(aes_state_regs_2_n59) );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_3_ ( .D(StateInxD[19]), .SI(
        aes_state_regs_2_n25), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_n24), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_3_ ( .D(aes_state_regs_2_S03xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n25), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_3_ ( .D(aes_state_regs_2_S23xDP_3_), 
        .SI(aes_state_regs_2_S20xDP_3_), .SE(aes_state_regs_2_n111), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[3]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_3_ ( .D(aes_state_regs_2_S20xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_3_), .QN(
        aes_state_regs_2_n102) );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_2_ ( .D(aes_state_regs_2_S01xDO_2_), 
        .SI(StateInxD[18]), .SE(aes_state_regs_2_n113), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_2_), .QN(aes_state_regs_2_n95) );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_2_ ( .D(aes_state_regs_2_n26), .SI(
        aes_state_regs_2_n29), .SE(aes_state_regs_2_n113), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S21xDP[2]), .QN(aes_state_regs_2_n52) );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_2_ ( .D(aes_state_regs_2_S02xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_2_ ( .D(aes_state_regs_2_n27), .SI(
        aes_state_regs_2_S23xDP_2_), .SE(aes_state_regs_2_n113), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_2_ ( .D(aes_state_regs_2_n29), .SI(
        aes_state_regs_2_n26), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S23xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_2_ ( .D(aes_state_regs_2_S02xDP_2_), 
        .SI(aes_state_regs_2_S01xDO_2_), .SE(aes_state_regs_2_n111), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n26), .QN() );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_2_ ( .D(aes_state_regs_2_S01xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_2_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_2_ ( .D(aes_state_regs_2_S21xDP[2]), 
        .SI(aes_state_regs_2_n27), .SE(aes_state_regs_2_n113), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_2_ ( .D(aes_state_regs_2_n28), .SI(
        aes_state_regs_2_S30xDP_2_), .SE(aes_state_regs_2_n112), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n27), .QN() );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_2_ ( .D(aes_state_regs_2_n30), .SI(
        aes_state_regs_2_S02xDP_2_), .SE(aes_state_regs_2_n113), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n28), .QN(aes_state_regs_2_n60) );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_2_ ( .D(StateInxD[18]), .SI(
        aes_state_regs_2_n30), .SE(aes_state_regs_2_n110), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_n29), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_2_ ( .D(aes_state_regs_2_S03xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n30), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_2_ ( .D(aes_state_regs_2_S23xDP_2_), 
        .SI(aes_state_regs_2_S20xDP_2_), .SE(aes_state_regs_2_n113), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[2]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_2_ ( .D(aes_state_regs_2_S20xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_2_), .QN(
        aes_state_regs_2_n103) );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_1_ ( .D(aes_state_regs_2_S01xDO_1_), 
        .SI(StateInxD[17]), .SE(aes_state_regs_2_n113), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_1_), .QN(aes_state_regs_2_n96) );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_1_ ( .D(aes_state_regs_2_n31), .SI(
        aes_state_regs_2_n34), .SE(aes_state_regs_2_n113), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S21xDP[1]), .QN(aes_state_regs_2_n53) );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_1_ ( .D(aes_state_regs_2_S02xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_1_ ( .D(aes_state_regs_2_n32), .SI(
        aes_state_regs_2_S23xDP_1_), .SE(aes_state_regs_2_n113), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_1_ ( .D(aes_state_regs_2_n34), .SI(
        aes_state_regs_2_n31), .SE(aes_state_regs_2_n111), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S23xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_1_ ( .D(aes_state_regs_2_S02xDP_1_), 
        .SI(aes_state_regs_2_S01xDO_1_), .SE(aes_state_regs_2_n112), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n31), .QN() );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_1_ ( .D(aes_state_regs_2_S01xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_1_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_1_ ( .D(aes_state_regs_2_S21xDP[1]), 
        .SI(aes_state_regs_2_n32), .SE(aes_state_regs_2_n113), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_1_ ( .D(aes_state_regs_2_n33), .SI(
        aes_state_regs_2_S30xDP_1_), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n32), .QN() );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_1_ ( .D(aes_state_regs_2_n35), .SI(
        aes_state_regs_2_S02xDP_1_), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n33), .QN(aes_state_regs_2_n61) );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_1_ ( .D(StateInxD[17]), .SI(
        aes_state_regs_2_n35), .SE(aes_state_regs_2_n112), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_n34), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_1_ ( .D(aes_state_regs_2_S03xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n35), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_1_ ( .D(aes_state_regs_2_S23xDP_1_), 
        .SI(aes_state_regs_2_S20xDP_1_), .SE(aes_state_regs_2_n112), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[1]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_1_ ( .D(aes_state_regs_2_S20xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_1_), .QN(
        aes_state_regs_2_n104) );
  SDFFR_X1 aes_state_regs_2_S00xDP_reg_0_ ( .D(
        aes_state_regs_2_MixColumnsS1xD[0]), .SI(aes_state_regs_2_S10xDP_0_), 
        .SE(aes_state_regs_2_n107), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_2_S00xDP[0]), .QN(aes_state_regs_2_n82) );
  DFFR_X1 aes_state_regs_2_S10xDP_reg_0_ ( .D(aes_state_regs_2_S10xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S10xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_2_S23xDP_reg_0_ ( .D(aes_state_regs_2_n37), .SI(
        aes_state_regs_2_S31xDP_0_), .SE(aes_state_regs_2_n112), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S23xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_2_S31xDP_reg_0_ ( .D(aes_state_regs_2_S02xDP_0_), 
        .SI(aes_state_regs_2_S01xDO_0_), .SE(aes_state_regs_2_n112), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S31xDP_0_), .QN() );
  DFFR_X1 aes_state_regs_2_S02xDP_reg_0_ ( .D(aes_state_regs_2_S02xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_2_S12xDP_reg_0_ ( .D(aes_state_regs_2_S22xDP_0_), 
        .SI(aes_state_regs_2_S23xDP_0_), .SE(aes_state_regs_2_n113), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S02xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_2_S22xDP_reg_0_ ( .D(aes_state_regs_2_n38), .SI(
        aes_state_regs_2_S30xDP_0_), .SE(aes_state_regs_2_n113), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S22xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_2_S30xDP_reg_0_ ( .D(aes_state_regs_2_S01xDO_0_), 
        .SI(StateInxD[16]), .SE(aes_state_regs_2_n113), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_2_S30xDP_0_), .QN(aes_state_regs_2_n97) );
  DFFR_X1 aes_state_regs_2_S01xDP_reg_0_ ( .D(aes_state_regs_2_S01xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S01xDO_0_), .QN() );
  SDFFR_X1 aes_state_regs_2_S11xDP_reg_0_ ( .D(aes_state_regs_2_n36), .SI(
        aes_state_regs_2_S22xDP_0_), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_S01xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_2_S21xDP_reg_0_ ( .D(aes_state_regs_2_S31xDP_0_), 
        .SI(aes_state_regs_2_n37), .SE(aes_state_regs_2_n110), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n36), .QN(aes_state_regs_2_n54) );
  SDFFR_X1 aes_state_regs_2_S33xDP_reg_0_ ( .D(StateInxD[16]), .SI(
        aes_state_regs_2_S03xDP_0_), .SE(aes_state_regs_2_n111), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_2_n37), .QN() );
  DFFR_X1 aes_state_regs_2_S03xDP_reg_0_ ( .D(aes_state_regs_2_S03xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_2_S13xDP_reg_0_ ( .D(aes_state_regs_2_S23xDP_0_), 
        .SI(aes_state_regs_2_S20xDP_0_), .SE(aes_state_regs_2_n112), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S03xDN[0]), .QN() );
  DFFR_X1 aes_state_regs_2_S20xDP_reg_0_ ( .D(aes_state_regs_2_S20xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_S20xDP_0_), .QN(
        aes_state_regs_2_n105) );
  SDFFR_X1 aes_state_regs_2_S32xDP_reg_0_ ( .D(aes_state_regs_2_S03xDP_0_), 
        .SI(aes_state_regs_2_S02xDP_0_), .SE(aes_state_regs_2_n113), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_2_n38), .QN(
        aes_state_regs_2_n62) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U119 ( .A(
        aes_state_regs_2_mix_columns_1_n210), .B(
        aes_state_regs_2_mix_columns_1_n209), .ZN(
        aes_state_regs_2_mix_columns_1_n218) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U118 ( .A(
        aes_state_regs_2_mix_columns_1_n203), .B(
        aes_state_regs_2_mix_columns_1_n244), .ZN(
        aes_state_regs_2_MixColumnsS1xD[0]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U117 ( .A(
        aes_state_regs_2_mix_columns_1_n205), .B(aes_state_regs_2_S00xDP[0]), 
        .ZN(aes_state_regs_2_mix_columns_1_n203) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U116 ( .A(
        aes_state_regs_2_mix_columns_1_n202), .B(
        aes_state_regs_2_mix_columns_1_n201), .ZN(
        aes_state_regs_2_MixColumnsS3xD[6]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U115 ( .A(aes_state_regs_2_S30xDP_5_), .B(aes_state_regs_2_S00xDP[5]), .ZN(aes_state_regs_2_mix_columns_1_n202) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U114 ( .A1(
        aes_state_regs_2_mix_columns_1_n243), .A2(aes_state_regs_2_S20xDP_6_), 
        .B1(aes_state_regs_2_mix_columns_1_n242), .B2(
        aes_state_regs_2_mix_columns_1_n200), .ZN(
        aes_state_regs_2_mix_columns_1_n201) );
  INV_X1 aes_state_regs_2_mix_columns_1_U113 ( .A(
        aes_state_regs_2_mix_columns_1_n243), .ZN(
        aes_state_regs_2_mix_columns_1_n200) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U112 ( .A(
        aes_state_regs_2_mix_columns_1_n198), .B(
        aes_state_regs_2_mix_columns_1_n199), .ZN(
        aes_state_regs_2_MixColumnsS1xD[2]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U111 ( .A(aes_state_regs_2_S20xDP_1_), .B(aes_state_regs_2_S20xDP_2_), .ZN(aes_state_regs_2_mix_columns_1_n199) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U110 ( .A(
        aes_state_regs_2_mix_columns_1_n216), .B(aes_state_regs_2_S10xDP_1_), 
        .Z(aes_state_regs_2_mix_columns_1_n198) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U109 ( .A(
        aes_state_regs_2_mix_columns_1_n197), .B(
        aes_state_regs_2_mix_columns_1_n213), .ZN(
        aes_state_regs_2_MixColumnsS1xD[1]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U108 ( .A(
        aes_state_regs_2_mix_columns_1_n206), .B(aes_state_regs_2_S00xDP[1]), 
        .ZN(aes_state_regs_2_mix_columns_1_n197) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U107 ( .A(
        aes_state_regs_2_mix_columns_1_n196), .B(
        aes_state_regs_2_mix_columns_1_n218), .ZN(
        aes_state_regs_2_MixColumnsS1xD[3]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U106 ( .A(aes_state_regs_2_S20xDP_3_), .B(aes_state_regs_2_mix_columns_1_n207), .ZN(
        aes_state_regs_2_mix_columns_1_n196) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U105 ( .A(
        aes_state_regs_2_mix_columns_1_n194), .B(
        aes_state_regs_2_mix_columns_1_n195), .ZN(
        aes_state_regs_2_MixColumnsS1xD[5]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U104 ( .A(aes_state_regs_2_S20xDP_4_), .B(aes_state_regs_2_mix_columns_1_n225), .ZN(
        aes_state_regs_2_mix_columns_1_n195) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U103 ( .A(aes_state_regs_2_S00xDP[5]), 
        .B(aes_state_regs_2_S10xDP_4_), .Z(aes_state_regs_2_mix_columns_1_n194) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U102 ( .A(
        aes_state_regs_2_mix_columns_1_n193), .B(
        aes_state_regs_2_mix_columns_1_n220), .ZN(
        aes_state_regs_2_MixColumnsS1xD[4]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U101 ( .A(
        aes_state_regs_2_mix_columns_1_n211), .B(aes_state_regs_2_S00xDP[4]), 
        .ZN(aes_state_regs_2_mix_columns_1_n193) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U100 ( .A(
        aes_state_regs_2_mix_columns_1_n191), .B(
        aes_state_regs_2_mix_columns_1_n192), .ZN(
        aes_state_regs_2_MixColumnsS1xD[6]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U99 ( .A(aes_state_regs_2_S20xDP_5_), 
        .B(aes_state_regs_2_mix_columns_1_n229), .ZN(
        aes_state_regs_2_mix_columns_1_n192) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U98 ( .A(aes_state_regs_2_S00xDP[6]), 
        .B(aes_state_regs_2_S10xDP_5_), .Z(aes_state_regs_2_mix_columns_1_n191) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U97 ( .A(
        aes_state_regs_2_mix_columns_1_n190), .B(
        aes_state_regs_2_mix_columns_1_n215), .ZN(
        aes_state_regs_2_MixColumnsS0xD[2]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U96 ( .A(aes_state_regs_2_S30xDP_2_), 
        .B(aes_state_regs_2_mix_columns_1_n236), .ZN(
        aes_state_regs_2_mix_columns_1_n190) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U95 ( .A(
        aes_state_regs_2_mix_columns_1_n189), .B(
        aes_state_regs_2_mix_columns_1_n188), .ZN(
        aes_state_regs_2_MixColumnsS1xD[7]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U94 ( .A(aes_state_regs_2_S10xDP_6_), 
        .B(aes_state_regs_2_mix_columns_1_n231), .ZN(
        aes_state_regs_2_mix_columns_1_n189) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U93 ( .A1(aes_state_regs_2_S20xDP_6_), .A2(aes_state_regs_2_S20xDP_7_), .B1(aes_state_regs_2_mix_columns_1_n212), 
        .B2(aes_state_regs_2_mix_columns_1_n242), .ZN(
        aes_state_regs_2_mix_columns_1_n188) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U92 ( .A(
        aes_state_regs_2_mix_columns_1_n187), .B(
        aes_state_regs_2_mix_columns_1_n207), .ZN(
        aes_state_regs_2_MixColumnsS0xD[3]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U91 ( .A(aes_state_regs_2_S30xDP_3_), 
        .B(aes_state_regs_2_mix_columns_1_n237), .ZN(
        aes_state_regs_2_mix_columns_1_n187) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U90 ( .A(
        aes_state_regs_2_mix_columns_1_n186), .B(
        aes_state_regs_2_mix_columns_1_n233), .ZN(
        aes_state_regs_2_MixColumnsS3xD[0]) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U89 ( .A1(aes_state_regs_2_S20xDP_0_), .A2(aes_state_regs_2_mix_columns_1_n232), .B1(
        aes_state_regs_2_mix_columns_1_n231), .B2(
        aes_state_regs_2_mix_columns_1_n230), .ZN(
        aes_state_regs_2_mix_columns_1_n186) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U88 ( .A(
        aes_state_regs_2_mix_columns_1_n185), .B(
        aes_state_regs_2_mix_columns_1_n229), .ZN(
        aes_state_regs_2_MixColumnsS0xD[6]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U87 ( .A(aes_state_regs_2_S10xDP_6_), 
        .B(aes_state_regs_2_mix_columns_1_n241), .ZN(
        aes_state_regs_2_mix_columns_1_n185) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U86 ( .A1(aes_state_regs_2_S20xDP_3_), .A2(aes_state_regs_2_S20xDP_7_), .B1(aes_state_regs_2_mix_columns_1_n212), 
        .B2(aes_state_regs_2_mix_columns_1_n184), .ZN(
        aes_state_regs_2_mix_columns_1_n220) );
  INV_X1 aes_state_regs_2_mix_columns_1_U85 ( .A(aes_state_regs_2_S20xDP_3_), 
        .ZN(aes_state_regs_2_mix_columns_1_n184) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U84 ( .A(
        aes_state_regs_2_mix_columns_1_n183), .B(
        aes_state_regs_2_mix_columns_1_n233), .ZN(
        aes_state_regs_2_MixColumnsS2xD[0]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U83 ( .A(aes_state_regs_2_S20xDP_7_), 
        .B(aes_state_regs_2_mix_columns_1_n214), .ZN(
        aes_state_regs_2_mix_columns_1_n183) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U82 ( .A(
        aes_state_regs_2_mix_columns_1_n182), .B(
        aes_state_regs_2_mix_columns_1_n211), .ZN(
        aes_state_regs_2_MixColumnsS0xD[4]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U81 ( .A(aes_state_regs_2_S10xDP_4_), 
        .B(aes_state_regs_2_mix_columns_1_n239), .ZN(
        aes_state_regs_2_mix_columns_1_n182) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U80 ( .A(
        aes_state_regs_2_mix_columns_1_n181), .B(
        aes_state_regs_2_mix_columns_1_n238), .ZN(
        aes_state_regs_2_MixColumnsS3xD[3]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U79 ( .A(
        aes_state_regs_2_mix_columns_1_n237), .B(aes_state_regs_2_S00xDP[3]), 
        .ZN(aes_state_regs_2_mix_columns_1_n181) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U78 ( .A(
        aes_state_regs_2_mix_columns_1_n180), .B(
        aes_state_regs_2_mix_columns_1_n225), .ZN(
        aes_state_regs_2_MixColumnsS0xD[5]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U77 ( .A(aes_state_regs_2_S10xDP_5_), 
        .B(aes_state_regs_2_mix_columns_1_n222), .ZN(
        aes_state_regs_2_mix_columns_1_n180) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U76 ( .A(
        aes_state_regs_2_mix_columns_1_n179), .B(
        aes_state_regs_2_mix_columns_1_n235), .ZN(
        aes_state_regs_2_MixColumnsS3xD[1]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U75 ( .A(
        aes_state_regs_2_mix_columns_1_n234), .B(aes_state_regs_2_S20xDP_1_), 
        .ZN(aes_state_regs_2_mix_columns_1_n179) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U74 ( .A(
        aes_state_regs_2_mix_columns_1_n222), .B(
        aes_state_regs_2_mix_columns_1_n178), .ZN(
        aes_state_regs_2_mix_columns_1_n240) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U73 ( .A1(aes_state_regs_2_S30xDP_3_), .A2(aes_state_regs_2_mix_columns_1_n221), .B1(aes_state_regs_2_S30xDP_7_), 
        .B2(aes_state_regs_2_mix_columns_1_n177), .ZN(
        aes_state_regs_2_mix_columns_1_n178) );
  INV_X1 aes_state_regs_2_mix_columns_1_U72 ( .A(aes_state_regs_2_S30xDP_3_), 
        .ZN(aes_state_regs_2_mix_columns_1_n177) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U71 ( .A(
        aes_state_regs_2_mix_columns_1_n176), .B(
        aes_state_regs_2_mix_columns_1_n223), .ZN(
        aes_state_regs_2_mix_columns_1_n211) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U70 ( .A(aes_state_regs_2_S10xDP_7_), 
        .B(aes_state_regs_2_S10xDP_3_), .ZN(
        aes_state_regs_2_mix_columns_1_n176) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U69 ( .A(
        aes_state_regs_2_mix_columns_1_n174), .B(
        aes_state_regs_2_mix_columns_1_n175), .ZN(
        aes_state_regs_2_MixColumnsS3xD[2]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U68 ( .A(aes_state_regs_2_S30xDP_1_), 
        .B(aes_state_regs_2_S00xDP[2]), .ZN(
        aes_state_regs_2_mix_columns_1_n175) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U67 ( .A(aes_state_regs_2_S00xDP[1]), 
        .B(aes_state_regs_2_mix_columns_1_n236), .Z(
        aes_state_regs_2_mix_columns_1_n174) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U66 ( .A(
        aes_state_regs_2_mix_columns_1_n173), .B(aes_state_regs_2_S30xDP_7_), 
        .ZN(aes_state_regs_2_MixColumnsS0xD[7]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U65 ( .A(
        aes_state_regs_2_mix_columns_1_n244), .B(
        aes_state_regs_2_mix_columns_1_n243), .ZN(
        aes_state_regs_2_mix_columns_1_n173) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U64 ( .A(
        aes_state_regs_2_mix_columns_1_n172), .B(
        aes_state_regs_2_mix_columns_1_n240), .ZN(
        aes_state_regs_2_MixColumnsS3xD[4]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U63 ( .A(
        aes_state_regs_2_mix_columns_1_n239), .B(aes_state_regs_2_S20xDP_4_), 
        .ZN(aes_state_regs_2_mix_columns_1_n172) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U62 ( .A(
        aes_state_regs_2_mix_columns_1_n170), .B(
        aes_state_regs_2_mix_columns_1_n171), .ZN(
        aes_state_regs_2_MixColumnsS3xD[5]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U61 ( .A(
        aes_state_regs_2_mix_columns_1_n241), .B(aes_state_regs_2_S20xDP_5_), 
        .ZN(aes_state_regs_2_mix_columns_1_n171) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U60 ( .A(aes_state_regs_2_S00xDP[4]), 
        .B(aes_state_regs_2_S30xDP_4_), .Z(aes_state_regs_2_mix_columns_1_n170) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U59 ( .A(
        aes_state_regs_2_mix_columns_1_n168), .B(
        aes_state_regs_2_mix_columns_1_n169), .ZN(
        aes_state_regs_2_mix_columns_1_n237) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U58 ( .A(aes_state_regs_2_S20xDP_3_), 
        .B(aes_state_regs_2_S10xDP_3_), .ZN(
        aes_state_regs_2_mix_columns_1_n169) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U57 ( .A(aes_state_regs_2_S00xDP[2]), 
        .B(aes_state_regs_2_S00xDP[7]), .Z(aes_state_regs_2_mix_columns_1_n168) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U56 ( .A(
        aes_state_regs_2_mix_columns_1_n167), .B(
        aes_state_regs_2_mix_columns_1_n166), .ZN(
        aes_state_regs_2_MixColumnsS3xD[7]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U55 ( .A(
        aes_state_regs_2_mix_columns_1_n244), .B(aes_state_regs_2_S30xDP_6_), 
        .ZN(aes_state_regs_2_mix_columns_1_n167) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U54 ( .A1(aes_state_regs_2_S00xDP[6]), .A2(aes_state_regs_2_S00xDP[7]), .B1(aes_state_regs_2_mix_columns_1_n245), 
        .B2(aes_state_regs_2_mix_columns_1_n165), .ZN(
        aes_state_regs_2_mix_columns_1_n166) );
  INV_X1 aes_state_regs_2_mix_columns_1_U53 ( .A(aes_state_regs_2_S00xDP[6]), 
        .ZN(aes_state_regs_2_mix_columns_1_n165) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U52 ( .A(
        aes_state_regs_2_mix_columns_1_n164), .B(
        aes_state_regs_2_mix_columns_1_n235), .ZN(
        aes_state_regs_2_MixColumnsS2xD[1]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U51 ( .A(aes_state_regs_2_S30xDP_1_), 
        .B(aes_state_regs_2_mix_columns_1_n213), .ZN(
        aes_state_regs_2_mix_columns_1_n164) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U50 ( .A(
        aes_state_regs_2_mix_columns_1_n216), .B(
        aes_state_regs_2_mix_columns_1_n163), .ZN(
        aes_state_regs_2_MixColumnsS2xD[2]) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U49 ( .A(
        aes_state_regs_2_mix_columns_1_n217), .B(aes_state_regs_2_S10xDP_2_), 
        .Z(aes_state_regs_2_mix_columns_1_n163) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U48 ( .A(
        aes_state_regs_2_mix_columns_1_n162), .B(
        aes_state_regs_2_mix_columns_1_n238), .ZN(
        aes_state_regs_2_MixColumnsS2xD[3]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U47 ( .A(aes_state_regs_2_S10xDP_3_), 
        .B(aes_state_regs_2_mix_columns_1_n218), .ZN(
        aes_state_regs_2_mix_columns_1_n162) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U46 ( .A(
        aes_state_regs_2_mix_columns_1_n161), .B(
        aes_state_regs_2_mix_columns_1_n206), .ZN(
        aes_state_regs_2_MixColumnsS0xD[1]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U45 ( .A(aes_state_regs_2_S10xDP_1_), 
        .B(aes_state_regs_2_mix_columns_1_n234), .ZN(
        aes_state_regs_2_mix_columns_1_n161) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U44 ( .A(
        aes_state_regs_2_mix_columns_1_n160), .B(
        aes_state_regs_2_mix_columns_1_n240), .ZN(
        aes_state_regs_2_MixColumnsS2xD[4]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U43 ( .A(aes_state_regs_2_S30xDP_4_), 
        .B(aes_state_regs_2_mix_columns_1_n220), .ZN(
        aes_state_regs_2_mix_columns_1_n160) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U42 ( .A(
        aes_state_regs_2_mix_columns_1_n159), .B(
        aes_state_regs_2_mix_columns_1_n205), .ZN(
        aes_state_regs_2_MixColumnsS0xD[0]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U41 ( .A(aes_state_regs_2_S00xDP[7]), 
        .B(aes_state_regs_2_mix_columns_1_n204), .ZN(
        aes_state_regs_2_mix_columns_1_n159) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U40 ( .A(
        aes_state_regs_2_mix_columns_1_n223), .B(aes_state_regs_2_S30xDP_5_), 
        .ZN(aes_state_regs_2_mix_columns_1_n224) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U39 ( .A(
        aes_state_regs_2_mix_columns_1_n224), .B(
        aes_state_regs_2_mix_columns_1_n241), .ZN(
        aes_state_regs_2_MixColumnsS2xD[5]) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U38 ( .A(
        aes_state_regs_2_mix_columns_1_n225), .B(aes_state_regs_2_S30xDP_6_), 
        .ZN(aes_state_regs_2_mix_columns_1_n226) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U37 ( .A(
        aes_state_regs_2_mix_columns_1_n226), .B(
        aes_state_regs_2_mix_columns_1_n243), .ZN(
        aes_state_regs_2_MixColumnsS2xD[6]) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U36 ( .A1(aes_state_regs_2_S10xDP_7_), .A2(aes_state_regs_2_mix_columns_1_n232), .B1(
        aes_state_regs_2_mix_columns_1_n231), .B2(
        aes_state_regs_2_mix_columns_1_n227), .ZN(
        aes_state_regs_2_mix_columns_1_n228) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U35 ( .A(
        aes_state_regs_2_mix_columns_1_n229), .B(
        aes_state_regs_2_mix_columns_1_n228), .ZN(
        aes_state_regs_2_MixColumnsS2xD[7]) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U34 ( .A(aes_state_regs_2_S10xDP_0_), 
        .B(aes_state_regs_2_S00xDP[0]), .Z(aes_state_regs_2_mix_columns_1_n233) );
  INV_X1 aes_state_regs_2_mix_columns_1_U33 ( .A(
        aes_state_regs_2_mix_columns_1_n231), .ZN(
        aes_state_regs_2_mix_columns_1_n232) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U32 ( .A1(aes_state_regs_2_S00xDP[7]), .A2(aes_state_regs_2_S30xDP_7_), .B1(aes_state_regs_2_mix_columns_1_n221), 
        .B2(aes_state_regs_2_mix_columns_1_n245), .ZN(
        aes_state_regs_2_mix_columns_1_n231) );
  INV_X1 aes_state_regs_2_mix_columns_1_U31 ( .A(aes_state_regs_2_S20xDP_0_), 
        .ZN(aes_state_regs_2_mix_columns_1_n230) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U30 ( .A(aes_state_regs_2_S30xDP_0_), 
        .B(aes_state_regs_2_mix_columns_1_n221), .ZN(
        aes_state_regs_2_mix_columns_1_n214) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U29 ( .A1(aes_state_regs_2_S10xDP_7_), .A2(aes_state_regs_2_S20xDP_7_), .B1(aes_state_regs_2_mix_columns_1_n212), 
        .B2(aes_state_regs_2_mix_columns_1_n227), .ZN(
        aes_state_regs_2_mix_columns_1_n244) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U28 ( .A(aes_state_regs_2_S30xDP_0_), 
        .B(aes_state_regs_2_S20xDP_0_), .Z(aes_state_regs_2_mix_columns_1_n205) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U27 ( .A(
        aes_state_regs_2_mix_columns_1_n215), .B(
        aes_state_regs_2_mix_columns_1_n214), .Z(
        aes_state_regs_2_mix_columns_1_n235) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U26 ( .A(aes_state_regs_2_S00xDP[7]), 
        .B(aes_state_regs_2_S00xDP[0]), .Z(aes_state_regs_2_mix_columns_1_n234) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U25 ( .A(aes_state_regs_2_S10xDP_2_), 
        .B(aes_state_regs_2_S20xDP_2_), .Z(aes_state_regs_2_mix_columns_1_n236) );
  INV_X1 aes_state_regs_2_mix_columns_1_U24 ( .A(aes_state_regs_2_S30xDP_2_), 
        .ZN(aes_state_regs_2_mix_columns_1_n219) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U23 ( .A1(aes_state_regs_2_S30xDP_2_), .A2(aes_state_regs_2_S30xDP_7_), .B1(aes_state_regs_2_mix_columns_1_n221), 
        .B2(aes_state_regs_2_mix_columns_1_n219), .ZN(
        aes_state_regs_2_mix_columns_1_n238) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U22 ( .A(aes_state_regs_2_S00xDP[7]), 
        .B(aes_state_regs_2_S00xDP[3]), .Z(aes_state_regs_2_mix_columns_1_n239) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U21 ( .A(aes_state_regs_2_S10xDP_5_), 
        .B(aes_state_regs_2_S00xDP[5]), .Z(aes_state_regs_2_mix_columns_1_n241) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U20 ( .A(aes_state_regs_2_S10xDP_6_), 
        .B(aes_state_regs_2_S00xDP[6]), .Z(aes_state_regs_2_mix_columns_1_n243) );
  INV_X1 aes_state_regs_2_mix_columns_1_U19 ( .A(aes_state_regs_2_S20xDP_6_), 
        .ZN(aes_state_regs_2_mix_columns_1_n242) );
  INV_X1 aes_state_regs_2_mix_columns_1_U18 ( .A(aes_state_regs_2_S00xDP[7]), 
        .ZN(aes_state_regs_2_mix_columns_1_n245) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U17 ( .A1(aes_state_regs_2_S20xDP_0_), .A2(aes_state_regs_2_S20xDP_7_), .B1(aes_state_regs_2_mix_columns_1_n212), 
        .B2(aes_state_regs_2_mix_columns_1_n230), .ZN(
        aes_state_regs_2_mix_columns_1_n213) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U16 ( .A(aes_state_regs_2_S30xDP_2_), 
        .B(aes_state_regs_2_S00xDP[2]), .Z(aes_state_regs_2_mix_columns_1_n216) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U15 ( .A(aes_state_regs_2_S30xDP_1_), 
        .B(aes_state_regs_2_S20xDP_1_), .ZN(
        aes_state_regs_2_mix_columns_1_n217) );
  INV_X1 aes_state_regs_2_mix_columns_1_U14 ( .A(aes_state_regs_2_S00xDP[3]), 
        .ZN(aes_state_regs_2_mix_columns_1_n208) );
  AOI22_X1 aes_state_regs_2_mix_columns_1_U13 ( .A1(aes_state_regs_2_S00xDP[3]), .A2(aes_state_regs_2_S20xDP_7_), .B1(aes_state_regs_2_mix_columns_1_n212), 
        .B2(aes_state_regs_2_mix_columns_1_n208), .ZN(
        aes_state_regs_2_mix_columns_1_n209) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U12 ( .A(aes_state_regs_2_S20xDP_2_), 
        .B(aes_state_regs_2_S30xDP_3_), .ZN(
        aes_state_regs_2_mix_columns_1_n210) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U11 ( .A(aes_state_regs_2_S30xDP_4_), 
        .B(aes_state_regs_2_S20xDP_4_), .Z(aes_state_regs_2_mix_columns_1_n223) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U10 ( .A(aes_state_regs_2_S30xDP_5_), 
        .B(aes_state_regs_2_S20xDP_5_), .Z(aes_state_regs_2_mix_columns_1_n225) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U9 ( .A(aes_state_regs_2_S30xDP_6_), 
        .B(aes_state_regs_2_S20xDP_6_), .Z(aes_state_regs_2_mix_columns_1_n229) );
  INV_X1 aes_state_regs_2_mix_columns_1_U8 ( .A(aes_state_regs_2_S10xDP_7_), 
        .ZN(aes_state_regs_2_mix_columns_1_n227) );
  XNOR2_X1 aes_state_regs_2_mix_columns_1_U7 ( .A(
        aes_state_regs_2_mix_columns_1_n204), .B(
        aes_state_regs_2_mix_columns_1_n217), .ZN(
        aes_state_regs_2_mix_columns_1_n206) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U6 ( .A(aes_state_regs_2_S10xDP_7_), 
        .B(aes_state_regs_2_S10xDP_2_), .Z(aes_state_regs_2_mix_columns_1_n207) );
  INV_X1 aes_state_regs_2_mix_columns_1_U5 ( .A(aes_state_regs_2_S20xDP_7_), 
        .ZN(aes_state_regs_2_mix_columns_1_n212) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U4 ( .A(aes_state_regs_2_S10xDP_4_), 
        .B(aes_state_regs_2_S00xDP[4]), .Z(aes_state_regs_2_mix_columns_1_n222) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U3 ( .A(aes_state_regs_2_S10xDP_1_), 
        .B(aes_state_regs_2_S00xDP[1]), .Z(aes_state_regs_2_mix_columns_1_n215) );
  INV_X1 aes_state_regs_2_mix_columns_1_U2 ( .A(aes_state_regs_2_S30xDP_7_), 
        .ZN(aes_state_regs_2_mix_columns_1_n221) );
  XOR2_X1 aes_state_regs_2_mix_columns_1_U1 ( .A(aes_state_regs_2_S10xDP_7_), 
        .B(aes_state_regs_2_S10xDP_0_), .Z(aes_state_regs_2_mix_columns_1_n204) );
  BUF_X1 aes_key_regs_1_U3 ( .A(n170), .Z(aes_key_regs_1_n4) );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_0_ ( .D(aes_key_regs_1_K00xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_0_ ( .D(aes_key_regs_1_K10xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_0_ ( .D(aes_key_regs_1_K20xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_0_ ( .D(aes_key_regs_1_K01xDP_0_), .SI(
        KeyOutxD[8]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_0_ ( .D(aes_key_regs_1_K01xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_0_ ( .D(aes_key_regs_1_K11xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_0_ ( .D(aes_key_regs_1_K21xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_0_ ( .D(aes_key_regs_1_K02xDP_0_), .SI(
        aes_key_regs_1_K01xDP_0_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_0_ ( .D(aes_key_regs_1_K02xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_0_ ( .D(aes_key_regs_1_K12xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_0_ ( .D(aes_key_regs_1_K22xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_0_ ( .D(K03xD[8]), .SI(
        aes_key_regs_1_K02xDP_0_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_1_ ( .D(aes_key_regs_1_K00xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_1_ ( .D(aes_key_regs_1_K10xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_1_ ( .D(aes_key_regs_1_K20xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_1_ ( .D(aes_key_regs_1_K01xDP_1_), .SI(
        KeyOutxD[9]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_1_ ( .D(aes_key_regs_1_K01xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_1_ ( .D(aes_key_regs_1_K11xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_1_ ( .D(aes_key_regs_1_K21xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_1_ ( .D(aes_key_regs_1_K02xDP_1_), .SI(
        aes_key_regs_1_K01xDP_1_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_1_ ( .D(aes_key_regs_1_K02xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_1_ ( .D(aes_key_regs_1_K12xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_1_ ( .D(aes_key_regs_1_K22xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_1_ ( .D(K03xD[9]), .SI(
        aes_key_regs_1_K02xDP_1_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_2_ ( .D(aes_key_regs_1_K00xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_2_ ( .D(aes_key_regs_1_K10xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_2_ ( .D(aes_key_regs_1_K20xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_2_ ( .D(aes_key_regs_1_K01xDP_2_), .SI(
        KeyOutxD[10]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_2_ ( .D(aes_key_regs_1_K01xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_2_ ( .D(aes_key_regs_1_K11xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_2_ ( .D(aes_key_regs_1_K21xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_2_ ( .D(aes_key_regs_1_K02xDP_2_), .SI(
        aes_key_regs_1_K01xDP_2_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_2_ ( .D(aes_key_regs_1_K02xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_2_ ( .D(aes_key_regs_1_K12xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_2_ ( .D(aes_key_regs_1_K22xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_2_ ( .D(K03xD[10]), .SI(
        aes_key_regs_1_K02xDP_2_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_3_ ( .D(aes_key_regs_1_K00xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_3_ ( .D(aes_key_regs_1_K10xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_3_ ( .D(aes_key_regs_1_K20xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_3_ ( .D(aes_key_regs_1_K01xDP_3_), .SI(
        KeyOutxD[11]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_3_ ( .D(aes_key_regs_1_K01xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_3_ ( .D(aes_key_regs_1_K11xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_3_ ( .D(aes_key_regs_1_K21xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_3_ ( .D(aes_key_regs_1_K02xDP_3_), .SI(
        aes_key_regs_1_K01xDP_3_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_3_ ( .D(aes_key_regs_1_K02xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_3_ ( .D(aes_key_regs_1_K12xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_3_ ( .D(aes_key_regs_1_K22xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_3_ ( .D(K03xD[11]), .SI(
        aes_key_regs_1_K02xDP_3_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_4_ ( .D(aes_key_regs_1_K00xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_4_ ( .D(aes_key_regs_1_K10xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_4_ ( .D(aes_key_regs_1_K20xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_4_ ( .D(aes_key_regs_1_K01xDP_4_), .SI(
        KeyOutxD[12]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_4_ ( .D(aes_key_regs_1_K01xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_4_ ( .D(aes_key_regs_1_K11xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_4_ ( .D(aes_key_regs_1_K21xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_4_ ( .D(aes_key_regs_1_K02xDP_4_), .SI(
        aes_key_regs_1_K01xDP_4_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_4_ ( .D(aes_key_regs_1_K02xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_4_ ( .D(aes_key_regs_1_K12xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_4_ ( .D(aes_key_regs_1_K22xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_4_ ( .D(K03xD[12]), .SI(
        aes_key_regs_1_K02xDP_4_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_5_ ( .D(aes_key_regs_1_K00xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_5_ ( .D(aes_key_regs_1_K10xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_5_ ( .D(aes_key_regs_1_K20xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_5_ ( .D(aes_key_regs_1_K01xDP_5_), .SI(
        KeyOutxD[13]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_5_ ( .D(aes_key_regs_1_K01xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_5_ ( .D(aes_key_regs_1_K11xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_5_ ( .D(aes_key_regs_1_K21xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_5_ ( .D(aes_key_regs_1_K02xDP_5_), .SI(
        aes_key_regs_1_K01xDP_5_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_5_ ( .D(aes_key_regs_1_K02xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_5_ ( .D(aes_key_regs_1_K12xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_5_ ( .D(aes_key_regs_1_K22xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_5_ ( .D(K03xD[13]), .SI(
        aes_key_regs_1_K02xDP_5_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_6_ ( .D(aes_key_regs_1_K00xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_6_ ( .D(aes_key_regs_1_K10xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_6_ ( .D(aes_key_regs_1_K20xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_6_ ( .D(aes_key_regs_1_K01xDP_6_), .SI(
        KeyOutxD[14]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_6_ ( .D(aes_key_regs_1_K01xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_6_ ( .D(aes_key_regs_1_K11xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_6_ ( .D(aes_key_regs_1_K21xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_6_ ( .D(aes_key_regs_1_K02xDP_6_), .SI(
        aes_key_regs_1_K01xDP_6_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_6_ ( .D(aes_key_regs_1_K02xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_6_ ( .D(aes_key_regs_1_K12xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_6_ ( .D(aes_key_regs_1_K22xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_6_ ( .D(K03xD[14]), .SI(
        aes_key_regs_1_K02xDP_6_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_7_ ( .D(aes_key_regs_1_K00xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_7_ ( .D(aes_key_regs_1_K10xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_7_ ( .D(aes_key_regs_1_K20xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_7_ ( .D(aes_key_regs_1_K01xDP_7_), .SI(
        KeyOutxD[15]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_7_ ( .D(aes_key_regs_1_K01xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_7_ ( .D(aes_key_regs_1_K11xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_7_ ( .D(aes_key_regs_1_K21xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_7_ ( .D(aes_key_regs_1_K02xDP_7_), .SI(
        aes_key_regs_1_K01xDP_7_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_7_ ( .D(aes_key_regs_1_K02xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_7_ ( .D(aes_key_regs_1_K12xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_7_ ( .D(aes_key_regs_1_K22xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_7_ ( .D(K03xD[15]), .SI(
        aes_key_regs_1_K02xDP_7_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_0_ ( .D(KeyInxD[8]), .SI(K03xD[8]), .SE(
        n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K23xDN[0]), 
        .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_0_ ( .D(KeyToSboxOutxD[8]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_0_ ( .D(aes_key_regs_1_K13xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_0_ ( .D(aes_key_regs_1_K23xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_1_ ( .D(KeyInxD[9]), .SI(K03xD[9]), .SE(
        aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_1_ ( .D(KeyToSboxOutxD[9]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_1_ ( .D(aes_key_regs_1_K13xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_1_ ( .D(aes_key_regs_1_K23xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_2_ ( .D(KeyInxD[10]), .SI(K03xD[10]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K23xDN[2]), 
        .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_2_ ( .D(KeyToSboxOutxD[10]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_2_ ( .D(aes_key_regs_1_K13xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_2_ ( .D(aes_key_regs_1_K23xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_3_ ( .D(KeyInxD[11]), .SI(K03xD[11]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K23xDN[3]), 
        .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_3_ ( .D(KeyToSboxOutxD[11]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_3_ ( .D(aes_key_regs_1_K13xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_3_ ( .D(aes_key_regs_1_K23xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_4_ ( .D(KeyInxD[12]), .SI(K03xD[12]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K23xDN[4]), 
        .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_4_ ( .D(KeyToSboxOutxD[12]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_4_ ( .D(aes_key_regs_1_K13xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_4_ ( .D(aes_key_regs_1_K23xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_5_ ( .D(KeyInxD[13]), .SI(K03xD[13]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K23xDN[5]), 
        .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_5_ ( .D(KeyToSboxOutxD[13]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_5_ ( .D(aes_key_regs_1_K13xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_5_ ( .D(aes_key_regs_1_K23xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_6_ ( .D(KeyInxD[14]), .SI(K03xD[14]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K23xDN[6]), 
        .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_6_ ( .D(KeyToSboxOutxD[14]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_6_ ( .D(aes_key_regs_1_K13xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_6_ ( .D(aes_key_regs_1_K23xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_7_ ( .D(KeyInxD[15]), .SI(K03xD[15]), 
        .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K23xDN[7]), 
        .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_7_ ( .D(KeyToSboxOutxD[15]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_7_ ( .D(aes_key_regs_1_K13xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_7_ ( .D(aes_key_regs_1_K23xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[7]), .QN() );
  OAI222_X1 aes_state_regs_1_U55 ( .A1(aes_state_regs_1_n190), .A2(
        aes_state_regs_1_n109), .B1(aes_state_regs_1_n197), .B2(
        aes_state_regs_1_n44), .C1(aes_state_regs_1_n183), .C2(
        aes_state_regs_1_n127), .ZN(aes_state_regs_1_S10xDN[7]) );
  INV_X1 aes_state_regs_1_U54 ( .A(aes_state_regs_1_MixColumnsS2xD[7]), .ZN(
        aes_state_regs_1_n190) );
  OAI222_X1 aes_state_regs_1_U53 ( .A1(aes_state_regs_1_n189), .A2(
        aes_state_regs_1_n109), .B1(aes_state_regs_1_n197), .B2(
        aes_state_regs_1_n45), .C1(aes_state_regs_1_n183), .C2(
        aes_state_regs_1_n126), .ZN(aes_state_regs_1_S10xDN[6]) );
  INV_X1 aes_state_regs_1_U52 ( .A(aes_state_regs_1_MixColumnsS2xD[6]), .ZN(
        aes_state_regs_1_n189) );
  OAI222_X1 aes_state_regs_1_U51 ( .A1(aes_state_regs_1_n188), .A2(
        aes_state_regs_1_n109), .B1(aes_state_regs_1_n197), .B2(
        aes_state_regs_1_n46), .C1(aes_state_regs_1_n183), .C2(
        aes_state_regs_1_n125), .ZN(aes_state_regs_1_S10xDN[5]) );
  INV_X1 aes_state_regs_1_U50 ( .A(aes_state_regs_1_MixColumnsS2xD[5]), .ZN(
        aes_state_regs_1_n188) );
  OAI222_X1 aes_state_regs_1_U49 ( .A1(aes_state_regs_1_n187), .A2(
        aes_state_regs_1_n109), .B1(aes_state_regs_1_n197), .B2(
        aes_state_regs_1_n47), .C1(aes_state_regs_1_n183), .C2(
        aes_state_regs_1_n124), .ZN(aes_state_regs_1_S10xDN[4]) );
  INV_X1 aes_state_regs_1_U48 ( .A(aes_state_regs_1_MixColumnsS2xD[4]), .ZN(
        aes_state_regs_1_n187) );
  OAI222_X1 aes_state_regs_1_U47 ( .A1(aes_state_regs_1_n186), .A2(
        aes_state_regs_1_n109), .B1(aes_state_regs_1_n197), .B2(
        aes_state_regs_1_n48), .C1(aes_state_regs_1_n183), .C2(
        aes_state_regs_1_n123), .ZN(aes_state_regs_1_S10xDN[3]) );
  INV_X1 aes_state_regs_1_U46 ( .A(aes_state_regs_1_MixColumnsS2xD[3]), .ZN(
        aes_state_regs_1_n186) );
  OAI222_X1 aes_state_regs_1_U45 ( .A1(aes_state_regs_1_n185), .A2(
        aes_state_regs_1_n109), .B1(aes_state_regs_1_n197), .B2(
        aes_state_regs_1_n49), .C1(aes_state_regs_1_n183), .C2(
        aes_state_regs_1_n122), .ZN(aes_state_regs_1_S10xDN[2]) );
  INV_X1 aes_state_regs_1_U44 ( .A(aes_state_regs_1_MixColumnsS2xD[2]), .ZN(
        aes_state_regs_1_n185) );
  OAI222_X1 aes_state_regs_1_U43 ( .A1(aes_state_regs_1_n184), .A2(
        aes_state_regs_1_n109), .B1(aes_state_regs_1_n197), .B2(
        aes_state_regs_1_n50), .C1(aes_state_regs_1_n183), .C2(
        aes_state_regs_1_n121), .ZN(aes_state_regs_1_S10xDN[1]) );
  INV_X1 aes_state_regs_1_U42 ( .A(aes_state_regs_1_MixColumnsS2xD[1]), .ZN(
        aes_state_regs_1_n184) );
  NAND2_X1 aes_state_regs_1_U41 ( .A1(doMixColumnsxS), .A2(
        aes_state_regs_1_n183), .ZN(aes_state_regs_1_n109) );
  INV_X1 aes_state_regs_1_U40 ( .A(n453), .ZN(aes_state_regs_1_n183) );
  INV_X8 aes_state_regs_1_U39 ( .A(aes_state_regs_1_n183), .ZN(
        aes_state_regs_1_n182) );
  OAI21_X1 aes_state_regs_1_U38 ( .B1(aes_state_regs_1_n43), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n180), .ZN(
        aes_state_regs_1_S20xDN[0]) );
  AOI22_X1 aes_state_regs_1_U37 ( .A1(aes_state_regs_1_MixColumnsS3xD[0]), 
        .A2(aes_state_regs_1_n202), .B1(aes_state_regs_1_n136), .B2(
        aes_state_regs_1_n182), .ZN(aes_state_regs_1_n180) );
  OAI21_X1 aes_state_regs_1_U36 ( .B1(aes_state_regs_1_n51), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n179), .ZN(
        aes_state_regs_1_S10xDN[0]) );
  AOI22_X1 aes_state_regs_1_U35 ( .A1(aes_state_regs_1_n182), .A2(
        aes_state_regs_1_n138), .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_MixColumnsS2xD[0]), .ZN(aes_state_regs_1_n179) );
  OAI21_X1 aes_state_regs_1_U34 ( .B1(aes_state_regs_1_n42), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n178), .ZN(
        aes_state_regs_1_S20xDN[1]) );
  AOI22_X1 aes_state_regs_1_U33 ( .A1(aes_state_regs_1_MixColumnsS3xD[1]), 
        .A2(aes_state_regs_1_n202), .B1(aes_state_regs_1_n141), .B2(
        aes_state_regs_1_n182), .ZN(aes_state_regs_1_n178) );
  OAI21_X1 aes_state_regs_1_U32 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n33), .A(aes_state_regs_1_n177), .ZN(StateOutxD[12])
         );
  NAND2_X1 aes_state_regs_1_U31 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[4]), .ZN(aes_state_regs_1_n177) );
  OAI21_X1 aes_state_regs_1_U30 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n29), .A(aes_state_regs_1_n176), .ZN(StateOutxD[15])
         );
  NAND2_X1 aes_state_regs_1_U29 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[7]), .ZN(aes_state_regs_1_n176) );
  OAI21_X1 aes_state_regs_1_U28 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n35), .A(aes_state_regs_1_n175), .ZN(StateOutxD[14])
         );
  NAND2_X1 aes_state_regs_1_U27 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[6]), .ZN(aes_state_regs_1_n175) );
  OAI21_X1 aes_state_regs_1_U26 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n31), .A(aes_state_regs_1_n174), .ZN(StateOutxD[10])
         );
  NAND2_X1 aes_state_regs_1_U25 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[2]), .ZN(aes_state_regs_1_n174) );
  AOI22_X1 aes_state_regs_1_U24 ( .A1(aes_state_regs_1_n182), .A2(
        aes_state_regs_1_n146), .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_MixColumnsS3xD[2]), .ZN(aes_state_regs_1_n191) );
  OAI21_X1 aes_state_regs_1_U23 ( .B1(aes_state_regs_1_n41), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n191), .ZN(
        aes_state_regs_1_S20xDN[2]) );
  AOI22_X1 aes_state_regs_1_U22 ( .A1(aes_state_regs_1_n182), .A2(
        aes_state_regs_1_n151), .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_MixColumnsS3xD[3]), .ZN(aes_state_regs_1_n192) );
  OAI21_X1 aes_state_regs_1_U21 ( .B1(aes_state_regs_1_n40), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n192), .ZN(
        aes_state_regs_1_S20xDN[3]) );
  AOI22_X1 aes_state_regs_1_U20 ( .A1(aes_state_regs_1_n182), .A2(
        aes_state_regs_1_n156), .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_MixColumnsS3xD[4]), .ZN(aes_state_regs_1_n193) );
  OAI21_X1 aes_state_regs_1_U19 ( .B1(aes_state_regs_1_n39), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n193), .ZN(
        aes_state_regs_1_S20xDN[4]) );
  AOI22_X1 aes_state_regs_1_U18 ( .A1(aes_state_regs_1_n182), .A2(
        aes_state_regs_1_n161), .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_MixColumnsS3xD[5]), .ZN(aes_state_regs_1_n194) );
  OAI21_X1 aes_state_regs_1_U17 ( .B1(aes_state_regs_1_n38), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n194), .ZN(
        aes_state_regs_1_S20xDN[5]) );
  AOI22_X1 aes_state_regs_1_U16 ( .A1(aes_state_regs_1_n182), .A2(
        aes_state_regs_1_n166), .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_MixColumnsS3xD[6]), .ZN(aes_state_regs_1_n195) );
  OAI21_X1 aes_state_regs_1_U15 ( .B1(aes_state_regs_1_n37), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n195), .ZN(
        aes_state_regs_1_S20xDN[6]) );
  AOI22_X1 aes_state_regs_1_U14 ( .A1(aes_state_regs_1_n182), .A2(
        aes_state_regs_1_n171), .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_MixColumnsS3xD[7]), .ZN(aes_state_regs_1_n196) );
  OAI21_X1 aes_state_regs_1_U13 ( .B1(aes_state_regs_1_n36), .B2(
        aes_state_regs_1_n197), .A(aes_state_regs_1_n196), .ZN(
        aes_state_regs_1_S20xDN[7]) );
  NAND2_X1 aes_state_regs_1_U12 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[5]), .ZN(aes_state_regs_1_n198) );
  OAI21_X1 aes_state_regs_1_U11 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n34), .A(aes_state_regs_1_n198), .ZN(StateOutxD[13])
         );
  NAND2_X1 aes_state_regs_1_U10 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[3]), .ZN(aes_state_regs_1_n199) );
  OAI21_X1 aes_state_regs_1_U9 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n32), .A(aes_state_regs_1_n199), .ZN(StateOutxD[11])
         );
  NAND2_X1 aes_state_regs_1_U8 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[1]), .ZN(aes_state_regs_1_n200) );
  OAI21_X1 aes_state_regs_1_U7 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n30), .A(aes_state_regs_1_n200), .ZN(StateOutxD[9])
         );
  NAND2_X1 aes_state_regs_1_U6 ( .A1(aes_state_regs_1_n202), .A2(
        aes_state_regs_1_MixColumnsS0xD[0]), .ZN(aes_state_regs_1_n201) );
  OAI21_X1 aes_state_regs_1_U5 ( .B1(aes_state_regs_1_n202), .B2(
        aes_state_regs_1_n28), .A(aes_state_regs_1_n201), .ZN(StateOutxD[8])
         );
  OR2_X1 aes_state_regs_1_U4 ( .A1(aes_state_regs_1_n182), .A2(doMixColumnsxS), 
        .ZN(aes_state_regs_1_n197) );
  INV_X2 aes_state_regs_1_U3 ( .A(aes_state_regs_1_n109), .ZN(
        aes_state_regs_1_n202) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_7_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[7]), .SI(aes_state_regs_1_S10xDP_7_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[7]), .QN(aes_state_regs_1_n29) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_6_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[6]), .SI(aes_state_regs_1_S10xDP_6_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[6]), .QN(aes_state_regs_1_n35) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_5_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[5]), .SI(aes_state_regs_1_S10xDP_5_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[5]), .QN(aes_state_regs_1_n34) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_4_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[4]), .SI(aes_state_regs_1_S10xDP_4_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[4]), .QN(aes_state_regs_1_n33) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_3_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[3]), .SI(aes_state_regs_1_S10xDP_3_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[3]), .QN(aes_state_regs_1_n32) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_2_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[2]), .SI(aes_state_regs_1_S10xDP_2_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[2]), .QN(aes_state_regs_1_n31) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_1_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[1]), .SI(aes_state_regs_1_S10xDP_1_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[1]), .QN(aes_state_regs_1_n30) );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_7_ ( .D(aes_state_regs_1_S10xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_7_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_6_ ( .D(aes_state_regs_1_S10xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_6_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_5_ ( .D(aes_state_regs_1_S10xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_5_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_4_ ( .D(aes_state_regs_1_S10xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_4_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_3_ ( .D(aes_state_regs_1_S10xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_3_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_2_ ( .D(aes_state_regs_1_S10xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_2_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_1_ ( .D(aes_state_regs_1_S10xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_7_ ( .D(aes_state_regs_1_S01xDO_7_), 
        .SI(StateInxD[15]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S30xDP_7_), .QN(aes_state_regs_1_n36) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_7_ ( .D(aes_state_regs_1_n173), .SI(
        aes_state_regs_1_n170), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[7]), .QN(aes_state_regs_1_n127) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_7_ ( .D(aes_state_regs_1_S02xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_7_ ( .D(aes_state_regs_1_n172), .SI(
        aes_state_regs_1_S23xDP_7_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_7_ ( .D(aes_state_regs_1_n170), .SI(
        aes_state_regs_1_n173), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_7_ ( .D(aes_state_regs_1_S02xDP_7_), 
        .SI(aes_state_regs_1_S01xDO_7_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n173), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_7_ ( .D(aes_state_regs_1_S01xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_7_ ( .D(aes_state_regs_1_S21xDP[7]), 
        .SI(aes_state_regs_1_n172), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_7_ ( .D(aes_state_regs_1_n171), .SI(
        aes_state_regs_1_S30xDP_7_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n172), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_7_ ( .D(aes_state_regs_1_n169), .SI(
        aes_state_regs_1_S02xDP_7_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n171), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_7_ ( .D(StateInxD[15]), .SI(
        aes_state_regs_1_n169), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n170), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_7_ ( .D(aes_state_regs_1_S03xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n169), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_7_ ( .D(aes_state_regs_1_S23xDP_7_), 
        .SI(aes_state_regs_1_S20xDP_7_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[7]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_7_ ( .D(aes_state_regs_1_S20xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_7_), .QN(
        aes_state_regs_1_n44) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_6_ ( .D(aes_state_regs_1_S01xDO_6_), 
        .SI(StateInxD[14]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S30xDP_6_), .QN(aes_state_regs_1_n37) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_6_ ( .D(aes_state_regs_1_n168), .SI(
        aes_state_regs_1_n165), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[6]), .QN(aes_state_regs_1_n126) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_6_ ( .D(aes_state_regs_1_S02xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_6_ ( .D(aes_state_regs_1_n167), .SI(
        aes_state_regs_1_S23xDP_6_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_6_ ( .D(aes_state_regs_1_n165), .SI(
        aes_state_regs_1_n168), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_6_ ( .D(aes_state_regs_1_S02xDP_6_), 
        .SI(aes_state_regs_1_S01xDO_6_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n168), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_6_ ( .D(aes_state_regs_1_S01xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_6_ ( .D(aes_state_regs_1_S21xDP[6]), 
        .SI(aes_state_regs_1_n167), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_6_ ( .D(aes_state_regs_1_n166), .SI(
        aes_state_regs_1_S30xDP_6_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n167), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_6_ ( .D(aes_state_regs_1_n164), .SI(
        aes_state_regs_1_S02xDP_6_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n166), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_6_ ( .D(StateInxD[14]), .SI(
        aes_state_regs_1_n164), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n165), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_6_ ( .D(aes_state_regs_1_S03xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n164), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_6_ ( .D(aes_state_regs_1_S23xDP_6_), 
        .SI(aes_state_regs_1_S20xDP_6_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[6]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_6_ ( .D(aes_state_regs_1_S20xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_6_), .QN(
        aes_state_regs_1_n45) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_5_ ( .D(aes_state_regs_1_S01xDO_5_), 
        .SI(StateInxD[13]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S30xDP_5_), .QN(aes_state_regs_1_n38) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_5_ ( .D(aes_state_regs_1_n163), .SI(
        aes_state_regs_1_n160), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[5]), .QN(aes_state_regs_1_n125) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_5_ ( .D(aes_state_regs_1_S02xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_5_ ( .D(aes_state_regs_1_n162), .SI(
        aes_state_regs_1_S23xDP_5_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_5_ ( .D(aes_state_regs_1_n160), .SI(
        aes_state_regs_1_n163), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_5_ ( .D(aes_state_regs_1_S02xDP_5_), 
        .SI(aes_state_regs_1_S01xDO_5_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n163), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_5_ ( .D(aes_state_regs_1_S01xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_5_ ( .D(aes_state_regs_1_S21xDP[5]), 
        .SI(aes_state_regs_1_n162), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_5_ ( .D(aes_state_regs_1_n161), .SI(
        aes_state_regs_1_S30xDP_5_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n162), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_5_ ( .D(aes_state_regs_1_n159), .SI(
        aes_state_regs_1_S02xDP_5_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n161), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_5_ ( .D(StateInxD[13]), .SI(
        aes_state_regs_1_n159), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n160), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_5_ ( .D(aes_state_regs_1_S03xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n159), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_5_ ( .D(aes_state_regs_1_S23xDP_5_), 
        .SI(aes_state_regs_1_S20xDP_5_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[5]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_5_ ( .D(aes_state_regs_1_S20xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_5_), .QN(
        aes_state_regs_1_n46) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_4_ ( .D(aes_state_regs_1_S01xDO_4_), 
        .SI(StateInxD[12]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S30xDP_4_), .QN(aes_state_regs_1_n39) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_4_ ( .D(aes_state_regs_1_n158), .SI(
        aes_state_regs_1_n155), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[4]), .QN(aes_state_regs_1_n124) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_4_ ( .D(aes_state_regs_1_S02xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_4_ ( .D(aes_state_regs_1_n157), .SI(
        aes_state_regs_1_S23xDP_4_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_4_ ( .D(aes_state_regs_1_n155), .SI(
        aes_state_regs_1_n158), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_4_ ( .D(aes_state_regs_1_S02xDP_4_), 
        .SI(aes_state_regs_1_S01xDO_4_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n158), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_4_ ( .D(aes_state_regs_1_S01xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_4_ ( .D(aes_state_regs_1_S21xDP[4]), 
        .SI(aes_state_regs_1_n157), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_4_ ( .D(aes_state_regs_1_n156), .SI(
        aes_state_regs_1_S30xDP_4_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n157), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_4_ ( .D(aes_state_regs_1_n154), .SI(
        aes_state_regs_1_S02xDP_4_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n156), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_4_ ( .D(StateInxD[12]), .SI(
        aes_state_regs_1_n154), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n155), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_4_ ( .D(aes_state_regs_1_S03xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n154), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_4_ ( .D(aes_state_regs_1_S23xDP_4_), 
        .SI(aes_state_regs_1_S20xDP_4_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[4]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_4_ ( .D(aes_state_regs_1_S20xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_4_), .QN(
        aes_state_regs_1_n47) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_3_ ( .D(aes_state_regs_1_S01xDO_3_), 
        .SI(StateInxD[11]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S30xDP_3_), .QN(aes_state_regs_1_n40) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_3_ ( .D(aes_state_regs_1_n153), .SI(
        aes_state_regs_1_n150), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[3]), .QN(aes_state_regs_1_n123) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_3_ ( .D(aes_state_regs_1_S02xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_3_ ( .D(aes_state_regs_1_n152), .SI(
        aes_state_regs_1_S23xDP_3_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_3_ ( .D(aes_state_regs_1_n150), .SI(
        aes_state_regs_1_n153), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_3_ ( .D(aes_state_regs_1_S02xDP_3_), 
        .SI(aes_state_regs_1_S01xDO_3_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n153), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_3_ ( .D(aes_state_regs_1_S01xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_3_ ( .D(aes_state_regs_1_S21xDP[3]), 
        .SI(aes_state_regs_1_n152), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_3_ ( .D(aes_state_regs_1_n151), .SI(
        aes_state_regs_1_S30xDP_3_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n152), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_3_ ( .D(aes_state_regs_1_n149), .SI(
        aes_state_regs_1_S02xDP_3_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n151), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_3_ ( .D(StateInxD[11]), .SI(
        aes_state_regs_1_n149), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n150), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_3_ ( .D(aes_state_regs_1_S03xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n149), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_3_ ( .D(aes_state_regs_1_S23xDP_3_), 
        .SI(aes_state_regs_1_S20xDP_3_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[3]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_3_ ( .D(aes_state_regs_1_S20xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_3_), .QN(
        aes_state_regs_1_n48) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_2_ ( .D(aes_state_regs_1_S01xDO_2_), 
        .SI(StateInxD[10]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S30xDP_2_), .QN(aes_state_regs_1_n41) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_2_ ( .D(aes_state_regs_1_n148), .SI(
        aes_state_regs_1_n145), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[2]), .QN(aes_state_regs_1_n122) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_2_ ( .D(aes_state_regs_1_S02xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_2_ ( .D(aes_state_regs_1_n147), .SI(
        aes_state_regs_1_S23xDP_2_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_2_ ( .D(aes_state_regs_1_n145), .SI(
        aes_state_regs_1_n148), .SE(n453), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S23xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_2_ ( .D(aes_state_regs_1_S02xDP_2_), 
        .SI(aes_state_regs_1_S01xDO_2_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n148), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_2_ ( .D(aes_state_regs_1_S01xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_2_ ( .D(aes_state_regs_1_S21xDP[2]), 
        .SI(aes_state_regs_1_n147), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_2_ ( .D(aes_state_regs_1_n146), .SI(
        aes_state_regs_1_S30xDP_2_), .SE(n453), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_n147), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_2_ ( .D(aes_state_regs_1_n144), .SI(
        aes_state_regs_1_S02xDP_2_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n146), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_2_ ( .D(StateInxD[10]), .SI(
        aes_state_regs_1_n144), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n145), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_2_ ( .D(aes_state_regs_1_S03xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n144), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_2_ ( .D(aes_state_regs_1_S23xDP_2_), 
        .SI(aes_state_regs_1_S20xDP_2_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[2]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_2_ ( .D(aes_state_regs_1_S20xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_2_), .QN(
        aes_state_regs_1_n49) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_1_ ( .D(aes_state_regs_1_S01xDO_1_), 
        .SI(StateInxD[9]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_1_), .QN(aes_state_regs_1_n42) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_1_ ( .D(aes_state_regs_1_n143), .SI(
        aes_state_regs_1_n140), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[1]), .QN(aes_state_regs_1_n121) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_1_ ( .D(aes_state_regs_1_S02xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_1_ ( .D(aes_state_regs_1_n142), .SI(
        aes_state_regs_1_S23xDP_1_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_1_ ( .D(aes_state_regs_1_n140), .SI(
        aes_state_regs_1_n143), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_1_ ( .D(aes_state_regs_1_S02xDP_1_), 
        .SI(aes_state_regs_1_S01xDO_1_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n143), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_1_ ( .D(aes_state_regs_1_S01xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_1_ ( .D(aes_state_regs_1_S21xDP[1]), 
        .SI(aes_state_regs_1_n142), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_1_ ( .D(aes_state_regs_1_n141), .SI(
        aes_state_regs_1_S30xDP_1_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n142), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_1_ ( .D(aes_state_regs_1_n139), .SI(
        aes_state_regs_1_S02xDP_1_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n141), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_1_ ( .D(StateInxD[9]), .SI(
        aes_state_regs_1_n139), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n140), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_1_ ( .D(aes_state_regs_1_S03xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n139), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_1_ ( .D(aes_state_regs_1_S23xDP_1_), 
        .SI(aes_state_regs_1_S20xDP_1_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[1]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_1_ ( .D(aes_state_regs_1_S20xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_1_), .QN(
        aes_state_regs_1_n50) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_0_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[0]), .SI(aes_state_regs_1_S10xDP_0_), 
        .SE(aes_state_regs_1_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[0]), .QN(aes_state_regs_1_n28) );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_0_ ( .D(aes_state_regs_1_S10xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_0_ ( .D(aes_state_regs_1_n137), .SI(
        aes_state_regs_1_S31xDP_0_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S23xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_0_ ( .D(aes_state_regs_1_S02xDP_0_), 
        .SI(aes_state_regs_1_S01xDO_0_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S31xDP_0_), .QN() );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_0_ ( .D(aes_state_regs_1_S02xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_0_ ( .D(aes_state_regs_1_S22xDP_0_), 
        .SI(aes_state_regs_1_S23xDP_0_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_0_ ( .D(aes_state_regs_1_n136), .SI(
        aes_state_regs_1_S30xDP_0_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S22xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_0_ ( .D(aes_state_regs_1_S01xDO_0_), 
        .SI(StateInxD[8]), .SE(aes_state_regs_1_n182), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_0_), .QN(aes_state_regs_1_n43) );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_0_ ( .D(aes_state_regs_1_S01xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_0_ ( .D(aes_state_regs_1_n138), .SI(
        aes_state_regs_1_S22xDP_0_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_0_ ( .D(aes_state_regs_1_S31xDP_0_), 
        .SI(aes_state_regs_1_n137), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n138), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_0_ ( .D(StateInxD[8]), .SI(
        aes_state_regs_1_S03xDP_0_), .SE(aes_state_regs_1_n182), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n137), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_0_ ( .D(aes_state_regs_1_S03xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_0_ ( .D(aes_state_regs_1_S23xDP_0_), 
        .SI(aes_state_regs_1_S20xDP_0_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[0]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_0_ ( .D(aes_state_regs_1_S20xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_0_), .QN(
        aes_state_regs_1_n51) );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_0_ ( .D(aes_state_regs_1_S03xDP_0_), 
        .SI(aes_state_regs_1_S02xDP_0_), .SE(aes_state_regs_1_n182), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n136), .QN() );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U119 ( .A(
        aes_state_regs_1_mix_columns_1_n245), .B(
        aes_state_regs_1_mix_columns_1_n244), .ZN(
        aes_state_regs_1_MixColumnsS3xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U118 ( .A(
        aes_state_regs_1_mix_columns_1_n240), .B(
        aes_state_regs_1_mix_columns_1_n239), .ZN(
        aes_state_regs_1_MixColumnsS3xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U117 ( .A(
        aes_state_regs_1_mix_columns_1_n235), .B(
        aes_state_regs_1_mix_columns_1_n234), .ZN(
        aes_state_regs_1_MixColumnsS3xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U116 ( .A(
        aes_state_regs_1_mix_columns_1_n226), .B(
        aes_state_regs_1_mix_columns_1_n225), .ZN(
        aes_state_regs_1_MixColumnsS3xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U115 ( .A(
        aes_state_regs_1_mix_columns_1_n187), .B(
        aes_state_regs_1_mix_columns_1_n241), .ZN(
        aes_state_regs_1_MixColumnsS1xD[0]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U114 ( .A(
        aes_state_regs_1_mix_columns_1_n193), .B(aes_state_regs_1_S00xDP[0]), 
        .ZN(aes_state_regs_1_mix_columns_1_n187) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U113 ( .A(
        aes_state_regs_1_mix_columns_1_n185), .B(
        aes_state_regs_1_mix_columns_1_n186), .ZN(
        aes_state_regs_1_MixColumnsS1xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U112 ( .A(aes_state_regs_1_S20xDP_1_), .B(aes_state_regs_1_S20xDP_2_), .ZN(aes_state_regs_1_mix_columns_1_n186) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U111 ( .A(
        aes_state_regs_1_mix_columns_1_n202), .B(aes_state_regs_1_S10xDP_1_), 
        .Z(aes_state_regs_1_mix_columns_1_n185) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U110 ( .A(
        aes_state_regs_1_mix_columns_1_n209), .B(
        aes_state_regs_1_mix_columns_1_n184), .ZN(
        aes_state_regs_1_mix_columns_1_n231) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U109 ( .A1(
        aes_state_regs_1_S30xDP_3_), .A2(aes_state_regs_1_mix_columns_1_n208), 
        .B1(aes_state_regs_1_S30xDP_7_), .B2(
        aes_state_regs_1_mix_columns_1_n183), .ZN(
        aes_state_regs_1_mix_columns_1_n184) );
  INV_X1 aes_state_regs_1_mix_columns_1_U108 ( .A(aes_state_regs_1_S30xDP_3_), 
        .ZN(aes_state_regs_1_mix_columns_1_n183) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U107 ( .A(
        aes_state_regs_1_mix_columns_1_n182), .B(
        aes_state_regs_1_mix_columns_1_n221), .ZN(
        aes_state_regs_1_MixColumnsS3xD[0]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U106 ( .A1(
        aes_state_regs_1_S20xDP_0_), .A2(aes_state_regs_1_mix_columns_1_n220), 
        .B1(aes_state_regs_1_mix_columns_1_n219), .B2(
        aes_state_regs_1_mix_columns_1_n218), .ZN(
        aes_state_regs_1_mix_columns_1_n182) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U105 ( .A(
        aes_state_regs_1_mix_columns_1_n181), .B(
        aes_state_regs_1_mix_columns_1_n205), .ZN(
        aes_state_regs_1_MixColumnsS1xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U104 ( .A(aes_state_regs_1_S20xDP_3_), .B(aes_state_regs_1_mix_columns_1_n195), .ZN(
        aes_state_regs_1_mix_columns_1_n181) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U103 ( .A(
        aes_state_regs_1_mix_columns_1_n179), .B(
        aes_state_regs_1_mix_columns_1_n180), .ZN(
        aes_state_regs_1_MixColumnsS1xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U102 ( .A(aes_state_regs_1_S20xDP_4_), .B(aes_state_regs_1_mix_columns_1_n213), .ZN(
        aes_state_regs_1_mix_columns_1_n180) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U101 ( .A(aes_state_regs_1_S00xDP[5]), 
        .B(aes_state_regs_1_S10xDP_4_), .Z(aes_state_regs_1_mix_columns_1_n179) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U100 ( .A(
        aes_state_regs_1_mix_columns_1_n178), .B(
        aes_state_regs_1_mix_columns_1_n221), .ZN(
        aes_state_regs_1_MixColumnsS2xD[0]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U99 ( .A(aes_state_regs_1_S20xDP_7_), 
        .B(aes_state_regs_1_mix_columns_1_n199), .ZN(
        aes_state_regs_1_mix_columns_1_n178) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U98 ( .A(
        aes_state_regs_1_mix_columns_1_n176), .B(
        aes_state_regs_1_mix_columns_1_n177), .ZN(
        aes_state_regs_1_MixColumnsS1xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U97 ( .A(aes_state_regs_1_S20xDP_5_), 
        .B(aes_state_regs_1_mix_columns_1_n217), .ZN(
        aes_state_regs_1_mix_columns_1_n177) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U96 ( .A(aes_state_regs_1_S00xDP[6]), 
        .B(aes_state_regs_1_S10xDP_5_), .Z(aes_state_regs_1_mix_columns_1_n176) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U95 ( .A(
        aes_state_regs_1_mix_columns_1_n175), .B(
        aes_state_regs_1_mix_columns_1_n211), .ZN(
        aes_state_regs_1_mix_columns_1_n196) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U94 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_3_), .ZN(
        aes_state_regs_1_mix_columns_1_n175) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U93 ( .A(
        aes_state_regs_1_mix_columns_1_n174), .B(
        aes_state_regs_1_mix_columns_1_n223), .ZN(
        aes_state_regs_1_MixColumnsS3xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U92 ( .A(
        aes_state_regs_1_mix_columns_1_n222), .B(aes_state_regs_1_S20xDP_1_), 
        .ZN(aes_state_regs_1_mix_columns_1_n174) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U91 ( .A(
        aes_state_regs_1_mix_columns_1_n173), .B(
        aes_state_regs_1_mix_columns_1_n198), .ZN(
        aes_state_regs_1_MixColumnsS1xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U90 ( .A(
        aes_state_regs_1_mix_columns_1_n194), .B(aes_state_regs_1_S00xDP[1]), 
        .ZN(aes_state_regs_1_mix_columns_1_n173) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U89 ( .A1(aes_state_regs_1_S30xDP_2_), .A2(aes_state_regs_1_S30xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n208), 
        .B2(aes_state_regs_1_mix_columns_1_n172), .ZN(
        aes_state_regs_1_mix_columns_1_n228) );
  INV_X1 aes_state_regs_1_mix_columns_1_U88 ( .A(aes_state_regs_1_S30xDP_2_), 
        .ZN(aes_state_regs_1_mix_columns_1_n172) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U87 ( .A(
        aes_state_regs_1_mix_columns_1_n171), .B(
        aes_state_regs_1_mix_columns_1_n207), .ZN(
        aes_state_regs_1_MixColumnsS1xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U86 ( .A(
        aes_state_regs_1_mix_columns_1_n196), .B(aes_state_regs_1_S00xDP[4]), 
        .ZN(aes_state_regs_1_mix_columns_1_n171) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U85 ( .A(
        aes_state_regs_1_mix_columns_1_n169), .B(
        aes_state_regs_1_mix_columns_1_n170), .ZN(
        aes_state_regs_1_MixColumnsS1xD[7]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U84 ( .A1(aes_state_regs_1_S20xDP_6_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n197), 
        .B2(aes_state_regs_1_mix_columns_1_n236), .ZN(
        aes_state_regs_1_mix_columns_1_n170) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U83 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_mix_columns_1_n219), .ZN(
        aes_state_regs_1_mix_columns_1_n169) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U82 ( .A(
        aes_state_regs_1_mix_columns_1_n167), .B(
        aes_state_regs_1_mix_columns_1_n168), .ZN(
        aes_state_regs_1_mix_columns_1_n227) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U81 ( .A(aes_state_regs_1_S20xDP_3_), 
        .B(aes_state_regs_1_S10xDP_3_), .ZN(
        aes_state_regs_1_mix_columns_1_n168) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U80 ( .A(aes_state_regs_1_S00xDP[2]), 
        .B(aes_state_regs_1_S00xDP[7]), .Z(aes_state_regs_1_mix_columns_1_n167) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U79 ( .A(
        aes_state_regs_1_mix_columns_1_n166), .B(
        aes_state_regs_1_mix_columns_1_n196), .ZN(
        aes_state_regs_1_MixColumnsS0xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U78 ( .A(aes_state_regs_1_S10xDP_4_), 
        .B(aes_state_regs_1_mix_columns_1_n230), .ZN(
        aes_state_regs_1_mix_columns_1_n166) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U77 ( .A(
        aes_state_regs_1_mix_columns_1_n163), .B(
        aes_state_regs_1_mix_columns_1_n165), .ZN(
        aes_state_regs_1_mix_columns_1_n205) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U76 ( .A1(aes_state_regs_1_S00xDP[3]), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n197), 
        .B2(aes_state_regs_1_mix_columns_1_n164), .ZN(
        aes_state_regs_1_mix_columns_1_n165) );
  INV_X1 aes_state_regs_1_mix_columns_1_U75 ( .A(aes_state_regs_1_S00xDP[3]), 
        .ZN(aes_state_regs_1_mix_columns_1_n164) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U74 ( .A(aes_state_regs_1_S20xDP_2_), 
        .B(aes_state_regs_1_S30xDP_3_), .ZN(
        aes_state_regs_1_mix_columns_1_n163) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U73 ( .A(
        aes_state_regs_1_mix_columns_1_n162), .B(aes_state_regs_1_S30xDP_7_), 
        .ZN(aes_state_regs_1_MixColumnsS0xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U72 ( .A(
        aes_state_regs_1_mix_columns_1_n241), .B(
        aes_state_regs_1_mix_columns_1_n238), .ZN(
        aes_state_regs_1_mix_columns_1_n162) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U71 ( .A(
        aes_state_regs_1_mix_columns_1_n161), .B(
        aes_state_regs_1_mix_columns_1_n217), .ZN(
        aes_state_regs_1_MixColumnsS0xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U70 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_mix_columns_1_n233), .ZN(
        aes_state_regs_1_mix_columns_1_n161) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U69 ( .A1(aes_state_regs_1_S20xDP_3_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n197), 
        .B2(aes_state_regs_1_mix_columns_1_n160), .ZN(
        aes_state_regs_1_mix_columns_1_n207) );
  INV_X1 aes_state_regs_1_mix_columns_1_U68 ( .A(aes_state_regs_1_S20xDP_3_), 
        .ZN(aes_state_regs_1_mix_columns_1_n160) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U67 ( .A(
        aes_state_regs_1_mix_columns_1_n159), .B(
        aes_state_regs_1_mix_columns_1_n200), .ZN(
        aes_state_regs_1_MixColumnsS0xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U66 ( .A(aes_state_regs_1_S30xDP_2_), 
        .B(aes_state_regs_1_mix_columns_1_n224), .ZN(
        aes_state_regs_1_mix_columns_1_n159) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U65 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_mix_columns_1_n224), .ZN(
        aes_state_regs_1_mix_columns_1_n225) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U64 ( .A(aes_state_regs_1_S00xDP[2]), 
        .B(aes_state_regs_1_S00xDP[1]), .Z(aes_state_regs_1_mix_columns_1_n226) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U63 ( .A(
        aes_state_regs_1_mix_columns_1_n227), .B(aes_state_regs_1_S00xDP[3]), 
        .ZN(aes_state_regs_1_mix_columns_1_n229) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U62 ( .A(
        aes_state_regs_1_mix_columns_1_n229), .B(
        aes_state_regs_1_mix_columns_1_n228), .ZN(
        aes_state_regs_1_MixColumnsS3xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U61 ( .A(
        aes_state_regs_1_mix_columns_1_n230), .B(aes_state_regs_1_S20xDP_4_), 
        .ZN(aes_state_regs_1_mix_columns_1_n232) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U60 ( .A(
        aes_state_regs_1_mix_columns_1_n232), .B(
        aes_state_regs_1_mix_columns_1_n231), .ZN(
        aes_state_regs_1_MixColumnsS3xD[4]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U59 ( .A(
        aes_state_regs_1_mix_columns_1_n233), .B(aes_state_regs_1_S20xDP_5_), 
        .Z(aes_state_regs_1_mix_columns_1_n235) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U58 ( .A(aes_state_regs_1_S30xDP_4_), 
        .B(aes_state_regs_1_S00xDP[4]), .ZN(
        aes_state_regs_1_mix_columns_1_n234) );
  INV_X1 aes_state_regs_1_mix_columns_1_U57 ( .A(
        aes_state_regs_1_mix_columns_1_n238), .ZN(
        aes_state_regs_1_mix_columns_1_n237) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U56 ( .A1(aes_state_regs_1_S20xDP_6_), .A2(aes_state_regs_1_mix_columns_1_n238), .B1(
        aes_state_regs_1_mix_columns_1_n237), .B2(
        aes_state_regs_1_mix_columns_1_n236), .ZN(
        aes_state_regs_1_mix_columns_1_n239) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U55 ( .A(aes_state_regs_1_S30xDP_5_), 
        .B(aes_state_regs_1_S00xDP[5]), .ZN(
        aes_state_regs_1_mix_columns_1_n240) );
  INV_X1 aes_state_regs_1_mix_columns_1_U54 ( .A(aes_state_regs_1_S00xDP[6]), 
        .ZN(aes_state_regs_1_mix_columns_1_n243) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U53 ( .A(aes_state_regs_1_S30xDP_6_), 
        .B(aes_state_regs_1_mix_columns_1_n241), .ZN(
        aes_state_regs_1_mix_columns_1_n245) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U52 ( .A1(aes_state_regs_1_S00xDP[7]), .A2(aes_state_regs_1_S00xDP[6]), .B1(aes_state_regs_1_mix_columns_1_n243), 
        .B2(aes_state_regs_1_mix_columns_1_n242), .ZN(
        aes_state_regs_1_mix_columns_1_n244) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U51 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_mix_columns_1_n198), .ZN(
        aes_state_regs_1_mix_columns_1_n201) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U50 ( .A(
        aes_state_regs_1_mix_columns_1_n201), .B(
        aes_state_regs_1_mix_columns_1_n223), .ZN(
        aes_state_regs_1_MixColumnsS2xD[1]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U49 ( .A(aes_state_regs_1_S10xDP_2_), 
        .B(aes_state_regs_1_mix_columns_1_n202), .Z(
        aes_state_regs_1_mix_columns_1_n203) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U48 ( .A(
        aes_state_regs_1_mix_columns_1_n204), .B(
        aes_state_regs_1_mix_columns_1_n203), .ZN(
        aes_state_regs_1_MixColumnsS2xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U47 ( .A(aes_state_regs_1_S10xDP_3_), 
        .B(aes_state_regs_1_mix_columns_1_n205), .ZN(
        aes_state_regs_1_mix_columns_1_n206) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U46 ( .A(
        aes_state_regs_1_mix_columns_1_n206), .B(
        aes_state_regs_1_mix_columns_1_n228), .ZN(
        aes_state_regs_1_MixColumnsS2xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U45 ( .A(aes_state_regs_1_S30xDP_4_), 
        .B(aes_state_regs_1_mix_columns_1_n207), .ZN(
        aes_state_regs_1_mix_columns_1_n210) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U44 ( .A(
        aes_state_regs_1_mix_columns_1_n210), .B(
        aes_state_regs_1_mix_columns_1_n231), .ZN(
        aes_state_regs_1_MixColumnsS2xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U43 ( .A(
        aes_state_regs_1_mix_columns_1_n211), .B(aes_state_regs_1_S30xDP_5_), 
        .ZN(aes_state_regs_1_mix_columns_1_n212) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U42 ( .A(
        aes_state_regs_1_mix_columns_1_n212), .B(
        aes_state_regs_1_mix_columns_1_n233), .ZN(
        aes_state_regs_1_MixColumnsS2xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U41 ( .A(
        aes_state_regs_1_mix_columns_1_n213), .B(aes_state_regs_1_S30xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n214) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U40 ( .A(
        aes_state_regs_1_mix_columns_1_n214), .B(
        aes_state_regs_1_mix_columns_1_n238), .ZN(
        aes_state_regs_1_MixColumnsS2xD[6]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U39 ( .A1(aes_state_regs_1_S10xDP_7_), .A2(aes_state_regs_1_mix_columns_1_n220), .B1(
        aes_state_regs_1_mix_columns_1_n219), .B2(
        aes_state_regs_1_mix_columns_1_n215), .ZN(
        aes_state_regs_1_mix_columns_1_n216) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U38 ( .A(
        aes_state_regs_1_mix_columns_1_n217), .B(
        aes_state_regs_1_mix_columns_1_n216), .ZN(
        aes_state_regs_1_MixColumnsS2xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U37 ( .A(aes_state_regs_1_S10xDP_5_), 
        .B(aes_state_regs_1_mix_columns_1_n209), .ZN(
        aes_state_regs_1_mix_columns_1_n192) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U36 ( .A(
        aes_state_regs_1_mix_columns_1_n192), .B(
        aes_state_regs_1_mix_columns_1_n213), .ZN(
        aes_state_regs_1_MixColumnsS0xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U35 ( .A(aes_state_regs_1_S30xDP_3_), 
        .B(aes_state_regs_1_mix_columns_1_n227), .ZN(
        aes_state_regs_1_mix_columns_1_n191) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U34 ( .A(
        aes_state_regs_1_mix_columns_1_n191), .B(
        aes_state_regs_1_mix_columns_1_n195), .ZN(
        aes_state_regs_1_MixColumnsS0xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U33 ( .A(aes_state_regs_1_S10xDP_1_), 
        .B(aes_state_regs_1_mix_columns_1_n222), .ZN(
        aes_state_regs_1_mix_columns_1_n190) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U32 ( .A(
        aes_state_regs_1_mix_columns_1_n190), .B(
        aes_state_regs_1_mix_columns_1_n194), .ZN(
        aes_state_regs_1_MixColumnsS0xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U31 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_mix_columns_1_n189), .ZN(
        aes_state_regs_1_mix_columns_1_n188) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U30 ( .A(
        aes_state_regs_1_mix_columns_1_n188), .B(
        aes_state_regs_1_mix_columns_1_n193), .ZN(
        aes_state_regs_1_MixColumnsS0xD[0]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U29 ( .A(aes_state_regs_1_S10xDP_0_), 
        .B(aes_state_regs_1_S00xDP[0]), .Z(aes_state_regs_1_mix_columns_1_n221) );
  INV_X1 aes_state_regs_1_mix_columns_1_U28 ( .A(
        aes_state_regs_1_mix_columns_1_n219), .ZN(
        aes_state_regs_1_mix_columns_1_n220) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U27 ( .A1(aes_state_regs_1_S00xDP[7]), .A2(aes_state_regs_1_S30xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n208), 
        .B2(aes_state_regs_1_mix_columns_1_n242), .ZN(
        aes_state_regs_1_mix_columns_1_n219) );
  INV_X1 aes_state_regs_1_mix_columns_1_U26 ( .A(aes_state_regs_1_S20xDP_0_), 
        .ZN(aes_state_regs_1_mix_columns_1_n218) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U25 ( .A(aes_state_regs_1_S30xDP_0_), 
        .B(aes_state_regs_1_mix_columns_1_n208), .ZN(
        aes_state_regs_1_mix_columns_1_n199) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U24 ( .A1(aes_state_regs_1_S10xDP_7_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n197), 
        .B2(aes_state_regs_1_mix_columns_1_n215), .ZN(
        aes_state_regs_1_mix_columns_1_n241) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U23 ( .A(aes_state_regs_1_S30xDP_0_), 
        .B(aes_state_regs_1_S20xDP_0_), .Z(aes_state_regs_1_mix_columns_1_n193) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U22 ( .A(
        aes_state_regs_1_mix_columns_1_n200), .B(
        aes_state_regs_1_mix_columns_1_n199), .Z(
        aes_state_regs_1_mix_columns_1_n223) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U21 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_S00xDP[0]), .Z(aes_state_regs_1_mix_columns_1_n222) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U20 ( .A(aes_state_regs_1_S10xDP_2_), 
        .B(aes_state_regs_1_S20xDP_2_), .Z(aes_state_regs_1_mix_columns_1_n224) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U19 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_S00xDP[3]), .Z(aes_state_regs_1_mix_columns_1_n230) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U18 ( .A(aes_state_regs_1_S10xDP_5_), 
        .B(aes_state_regs_1_S00xDP[5]), .Z(aes_state_regs_1_mix_columns_1_n233) );
  INV_X1 aes_state_regs_1_mix_columns_1_U17 ( .A(aes_state_regs_1_S20xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n236) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U16 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_S00xDP[6]), .Z(aes_state_regs_1_mix_columns_1_n238) );
  INV_X1 aes_state_regs_1_mix_columns_1_U15 ( .A(aes_state_regs_1_S00xDP[7]), 
        .ZN(aes_state_regs_1_mix_columns_1_n242) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U14 ( .A1(aes_state_regs_1_S20xDP_0_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n197), 
        .B2(aes_state_regs_1_mix_columns_1_n218), .ZN(
        aes_state_regs_1_mix_columns_1_n198) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U13 ( .A(aes_state_regs_1_S30xDP_2_), 
        .B(aes_state_regs_1_S00xDP[2]), .Z(aes_state_regs_1_mix_columns_1_n202) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U12 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_S20xDP_1_), .ZN(
        aes_state_regs_1_mix_columns_1_n204) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U11 ( .A(aes_state_regs_1_S30xDP_4_), 
        .B(aes_state_regs_1_S20xDP_4_), .Z(aes_state_regs_1_mix_columns_1_n211) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U10 ( .A(aes_state_regs_1_S30xDP_5_), 
        .B(aes_state_regs_1_S20xDP_5_), .Z(aes_state_regs_1_mix_columns_1_n213) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U9 ( .A(aes_state_regs_1_S30xDP_6_), 
        .B(aes_state_regs_1_S20xDP_6_), .Z(aes_state_regs_1_mix_columns_1_n217) );
  INV_X1 aes_state_regs_1_mix_columns_1_U8 ( .A(aes_state_regs_1_S10xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n215) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U7 ( .A(
        aes_state_regs_1_mix_columns_1_n189), .B(
        aes_state_regs_1_mix_columns_1_n204), .ZN(
        aes_state_regs_1_mix_columns_1_n194) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U6 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_2_), .Z(aes_state_regs_1_mix_columns_1_n195) );
  INV_X1 aes_state_regs_1_mix_columns_1_U5 ( .A(aes_state_regs_1_S20xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n197) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U4 ( .A(aes_state_regs_1_S10xDP_4_), 
        .B(aes_state_regs_1_S00xDP[4]), .Z(aes_state_regs_1_mix_columns_1_n209) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U3 ( .A(aes_state_regs_1_S10xDP_1_), 
        .B(aes_state_regs_1_S00xDP[1]), .Z(aes_state_regs_1_mix_columns_1_n200) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U2 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_0_), .Z(aes_state_regs_1_mix_columns_1_n189) );
  INV_X1 aes_state_regs_1_mix_columns_1_U1 ( .A(aes_state_regs_1_S30xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n208) );
  BUF_X1 aes_key_regs_0_U3 ( .A(n170), .Z(aes_key_regs_0_n4) );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_0_ ( .D(aes_key_regs_0_K00xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_0_ ( .D(aes_key_regs_0_K10xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_0_ ( .D(aes_key_regs_0_K20xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_0_ ( .D(aes_key_regs_0_K01xDP_0_), .SI(
        KeyOutxD[0]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_0_ ( .D(aes_key_regs_0_K01xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_0_ ( .D(aes_key_regs_0_K11xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_0_ ( .D(aes_key_regs_0_K21xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_0_ ( .D(aes_key_regs_0_K02xDP_0_), .SI(
        aes_key_regs_0_K01xDP_0_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_0_ ( .D(aes_key_regs_0_K02xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_0_ ( .D(aes_key_regs_0_K12xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_0_ ( .D(aes_key_regs_0_K22xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_0_ ( .D(K03xD[0]), .SI(
        aes_key_regs_0_K02xDP_0_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_1_ ( .D(aes_key_regs_0_K00xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_1_ ( .D(aes_key_regs_0_K10xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_1_ ( .D(aes_key_regs_0_K20xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_1_ ( .D(aes_key_regs_0_K01xDP_1_), .SI(
        KeyOutxD[1]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_1_ ( .D(aes_key_regs_0_K01xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_1_ ( .D(aes_key_regs_0_K11xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_1_ ( .D(aes_key_regs_0_K21xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_1_ ( .D(aes_key_regs_0_K02xDP_1_), .SI(
        aes_key_regs_0_K01xDP_1_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_1_ ( .D(aes_key_regs_0_K02xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_1_ ( .D(aes_key_regs_0_K12xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_1_ ( .D(aes_key_regs_0_K22xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_1_ ( .D(K03xD[1]), .SI(
        aes_key_regs_0_K02xDP_1_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_2_ ( .D(aes_key_regs_0_K00xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_2_ ( .D(aes_key_regs_0_K10xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_2_ ( .D(aes_key_regs_0_K20xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_2_ ( .D(aes_key_regs_0_K01xDP_2_), .SI(
        KeyOutxD[2]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_2_ ( .D(aes_key_regs_0_K01xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_2_ ( .D(aes_key_regs_0_K11xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_2_ ( .D(aes_key_regs_0_K21xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_2_ ( .D(aes_key_regs_0_K02xDP_2_), .SI(
        aes_key_regs_0_K01xDP_2_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_2_ ( .D(aes_key_regs_0_K02xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_2_ ( .D(aes_key_regs_0_K12xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_2_ ( .D(aes_key_regs_0_K22xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_2_ ( .D(K03xD[2]), .SI(
        aes_key_regs_0_K02xDP_2_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_3_ ( .D(aes_key_regs_0_K00xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_3_ ( .D(aes_key_regs_0_K10xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_3_ ( .D(aes_key_regs_0_K20xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_3_ ( .D(aes_key_regs_0_K01xDP_3_), .SI(
        KeyOutxD[3]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_3_ ( .D(aes_key_regs_0_K01xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_3_ ( .D(aes_key_regs_0_K11xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_3_ ( .D(aes_key_regs_0_K21xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_3_ ( .D(aes_key_regs_0_K02xDP_3_), .SI(
        aes_key_regs_0_K01xDP_3_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_3_ ( .D(aes_key_regs_0_K02xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_3_ ( .D(aes_key_regs_0_K12xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_3_ ( .D(aes_key_regs_0_K22xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_3_ ( .D(K03xD[3]), .SI(
        aes_key_regs_0_K02xDP_3_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_4_ ( .D(aes_key_regs_0_K00xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_4_ ( .D(aes_key_regs_0_K10xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_4_ ( .D(aes_key_regs_0_K20xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_4_ ( .D(aes_key_regs_0_K01xDP_4_), .SI(
        KeyOutxD[4]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_4_ ( .D(aes_key_regs_0_K01xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_4_ ( .D(aes_key_regs_0_K11xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_4_ ( .D(aes_key_regs_0_K21xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_4_ ( .D(aes_key_regs_0_K02xDP_4_), .SI(
        aes_key_regs_0_K01xDP_4_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_4_ ( .D(aes_key_regs_0_K02xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_4_ ( .D(aes_key_regs_0_K12xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_4_ ( .D(aes_key_regs_0_K22xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_4_ ( .D(K03xD[4]), .SI(
        aes_key_regs_0_K02xDP_4_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_5_ ( .D(aes_key_regs_0_K00xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_5_ ( .D(aes_key_regs_0_K10xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_5_ ( .D(aes_key_regs_0_K20xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_5_ ( .D(aes_key_regs_0_K01xDP_5_), .SI(
        KeyOutxD[5]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_5_ ( .D(aes_key_regs_0_K01xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_5_ ( .D(aes_key_regs_0_K11xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_5_ ( .D(aes_key_regs_0_K21xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_5_ ( .D(aes_key_regs_0_K02xDP_5_), .SI(
        aes_key_regs_0_K01xDP_5_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_5_ ( .D(aes_key_regs_0_K02xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_5_ ( .D(aes_key_regs_0_K12xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_5_ ( .D(aes_key_regs_0_K22xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_5_ ( .D(K03xD[5]), .SI(
        aes_key_regs_0_K02xDP_5_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_6_ ( .D(aes_key_regs_0_K00xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_6_ ( .D(aes_key_regs_0_K10xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_6_ ( .D(aes_key_regs_0_K20xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_6_ ( .D(aes_key_regs_0_K01xDP_6_), .SI(
        KeyOutxD[6]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_6_ ( .D(aes_key_regs_0_K01xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_6_ ( .D(aes_key_regs_0_K11xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_6_ ( .D(aes_key_regs_0_K21xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_6_ ( .D(aes_key_regs_0_K02xDP_6_), .SI(
        aes_key_regs_0_K01xDP_6_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_6_ ( .D(aes_key_regs_0_K02xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_6_ ( .D(aes_key_regs_0_K12xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_6_ ( .D(aes_key_regs_0_K22xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_6_ ( .D(K03xD[6]), .SI(
        aes_key_regs_0_K02xDP_6_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_7_ ( .D(aes_key_regs_0_K00xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_7_ ( .D(aes_key_regs_0_K10xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_7_ ( .D(aes_key_regs_0_K20xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_7_ ( .D(aes_key_regs_0_K01xDP_7_), .SI(
        KeyOutxD[7]), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_7_ ( .D(aes_key_regs_0_K01xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_7_ ( .D(aes_key_regs_0_K11xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_7_ ( .D(aes_key_regs_0_K21xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_7_ ( .D(aes_key_regs_0_K02xDP_7_), .SI(
        aes_key_regs_0_K01xDP_7_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_7_ ( .D(aes_key_regs_0_K02xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_7_ ( .D(aes_key_regs_0_K12xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_7_ ( .D(aes_key_regs_0_K22xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_7_ ( .D(K03xD[7]), .SI(
        aes_key_regs_0_K02xDP_7_), .SE(n170), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_0_ ( .D(KeyInxD[0]), .SI(K03xD[0]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_0_ ( .D(KeyToSboxOutxD[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_0_ ( .D(aes_key_regs_0_K13xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_0_ ( .D(aes_key_regs_0_K23xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_1_ ( .D(KeyInxD[1]), .SI(K03xD[1]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_1_ ( .D(KeyToSboxOutxD[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_1_ ( .D(aes_key_regs_0_K13xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_1_ ( .D(aes_key_regs_0_K23xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_2_ ( .D(KeyInxD[2]), .SI(K03xD[2]), .SE(
        n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[2]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_2_ ( .D(KeyToSboxOutxD[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_2_ ( .D(aes_key_regs_0_K13xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_2_ ( .D(aes_key_regs_0_K23xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_3_ ( .D(KeyInxD[3]), .SI(K03xD[3]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_3_ ( .D(KeyToSboxOutxD[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_3_ ( .D(aes_key_regs_0_K13xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_3_ ( .D(aes_key_regs_0_K23xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_4_ ( .D(KeyInxD[4]), .SI(K03xD[4]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_4_ ( .D(KeyToSboxOutxD[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_4_ ( .D(aes_key_regs_0_K13xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_4_ ( .D(aes_key_regs_0_K23xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_5_ ( .D(KeyInxD[5]), .SI(K03xD[5]), .SE(
        n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[5]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_5_ ( .D(KeyToSboxOutxD[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_5_ ( .D(aes_key_regs_0_K13xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_5_ ( .D(aes_key_regs_0_K23xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_6_ ( .D(KeyInxD[6]), .SI(K03xD[6]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_6_ ( .D(KeyToSboxOutxD[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_6_ ( .D(aes_key_regs_0_K13xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_6_ ( .D(aes_key_regs_0_K23xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_7_ ( .D(KeyInxD[7]), .SI(K03xD[7]), .SE(
        n170), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K23xDN[7]), 
        .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_7_ ( .D(KeyToSboxOutxD[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_7_ ( .D(aes_key_regs_0_K13xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_7_ ( .D(aes_key_regs_0_K23xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[7]), .QN() );
  AOI22_X1 aes_state_regs_0_U56 ( .A1(aes_state_regs_0_n178), .A2(
        aes_state_regs_0_n171), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[7]), .ZN(aes_state_regs_0_n196) );
  AOI22_X1 aes_state_regs_0_U55 ( .A1(aes_state_regs_0_n178), .A2(
        aes_state_regs_0_n166), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[6]), .ZN(aes_state_regs_0_n195) );
  AOI22_X1 aes_state_regs_0_U54 ( .A1(aes_state_regs_0_n178), .A2(
        aes_state_regs_0_n161), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[5]), .ZN(aes_state_regs_0_n194) );
  AOI22_X1 aes_state_regs_0_U53 ( .A1(aes_state_regs_0_n179), .A2(
        aes_state_regs_0_n151), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[3]), .ZN(aes_state_regs_0_n192) );
  AOI22_X1 aes_state_regs_0_U52 ( .A1(aes_state_regs_0_n179), .A2(
        aes_state_regs_0_n146), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[2]), .ZN(aes_state_regs_0_n191) );
  AOI22_X1 aes_state_regs_0_U51 ( .A1(aes_state_regs_0_n179), .A2(
        aes_state_regs_0_n141), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[1]), .ZN(aes_state_regs_0_n190) );
  AOI22_X1 aes_state_regs_0_U50 ( .A1(aes_state_regs_0_n179), .A2(
        aes_state_regs_0_n136), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[0]), .ZN(aes_state_regs_0_n189) );
  OAI222_X1 aes_state_regs_0_U49 ( .A1(aes_state_regs_0_n188), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n197), .B2(
        aes_state_regs_0_n44), .C1(aes_state_regs_0_n180), .C2(
        aes_state_regs_0_n127), .ZN(aes_state_regs_0_S10xDN[7]) );
  INV_X1 aes_state_regs_0_U48 ( .A(aes_state_regs_0_MixColumnsS2xD[7]), .ZN(
        aes_state_regs_0_n188) );
  OAI222_X1 aes_state_regs_0_U47 ( .A1(aes_state_regs_0_n187), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n197), .B2(
        aes_state_regs_0_n45), .C1(aes_state_regs_0_n180), .C2(
        aes_state_regs_0_n126), .ZN(aes_state_regs_0_S10xDN[6]) );
  INV_X1 aes_state_regs_0_U46 ( .A(aes_state_regs_0_MixColumnsS2xD[6]), .ZN(
        aes_state_regs_0_n187) );
  OAI222_X1 aes_state_regs_0_U45 ( .A1(aes_state_regs_0_n186), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n197), .B2(
        aes_state_regs_0_n46), .C1(aes_state_regs_0_n180), .C2(
        aes_state_regs_0_n125), .ZN(aes_state_regs_0_S10xDN[5]) );
  INV_X1 aes_state_regs_0_U44 ( .A(aes_state_regs_0_MixColumnsS2xD[5]), .ZN(
        aes_state_regs_0_n186) );
  OAI222_X1 aes_state_regs_0_U43 ( .A1(aes_state_regs_0_n185), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n197), .B2(
        aes_state_regs_0_n47), .C1(aes_state_regs_0_n180), .C2(
        aes_state_regs_0_n124), .ZN(aes_state_regs_0_S10xDN[4]) );
  INV_X1 aes_state_regs_0_U42 ( .A(aes_state_regs_0_MixColumnsS2xD[4]), .ZN(
        aes_state_regs_0_n185) );
  OAI222_X1 aes_state_regs_0_U41 ( .A1(aes_state_regs_0_n184), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n197), .B2(
        aes_state_regs_0_n48), .C1(aes_state_regs_0_n180), .C2(
        aes_state_regs_0_n123), .ZN(aes_state_regs_0_S10xDN[3]) );
  INV_X1 aes_state_regs_0_U40 ( .A(aes_state_regs_0_MixColumnsS2xD[3]), .ZN(
        aes_state_regs_0_n184) );
  OAI222_X1 aes_state_regs_0_U39 ( .A1(aes_state_regs_0_n183), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n197), .B2(
        aes_state_regs_0_n49), .C1(aes_state_regs_0_n180), .C2(
        aes_state_regs_0_n122), .ZN(aes_state_regs_0_S10xDN[2]) );
  INV_X1 aes_state_regs_0_U38 ( .A(aes_state_regs_0_MixColumnsS2xD[2]), .ZN(
        aes_state_regs_0_n183) );
  OAI222_X1 aes_state_regs_0_U37 ( .A1(aes_state_regs_0_n182), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n197), .B2(
        aes_state_regs_0_n50), .C1(aes_state_regs_0_n180), .C2(
        aes_state_regs_0_n121), .ZN(aes_state_regs_0_S10xDN[1]) );
  INV_X1 aes_state_regs_0_U36 ( .A(aes_state_regs_0_MixColumnsS2xD[1]), .ZN(
        aes_state_regs_0_n182) );
  AOI22_X1 aes_state_regs_0_U35 ( .A1(aes_state_regs_0_n179), .A2(
        aes_state_regs_0_n138), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS2xD[0]), .ZN(aes_state_regs_0_n181) );
  INV_X1 aes_state_regs_0_U34 ( .A(aes_state_regs_0_n180), .ZN(
        aes_state_regs_0_n179) );
  INV_X1 aes_state_regs_0_U33 ( .A(n453), .ZN(aes_state_regs_0_n180) );
  INV_X4 aes_state_regs_0_U32 ( .A(aes_state_regs_0_n180), .ZN(
        aes_state_regs_0_n178) );
  OAI21_X1 aes_state_regs_0_U31 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n30), .A(aes_state_regs_0_n176), .ZN(StateOutxD[7])
         );
  NAND2_X1 aes_state_regs_0_U30 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[7]), .ZN(aes_state_regs_0_n176) );
  OAI21_X1 aes_state_regs_0_U29 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n29), .A(aes_state_regs_0_n175), .ZN(StateOutxD[6])
         );
  NAND2_X1 aes_state_regs_0_U28 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[6]), .ZN(aes_state_regs_0_n175) );
  OAI21_X1 aes_state_regs_0_U27 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n32), .A(aes_state_regs_0_n174), .ZN(StateOutxD[2])
         );
  NAND2_X1 aes_state_regs_0_U26 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[2]), .ZN(aes_state_regs_0_n174) );
  OAI21_X1 aes_state_regs_0_U25 ( .B1(aes_state_regs_0_n43), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n189), .ZN(
        aes_state_regs_0_S20xDN[0]) );
  OAI21_X1 aes_state_regs_0_U24 ( .B1(aes_state_regs_0_n51), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n181), .ZN(
        aes_state_regs_0_S10xDN[0]) );
  NAND2_X1 aes_state_regs_0_U23 ( .A1(doMixColumnsxS), .A2(
        aes_state_regs_0_n180), .ZN(aes_state_regs_0_n109) );
  OAI21_X1 aes_state_regs_0_U22 ( .B1(aes_state_regs_0_n42), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n190), .ZN(
        aes_state_regs_0_S20xDN[1]) );
  OAI21_X1 aes_state_regs_0_U21 ( .B1(aes_state_regs_0_n41), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n191), .ZN(
        aes_state_regs_0_S20xDN[2]) );
  OAI21_X1 aes_state_regs_0_U20 ( .B1(aes_state_regs_0_n40), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n192), .ZN(
        aes_state_regs_0_S20xDN[3]) );
  AOI22_X1 aes_state_regs_0_U19 ( .A1(aes_state_regs_0_n178), .A2(
        aes_state_regs_0_n156), .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_MixColumnsS3xD[4]), .ZN(aes_state_regs_0_n193) );
  OAI21_X1 aes_state_regs_0_U18 ( .B1(aes_state_regs_0_n39), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n193), .ZN(
        aes_state_regs_0_S20xDN[4]) );
  OAI21_X1 aes_state_regs_0_U17 ( .B1(aes_state_regs_0_n38), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n194), .ZN(
        aes_state_regs_0_S20xDN[5]) );
  OAI21_X1 aes_state_regs_0_U16 ( .B1(aes_state_regs_0_n37), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n195), .ZN(
        aes_state_regs_0_S20xDN[6]) );
  OAI21_X1 aes_state_regs_0_U15 ( .B1(aes_state_regs_0_n36), .B2(
        aes_state_regs_0_n197), .A(aes_state_regs_0_n196), .ZN(
        aes_state_regs_0_S20xDN[7]) );
  NAND2_X1 aes_state_regs_0_U14 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[5]), .ZN(aes_state_regs_0_n198) );
  OAI21_X1 aes_state_regs_0_U13 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n35), .A(aes_state_regs_0_n198), .ZN(StateOutxD[5])
         );
  NAND2_X1 aes_state_regs_0_U12 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[4]), .ZN(aes_state_regs_0_n199) );
  OAI21_X1 aes_state_regs_0_U11 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n34), .A(aes_state_regs_0_n199), .ZN(StateOutxD[4])
         );
  NAND2_X1 aes_state_regs_0_U10 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[3]), .ZN(aes_state_regs_0_n200) );
  OAI21_X1 aes_state_regs_0_U9 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n33), .A(aes_state_regs_0_n200), .ZN(StateOutxD[3])
         );
  NAND2_X1 aes_state_regs_0_U8 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[1]), .ZN(aes_state_regs_0_n201) );
  OAI21_X1 aes_state_regs_0_U7 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n31), .A(aes_state_regs_0_n201), .ZN(StateOutxD[1])
         );
  NAND2_X1 aes_state_regs_0_U6 ( .A1(aes_state_regs_0_n203), .A2(
        aes_state_regs_0_MixColumnsS0xD[0]), .ZN(aes_state_regs_0_n202) );
  OAI21_X1 aes_state_regs_0_U5 ( .B1(aes_state_regs_0_n203), .B2(
        aes_state_regs_0_n28), .A(aes_state_regs_0_n202), .ZN(StateOutxD[0])
         );
  OR2_X1 aes_state_regs_0_U4 ( .A1(aes_state_regs_0_n179), .A2(doMixColumnsxS), 
        .ZN(aes_state_regs_0_n197) );
  INV_X2 aes_state_regs_0_U3 ( .A(aes_state_regs_0_n109), .ZN(
        aes_state_regs_0_n203) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_7_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[7]), .SI(aes_state_regs_0_S10xDP_7_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[7]), .QN(aes_state_regs_0_n30) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_6_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[6]), .SI(aes_state_regs_0_S10xDP_6_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[6]), .QN(aes_state_regs_0_n29) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_5_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[5]), .SI(aes_state_regs_0_S10xDP_5_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[5]), .QN(aes_state_regs_0_n35) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_4_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[4]), .SI(aes_state_regs_0_S10xDP_4_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[4]), .QN(aes_state_regs_0_n34) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_3_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[3]), .SI(aes_state_regs_0_S10xDP_3_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[3]), .QN(aes_state_regs_0_n33) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_2_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[2]), .SI(aes_state_regs_0_S10xDP_2_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[2]), .QN(aes_state_regs_0_n32) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_1_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[1]), .SI(aes_state_regs_0_S10xDP_1_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[1]), .QN(aes_state_regs_0_n31) );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_7_ ( .D(aes_state_regs_0_S10xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_7_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_6_ ( .D(aes_state_regs_0_S10xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_6_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_5_ ( .D(aes_state_regs_0_S10xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_5_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_4_ ( .D(aes_state_regs_0_S10xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_4_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_3_ ( .D(aes_state_regs_0_S10xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_3_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_2_ ( .D(aes_state_regs_0_S10xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_2_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_1_ ( .D(aes_state_regs_0_S10xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_7_ ( .D(aes_state_regs_0_S01xDO_7_), 
        .SI(StateInxD[7]), .SE(aes_state_regs_0_n179), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_7_), .QN(aes_state_regs_0_n36) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_7_ ( .D(aes_state_regs_0_n173), .SI(
        aes_state_regs_0_n170), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[7]), .QN(aes_state_regs_0_n127) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_7_ ( .D(aes_state_regs_0_S02xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_7_ ( .D(aes_state_regs_0_n172), .SI(
        aes_state_regs_0_S23xDP_7_), .SE(aes_state_regs_0_n179), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_7_ ( .D(aes_state_regs_0_n170), .SI(
        aes_state_regs_0_n173), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_7_ ( .D(aes_state_regs_0_S02xDP_7_), 
        .SI(aes_state_regs_0_S01xDO_7_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n173), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_7_ ( .D(aes_state_regs_0_S01xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_7_ ( .D(aes_state_regs_0_S21xDP[7]), 
        .SI(aes_state_regs_0_n172), .SE(aes_state_regs_0_n179), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_7_ ( .D(aes_state_regs_0_n171), .SI(
        aes_state_regs_0_S30xDP_7_), .SE(aes_state_regs_0_n179), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n172), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_7_ ( .D(aes_state_regs_0_n169), .SI(
        aes_state_regs_0_S02xDP_7_), .SE(aes_state_regs_0_n179), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n171), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_7_ ( .D(StateInxD[7]), .SI(
        aes_state_regs_0_n169), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n170), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_7_ ( .D(aes_state_regs_0_S03xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n169), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_7_ ( .D(aes_state_regs_0_S23xDP_7_), 
        .SI(aes_state_regs_0_S20xDP_7_), .SE(aes_state_regs_0_n179), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[7]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_7_ ( .D(aes_state_regs_0_S20xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_7_), .QN(
        aes_state_regs_0_n44) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_6_ ( .D(aes_state_regs_0_S01xDO_6_), 
        .SI(StateInxD[6]), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_6_), .QN(aes_state_regs_0_n37) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_6_ ( .D(aes_state_regs_0_n168), .SI(
        aes_state_regs_0_n165), .SE(aes_state_regs_0_n179), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[6]), .QN(aes_state_regs_0_n126) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_6_ ( .D(aes_state_regs_0_S02xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_6_ ( .D(aes_state_regs_0_n167), .SI(
        aes_state_regs_0_S23xDP_6_), .SE(aes_state_regs_0_n179), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_6_ ( .D(aes_state_regs_0_n165), .SI(
        aes_state_regs_0_n168), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_6_ ( .D(aes_state_regs_0_S02xDP_6_), 
        .SI(aes_state_regs_0_S01xDO_6_), .SE(aes_state_regs_0_n179), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n168), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_6_ ( .D(aes_state_regs_0_S01xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_6_ ( .D(aes_state_regs_0_S21xDP[6]), 
        .SI(aes_state_regs_0_n167), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_6_ ( .D(aes_state_regs_0_n166), .SI(
        aes_state_regs_0_S30xDP_6_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n167), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_6_ ( .D(aes_state_regs_0_n164), .SI(
        aes_state_regs_0_S02xDP_6_), .SE(aes_state_regs_0_n179), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n166), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_6_ ( .D(StateInxD[6]), .SI(
        aes_state_regs_0_n164), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n165), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_6_ ( .D(aes_state_regs_0_S03xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n164), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_6_ ( .D(aes_state_regs_0_S23xDP_6_), 
        .SI(aes_state_regs_0_S20xDP_6_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[6]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_6_ ( .D(aes_state_regs_0_S20xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_6_), .QN(
        aes_state_regs_0_n45) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_5_ ( .D(aes_state_regs_0_S01xDO_5_), 
        .SI(StateInxD[5]), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_5_), .QN(aes_state_regs_0_n38) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_5_ ( .D(aes_state_regs_0_n163), .SI(
        aes_state_regs_0_n160), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[5]), .QN(aes_state_regs_0_n125) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_5_ ( .D(aes_state_regs_0_S02xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_5_ ( .D(aes_state_regs_0_n162), .SI(
        aes_state_regs_0_S23xDP_5_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_5_ ( .D(aes_state_regs_0_n160), .SI(
        aes_state_regs_0_n163), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_5_ ( .D(aes_state_regs_0_S02xDP_5_), 
        .SI(aes_state_regs_0_S01xDO_5_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n163), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_5_ ( .D(aes_state_regs_0_S01xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_5_ ( .D(aes_state_regs_0_S21xDP[5]), 
        .SI(aes_state_regs_0_n162), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_5_ ( .D(aes_state_regs_0_n161), .SI(
        aes_state_regs_0_S30xDP_5_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n162), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_5_ ( .D(aes_state_regs_0_n159), .SI(
        aes_state_regs_0_S02xDP_5_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n161), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_5_ ( .D(StateInxD[5]), .SI(
        aes_state_regs_0_n159), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n160), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_5_ ( .D(aes_state_regs_0_S03xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n159), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_5_ ( .D(aes_state_regs_0_S23xDP_5_), 
        .SI(aes_state_regs_0_S20xDP_5_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[5]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_5_ ( .D(aes_state_regs_0_S20xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_5_), .QN(
        aes_state_regs_0_n46) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_4_ ( .D(aes_state_regs_0_S01xDO_4_), 
        .SI(StateInxD[4]), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_4_), .QN(aes_state_regs_0_n39) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_4_ ( .D(aes_state_regs_0_n158), .SI(
        aes_state_regs_0_n155), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[4]), .QN(aes_state_regs_0_n124) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_4_ ( .D(aes_state_regs_0_S02xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_4_ ( .D(aes_state_regs_0_n157), .SI(
        aes_state_regs_0_S23xDP_4_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_4_ ( .D(aes_state_regs_0_n155), .SI(
        aes_state_regs_0_n158), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_4_ ( .D(aes_state_regs_0_S02xDP_4_), 
        .SI(aes_state_regs_0_S01xDO_4_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n158), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_4_ ( .D(aes_state_regs_0_S01xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_4_ ( .D(aes_state_regs_0_S21xDP[4]), 
        .SI(aes_state_regs_0_n157), .SE(n453), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S01xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_4_ ( .D(aes_state_regs_0_n156), .SI(
        aes_state_regs_0_S30xDP_4_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n157), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_4_ ( .D(aes_state_regs_0_n154), .SI(
        aes_state_regs_0_S02xDP_4_), .SE(n453), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_n156), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_4_ ( .D(StateInxD[4]), .SI(
        aes_state_regs_0_n154), .SE(aes_state_regs_0_n179), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n155), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_4_ ( .D(aes_state_regs_0_S03xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n154), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_4_ ( .D(aes_state_regs_0_S23xDP_4_), 
        .SI(aes_state_regs_0_S20xDP_4_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[4]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_4_ ( .D(aes_state_regs_0_S20xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_4_), .QN(
        aes_state_regs_0_n47) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_3_ ( .D(aes_state_regs_0_S01xDO_3_), 
        .SI(StateInxD[3]), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_3_), .QN(aes_state_regs_0_n40) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_3_ ( .D(aes_state_regs_0_n153), .SI(
        aes_state_regs_0_n150), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[3]), .QN(aes_state_regs_0_n123) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_3_ ( .D(aes_state_regs_0_S02xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_3_ ( .D(aes_state_regs_0_n152), .SI(
        aes_state_regs_0_S23xDP_3_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_3_ ( .D(aes_state_regs_0_n150), .SI(
        aes_state_regs_0_n153), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_3_ ( .D(aes_state_regs_0_S02xDP_3_), 
        .SI(aes_state_regs_0_S01xDO_3_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n153), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_3_ ( .D(aes_state_regs_0_S01xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_3_ ( .D(aes_state_regs_0_S21xDP[3]), 
        .SI(aes_state_regs_0_n152), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_3_ ( .D(aes_state_regs_0_n151), .SI(
        aes_state_regs_0_S30xDP_3_), .SE(aes_state_regs_0_n179), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n152), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_3_ ( .D(aes_state_regs_0_n149), .SI(
        aes_state_regs_0_S02xDP_3_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n151), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_3_ ( .D(StateInxD[3]), .SI(
        aes_state_regs_0_n149), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n150), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_3_ ( .D(aes_state_regs_0_S03xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n149), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_3_ ( .D(aes_state_regs_0_S23xDP_3_), 
        .SI(aes_state_regs_0_S20xDP_3_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[3]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_3_ ( .D(aes_state_regs_0_S20xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_3_), .QN(
        aes_state_regs_0_n48) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_2_ ( .D(aes_state_regs_0_S01xDO_2_), 
        .SI(StateInxD[2]), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_2_), .QN(aes_state_regs_0_n41) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_2_ ( .D(aes_state_regs_0_n148), .SI(
        aes_state_regs_0_n145), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[2]), .QN(aes_state_regs_0_n122) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_2_ ( .D(aes_state_regs_0_S02xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_2_ ( .D(aes_state_regs_0_n147), .SI(
        aes_state_regs_0_S23xDP_2_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_2_ ( .D(aes_state_regs_0_n145), .SI(
        aes_state_regs_0_n148), .SE(aes_state_regs_0_n179), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_2_ ( .D(aes_state_regs_0_S02xDP_2_), 
        .SI(aes_state_regs_0_S01xDO_2_), .SE(aes_state_regs_0_n179), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n148), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_2_ ( .D(aes_state_regs_0_S01xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_2_ ( .D(aes_state_regs_0_S21xDP[2]), 
        .SI(aes_state_regs_0_n147), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_2_ ( .D(aes_state_regs_0_n146), .SI(
        aes_state_regs_0_S30xDP_2_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n147), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_2_ ( .D(aes_state_regs_0_n144), .SI(
        aes_state_regs_0_S02xDP_2_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n146), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_2_ ( .D(StateInxD[2]), .SI(
        aes_state_regs_0_n144), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n145), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_2_ ( .D(aes_state_regs_0_S03xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n144), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_2_ ( .D(aes_state_regs_0_S23xDP_2_), 
        .SI(aes_state_regs_0_S20xDP_2_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[2]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_2_ ( .D(aes_state_regs_0_S20xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_2_), .QN(
        aes_state_regs_0_n49) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_1_ ( .D(aes_state_regs_0_S01xDO_1_), 
        .SI(StateInxD[1]), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_1_), .QN(aes_state_regs_0_n42) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_1_ ( .D(aes_state_regs_0_n143), .SI(
        aes_state_regs_0_n140), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[1]), .QN(aes_state_regs_0_n121) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_1_ ( .D(aes_state_regs_0_S02xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_1_ ( .D(aes_state_regs_0_n142), .SI(
        aes_state_regs_0_S23xDP_1_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_1_ ( .D(aes_state_regs_0_n140), .SI(
        aes_state_regs_0_n143), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_1_ ( .D(aes_state_regs_0_S02xDP_1_), 
        .SI(aes_state_regs_0_S01xDO_1_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n143), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_1_ ( .D(aes_state_regs_0_S01xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_1_ ( .D(aes_state_regs_0_S21xDP[1]), 
        .SI(aes_state_regs_0_n142), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_1_ ( .D(aes_state_regs_0_n141), .SI(
        aes_state_regs_0_S30xDP_1_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n142), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_1_ ( .D(aes_state_regs_0_n139), .SI(
        aes_state_regs_0_S02xDP_1_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n141), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_1_ ( .D(StateInxD[1]), .SI(
        aes_state_regs_0_n139), .SE(aes_state_regs_0_n178), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n140), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_1_ ( .D(aes_state_regs_0_S03xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n139), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_1_ ( .D(aes_state_regs_0_S23xDP_1_), 
        .SI(aes_state_regs_0_S20xDP_1_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[1]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_1_ ( .D(aes_state_regs_0_S20xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_1_), .QN(
        aes_state_regs_0_n50) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_0_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[0]), .SI(aes_state_regs_0_S10xDP_0_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[0]), .QN(aes_state_regs_0_n28) );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_0_ ( .D(aes_state_regs_0_S10xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_0_ ( .D(aes_state_regs_0_n137), .SI(
        aes_state_regs_0_S31xDP_0_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S23xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_0_ ( .D(aes_state_regs_0_S02xDP_0_), 
        .SI(aes_state_regs_0_S01xDO_0_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S31xDP_0_), .QN() );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_0_ ( .D(aes_state_regs_0_S02xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_0_ ( .D(aes_state_regs_0_S22xDP_0_), 
        .SI(aes_state_regs_0_S23xDP_0_), .SE(aes_state_regs_0_n179), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_0_ ( .D(aes_state_regs_0_n136), .SI(
        aes_state_regs_0_S30xDP_0_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S22xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_0_ ( .D(aes_state_regs_0_S01xDO_0_), 
        .SI(StateInxD[0]), .SE(aes_state_regs_0_n179), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_0_), .QN(aes_state_regs_0_n43) );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_0_ ( .D(aes_state_regs_0_S01xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_0_ ( .D(aes_state_regs_0_n138), .SI(
        aes_state_regs_0_S22xDP_0_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_0_ ( .D(aes_state_regs_0_S31xDP_0_), 
        .SI(aes_state_regs_0_n137), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n138), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_0_ ( .D(StateInxD[0]), .SI(
        aes_state_regs_0_S03xDP_0_), .SE(aes_state_regs_0_n178), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n137), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_0_ ( .D(aes_state_regs_0_S03xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_0_ ( .D(aes_state_regs_0_S23xDP_0_), 
        .SI(aes_state_regs_0_S20xDP_0_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[0]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_0_ ( .D(aes_state_regs_0_S20xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_0_), .QN(
        aes_state_regs_0_n51) );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_0_ ( .D(aes_state_regs_0_S03xDP_0_), 
        .SI(aes_state_regs_0_S02xDP_0_), .SE(aes_state_regs_0_n178), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n136), .QN() );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U119 ( .A(
        aes_state_regs_0_mix_columns_1_n245), .B(
        aes_state_regs_0_mix_columns_1_n244), .ZN(
        aes_state_regs_0_MixColumnsS3xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U118 ( .A(
        aes_state_regs_0_mix_columns_1_n240), .B(
        aes_state_regs_0_mix_columns_1_n239), .ZN(
        aes_state_regs_0_MixColumnsS3xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U117 ( .A(
        aes_state_regs_0_mix_columns_1_n235), .B(
        aes_state_regs_0_mix_columns_1_n234), .ZN(
        aes_state_regs_0_MixColumnsS3xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U116 ( .A(
        aes_state_regs_0_mix_columns_1_n226), .B(
        aes_state_regs_0_mix_columns_1_n225), .ZN(
        aes_state_regs_0_MixColumnsS3xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U115 ( .A(
        aes_state_regs_0_mix_columns_1_n183), .B(
        aes_state_regs_0_mix_columns_1_n241), .ZN(
        aes_state_regs_0_MixColumnsS1xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U114 ( .A(
        aes_state_regs_0_mix_columns_1_n190), .B(aes_state_regs_0_S00xDP[0]), 
        .ZN(aes_state_regs_0_mix_columns_1_n183) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U113 ( .A(
        aes_state_regs_0_mix_columns_1_n181), .B(
        aes_state_regs_0_mix_columns_1_n182), .ZN(
        aes_state_regs_0_MixColumnsS1xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U112 ( .A(aes_state_regs_0_S20xDP_1_), .B(aes_state_regs_0_S20xDP_2_), .ZN(aes_state_regs_0_mix_columns_1_n182) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U111 ( .A(
        aes_state_regs_0_mix_columns_1_n200), .B(aes_state_regs_0_S10xDP_1_), 
        .Z(aes_state_regs_0_mix_columns_1_n181) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U110 ( .A(
        aes_state_regs_0_mix_columns_1_n207), .B(
        aes_state_regs_0_mix_columns_1_n180), .ZN(
        aes_state_regs_0_mix_columns_1_n231) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U109 ( .A1(
        aes_state_regs_0_S30xDP_3_), .A2(aes_state_regs_0_mix_columns_1_n206), 
        .B1(aes_state_regs_0_S30xDP_7_), .B2(
        aes_state_regs_0_mix_columns_1_n179), .ZN(
        aes_state_regs_0_mix_columns_1_n180) );
  INV_X1 aes_state_regs_0_mix_columns_1_U108 ( .A(aes_state_regs_0_S30xDP_3_), 
        .ZN(aes_state_regs_0_mix_columns_1_n179) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U107 ( .A(
        aes_state_regs_0_mix_columns_1_n178), .B(
        aes_state_regs_0_mix_columns_1_n196), .ZN(
        aes_state_regs_0_MixColumnsS1xD[1]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U106 ( .A(
        aes_state_regs_0_mix_columns_1_n191), .B(aes_state_regs_0_S00xDP[1]), 
        .ZN(aes_state_regs_0_mix_columns_1_n178) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U105 ( .A(
        aes_state_regs_0_mix_columns_1_n177), .B(
        aes_state_regs_0_mix_columns_1_n203), .ZN(
        aes_state_regs_0_MixColumnsS1xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U104 ( .A(aes_state_regs_0_S20xDP_3_), .B(aes_state_regs_0_mix_columns_1_n192), .ZN(
        aes_state_regs_0_mix_columns_1_n177) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U103 ( .A(
        aes_state_regs_0_mix_columns_1_n176), .B(
        aes_state_regs_0_mix_columns_1_n205), .ZN(
        aes_state_regs_0_MixColumnsS1xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U102 ( .A(
        aes_state_regs_0_mix_columns_1_n193), .B(aes_state_regs_0_S00xDP[4]), 
        .ZN(aes_state_regs_0_mix_columns_1_n176) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U101 ( .A1(
        aes_state_regs_0_S30xDP_2_), .A2(aes_state_regs_0_S30xDP_7_), .B1(
        aes_state_regs_0_mix_columns_1_n206), .B2(
        aes_state_regs_0_mix_columns_1_n175), .ZN(
        aes_state_regs_0_mix_columns_1_n228) );
  INV_X1 aes_state_regs_0_mix_columns_1_U100 ( .A(aes_state_regs_0_S30xDP_2_), 
        .ZN(aes_state_regs_0_mix_columns_1_n175) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U99 ( .A(
        aes_state_regs_0_mix_columns_1_n173), .B(
        aes_state_regs_0_mix_columns_1_n174), .ZN(
        aes_state_regs_0_MixColumnsS1xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U98 ( .A(aes_state_regs_0_S20xDP_4_), 
        .B(aes_state_regs_0_mix_columns_1_n211), .ZN(
        aes_state_regs_0_mix_columns_1_n174) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U97 ( .A(aes_state_regs_0_S00xDP[5]), 
        .B(aes_state_regs_0_S10xDP_4_), .Z(aes_state_regs_0_mix_columns_1_n173) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U96 ( .A(
        aes_state_regs_0_mix_columns_1_n171), .B(
        aes_state_regs_0_mix_columns_1_n172), .ZN(
        aes_state_regs_0_MixColumnsS1xD[7]) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U95 ( .A1(aes_state_regs_0_S20xDP_6_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n236), .ZN(
        aes_state_regs_0_mix_columns_1_n172) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U94 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n217), .ZN(
        aes_state_regs_0_mix_columns_1_n171) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U93 ( .A(
        aes_state_regs_0_mix_columns_1_n169), .B(
        aes_state_regs_0_mix_columns_1_n170), .ZN(
        aes_state_regs_0_MixColumnsS1xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U92 ( .A(aes_state_regs_0_S20xDP_5_), 
        .B(aes_state_regs_0_mix_columns_1_n215), .ZN(
        aes_state_regs_0_mix_columns_1_n170) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U91 ( .A(aes_state_regs_0_S00xDP[6]), 
        .B(aes_state_regs_0_S10xDP_5_), .Z(aes_state_regs_0_mix_columns_1_n169) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U90 ( .A1(aes_state_regs_0_S20xDP_3_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n168), .ZN(
        aes_state_regs_0_mix_columns_1_n205) );
  INV_X1 aes_state_regs_0_mix_columns_1_U89 ( .A(aes_state_regs_0_S20xDP_3_), 
        .ZN(aes_state_regs_0_mix_columns_1_n168) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U88 ( .A(
        aes_state_regs_0_mix_columns_1_n167), .B(
        aes_state_regs_0_mix_columns_1_n209), .ZN(
        aes_state_regs_0_mix_columns_1_n193) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U87 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_3_), .ZN(
        aes_state_regs_0_mix_columns_1_n167) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U86 ( .A(
        aes_state_regs_0_mix_columns_1_n165), .B(
        aes_state_regs_0_mix_columns_1_n166), .ZN(
        aes_state_regs_0_mix_columns_1_n227) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U85 ( .A(aes_state_regs_0_S20xDP_3_), 
        .B(aes_state_regs_0_S10xDP_3_), .ZN(
        aes_state_regs_0_mix_columns_1_n166) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U84 ( .A(aes_state_regs_0_S00xDP[2]), 
        .B(aes_state_regs_0_S00xDP[7]), .Z(aes_state_regs_0_mix_columns_1_n165) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U83 ( .A(
        aes_state_regs_0_mix_columns_1_n164), .B(
        aes_state_regs_0_mix_columns_1_n163), .ZN(
        aes_state_regs_0_mix_columns_1_n203) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U82 ( .A(aes_state_regs_0_S20xDP_2_), 
        .B(aes_state_regs_0_S30xDP_3_), .ZN(
        aes_state_regs_0_mix_columns_1_n164) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U81 ( .A1(aes_state_regs_0_S00xDP[3]), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n162), .ZN(
        aes_state_regs_0_mix_columns_1_n163) );
  INV_X1 aes_state_regs_0_mix_columns_1_U80 ( .A(aes_state_regs_0_S00xDP[3]), 
        .ZN(aes_state_regs_0_mix_columns_1_n162) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U79 ( .A(
        aes_state_regs_0_mix_columns_1_n161), .B(aes_state_regs_0_S30xDP_7_), 
        .ZN(aes_state_regs_0_MixColumnsS0xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U78 ( .A(
        aes_state_regs_0_mix_columns_1_n241), .B(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_mix_columns_1_n161) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U77 ( .A(
        aes_state_regs_0_mix_columns_1_n160), .B(
        aes_state_regs_0_mix_columns_1_n215), .ZN(
        aes_state_regs_0_MixColumnsS0xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U76 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n233), .ZN(
        aes_state_regs_0_mix_columns_1_n160) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U75 ( .A(
        aes_state_regs_0_mix_columns_1_n159), .B(
        aes_state_regs_0_mix_columns_1_n198), .ZN(
        aes_state_regs_0_MixColumnsS0xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U74 ( .A(aes_state_regs_0_S30xDP_2_), 
        .B(aes_state_regs_0_mix_columns_1_n224), .ZN(
        aes_state_regs_0_mix_columns_1_n159) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U73 ( .A1(aes_state_regs_0_S20xDP_0_), .A2(aes_state_regs_0_mix_columns_1_n218), .B1(
        aes_state_regs_0_mix_columns_1_n217), .B2(
        aes_state_regs_0_mix_columns_1_n216), .ZN(
        aes_state_regs_0_mix_columns_1_n219) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U72 ( .A(
        aes_state_regs_0_mix_columns_1_n220), .B(
        aes_state_regs_0_mix_columns_1_n219), .ZN(
        aes_state_regs_0_MixColumnsS3xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U71 ( .A(aes_state_regs_0_S20xDP_7_), 
        .B(aes_state_regs_0_mix_columns_1_n197), .ZN(
        aes_state_regs_0_mix_columns_1_n195) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U70 ( .A(
        aes_state_regs_0_mix_columns_1_n195), .B(
        aes_state_regs_0_mix_columns_1_n220), .ZN(
        aes_state_regs_0_MixColumnsS2xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U69 ( .A(
        aes_state_regs_0_mix_columns_1_n221), .B(aes_state_regs_0_S20xDP_1_), 
        .ZN(aes_state_regs_0_mix_columns_1_n223) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U68 ( .A(
        aes_state_regs_0_mix_columns_1_n223), .B(
        aes_state_regs_0_mix_columns_1_n222), .ZN(
        aes_state_regs_0_MixColumnsS3xD[1]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U67 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n224), .ZN(
        aes_state_regs_0_mix_columns_1_n225) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U66 ( .A(aes_state_regs_0_S00xDP[2]), 
        .B(aes_state_regs_0_S00xDP[1]), .Z(aes_state_regs_0_mix_columns_1_n226) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U65 ( .A(
        aes_state_regs_0_mix_columns_1_n227), .B(aes_state_regs_0_S00xDP[3]), 
        .ZN(aes_state_regs_0_mix_columns_1_n229) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U64 ( .A(
        aes_state_regs_0_mix_columns_1_n229), .B(
        aes_state_regs_0_mix_columns_1_n228), .ZN(
        aes_state_regs_0_MixColumnsS3xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U63 ( .A(
        aes_state_regs_0_mix_columns_1_n230), .B(aes_state_regs_0_S20xDP_4_), 
        .ZN(aes_state_regs_0_mix_columns_1_n232) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U62 ( .A(
        aes_state_regs_0_mix_columns_1_n232), .B(
        aes_state_regs_0_mix_columns_1_n231), .ZN(
        aes_state_regs_0_MixColumnsS3xD[4]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U61 ( .A(
        aes_state_regs_0_mix_columns_1_n233), .B(aes_state_regs_0_S20xDP_5_), 
        .Z(aes_state_regs_0_mix_columns_1_n235) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U60 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_S00xDP[4]), .ZN(
        aes_state_regs_0_mix_columns_1_n234) );
  INV_X1 aes_state_regs_0_mix_columns_1_U59 ( .A(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_mix_columns_1_n237) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U58 ( .A1(aes_state_regs_0_S20xDP_6_), .A2(aes_state_regs_0_mix_columns_1_n238), .B1(
        aes_state_regs_0_mix_columns_1_n237), .B2(
        aes_state_regs_0_mix_columns_1_n236), .ZN(
        aes_state_regs_0_mix_columns_1_n239) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U57 ( .A(aes_state_regs_0_S30xDP_5_), 
        .B(aes_state_regs_0_S00xDP[5]), .ZN(
        aes_state_regs_0_mix_columns_1_n240) );
  INV_X1 aes_state_regs_0_mix_columns_1_U56 ( .A(aes_state_regs_0_S00xDP[6]), 
        .ZN(aes_state_regs_0_mix_columns_1_n243) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U55 ( .A(aes_state_regs_0_S30xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n241), .ZN(
        aes_state_regs_0_mix_columns_1_n245) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U54 ( .A1(aes_state_regs_0_S00xDP[7]), .A2(aes_state_regs_0_S00xDP[6]), .B1(aes_state_regs_0_mix_columns_1_n243), 
        .B2(aes_state_regs_0_mix_columns_1_n242), .ZN(
        aes_state_regs_0_mix_columns_1_n244) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U53 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n196), .ZN(
        aes_state_regs_0_mix_columns_1_n199) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U52 ( .A(
        aes_state_regs_0_mix_columns_1_n199), .B(
        aes_state_regs_0_mix_columns_1_n222), .ZN(
        aes_state_regs_0_MixColumnsS2xD[1]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U51 ( .A(aes_state_regs_0_S10xDP_2_), 
        .B(aes_state_regs_0_mix_columns_1_n200), .Z(
        aes_state_regs_0_mix_columns_1_n201) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U50 ( .A(
        aes_state_regs_0_mix_columns_1_n202), .B(
        aes_state_regs_0_mix_columns_1_n201), .ZN(
        aes_state_regs_0_MixColumnsS2xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U49 ( .A(aes_state_regs_0_S10xDP_3_), 
        .B(aes_state_regs_0_mix_columns_1_n203), .ZN(
        aes_state_regs_0_mix_columns_1_n204) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U48 ( .A(
        aes_state_regs_0_mix_columns_1_n204), .B(
        aes_state_regs_0_mix_columns_1_n228), .ZN(
        aes_state_regs_0_MixColumnsS2xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U47 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_mix_columns_1_n205), .ZN(
        aes_state_regs_0_mix_columns_1_n208) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U46 ( .A(
        aes_state_regs_0_mix_columns_1_n208), .B(
        aes_state_regs_0_mix_columns_1_n231), .ZN(
        aes_state_regs_0_MixColumnsS2xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U45 ( .A(
        aes_state_regs_0_mix_columns_1_n209), .B(aes_state_regs_0_S30xDP_5_), 
        .ZN(aes_state_regs_0_mix_columns_1_n210) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U44 ( .A(
        aes_state_regs_0_mix_columns_1_n210), .B(
        aes_state_regs_0_mix_columns_1_n233), .ZN(
        aes_state_regs_0_MixColumnsS2xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U43 ( .A(
        aes_state_regs_0_mix_columns_1_n211), .B(aes_state_regs_0_S30xDP_6_), 
        .ZN(aes_state_regs_0_mix_columns_1_n212) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U42 ( .A(
        aes_state_regs_0_mix_columns_1_n212), .B(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_MixColumnsS2xD[6]) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U41 ( .A1(aes_state_regs_0_S10xDP_7_), .A2(aes_state_regs_0_mix_columns_1_n218), .B1(
        aes_state_regs_0_mix_columns_1_n217), .B2(
        aes_state_regs_0_mix_columns_1_n213), .ZN(
        aes_state_regs_0_mix_columns_1_n214) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U40 ( .A(
        aes_state_regs_0_mix_columns_1_n215), .B(
        aes_state_regs_0_mix_columns_1_n214), .ZN(
        aes_state_regs_0_MixColumnsS2xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U39 ( .A(aes_state_regs_0_S10xDP_5_), 
        .B(aes_state_regs_0_mix_columns_1_n207), .ZN(
        aes_state_regs_0_mix_columns_1_n189) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U38 ( .A(
        aes_state_regs_0_mix_columns_1_n189), .B(
        aes_state_regs_0_mix_columns_1_n211), .ZN(
        aes_state_regs_0_MixColumnsS0xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U37 ( .A(aes_state_regs_0_S10xDP_4_), 
        .B(aes_state_regs_0_mix_columns_1_n230), .ZN(
        aes_state_regs_0_mix_columns_1_n188) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U36 ( .A(
        aes_state_regs_0_mix_columns_1_n188), .B(
        aes_state_regs_0_mix_columns_1_n193), .ZN(
        aes_state_regs_0_MixColumnsS0xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U35 ( .A(aes_state_regs_0_S30xDP_3_), 
        .B(aes_state_regs_0_mix_columns_1_n227), .ZN(
        aes_state_regs_0_mix_columns_1_n187) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U34 ( .A(
        aes_state_regs_0_mix_columns_1_n187), .B(
        aes_state_regs_0_mix_columns_1_n192), .ZN(
        aes_state_regs_0_MixColumnsS0xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U33 ( .A(aes_state_regs_0_S10xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n221), .ZN(
        aes_state_regs_0_mix_columns_1_n186) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U32 ( .A(
        aes_state_regs_0_mix_columns_1_n186), .B(
        aes_state_regs_0_mix_columns_1_n191), .ZN(
        aes_state_regs_0_MixColumnsS0xD[1]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U31 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_mix_columns_1_n185), .ZN(
        aes_state_regs_0_mix_columns_1_n184) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U30 ( .A(
        aes_state_regs_0_mix_columns_1_n184), .B(
        aes_state_regs_0_mix_columns_1_n190), .ZN(
        aes_state_regs_0_MixColumnsS0xD[0]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U29 ( .A(aes_state_regs_0_S10xDP_0_), 
        .B(aes_state_regs_0_S00xDP[0]), .Z(aes_state_regs_0_mix_columns_1_n220) );
  INV_X1 aes_state_regs_0_mix_columns_1_U28 ( .A(
        aes_state_regs_0_mix_columns_1_n217), .ZN(
        aes_state_regs_0_mix_columns_1_n218) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U27 ( .A1(aes_state_regs_0_S00xDP[7]), .A2(aes_state_regs_0_S30xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n206), 
        .B2(aes_state_regs_0_mix_columns_1_n242), .ZN(
        aes_state_regs_0_mix_columns_1_n217) );
  INV_X1 aes_state_regs_0_mix_columns_1_U26 ( .A(aes_state_regs_0_S20xDP_0_), 
        .ZN(aes_state_regs_0_mix_columns_1_n216) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U25 ( .A(aes_state_regs_0_S30xDP_0_), 
        .B(aes_state_regs_0_mix_columns_1_n206), .ZN(
        aes_state_regs_0_mix_columns_1_n197) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U24 ( .A(aes_state_regs_0_S30xDP_0_), 
        .B(aes_state_regs_0_S20xDP_0_), .Z(aes_state_regs_0_mix_columns_1_n190) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U23 ( .A1(aes_state_regs_0_S10xDP_7_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n213), .ZN(
        aes_state_regs_0_mix_columns_1_n241) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U22 ( .A(
        aes_state_regs_0_mix_columns_1_n198), .B(
        aes_state_regs_0_mix_columns_1_n197), .Z(
        aes_state_regs_0_mix_columns_1_n222) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U21 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_S00xDP[0]), .Z(aes_state_regs_0_mix_columns_1_n221) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U20 ( .A(aes_state_regs_0_S10xDP_2_), 
        .B(aes_state_regs_0_S20xDP_2_), .Z(aes_state_regs_0_mix_columns_1_n224) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U19 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_S00xDP[3]), .Z(aes_state_regs_0_mix_columns_1_n230) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U18 ( .A(aes_state_regs_0_S10xDP_5_), 
        .B(aes_state_regs_0_S00xDP[5]), .Z(aes_state_regs_0_mix_columns_1_n233) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U17 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_S00xDP[6]), .Z(aes_state_regs_0_mix_columns_1_n238) );
  INV_X1 aes_state_regs_0_mix_columns_1_U16 ( .A(aes_state_regs_0_S20xDP_6_), 
        .ZN(aes_state_regs_0_mix_columns_1_n236) );
  INV_X1 aes_state_regs_0_mix_columns_1_U15 ( .A(aes_state_regs_0_S00xDP[7]), 
        .ZN(aes_state_regs_0_mix_columns_1_n242) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U14 ( .A1(aes_state_regs_0_S20xDP_0_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n216), .ZN(
        aes_state_regs_0_mix_columns_1_n196) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U13 ( .A(aes_state_regs_0_S30xDP_2_), 
        .B(aes_state_regs_0_S00xDP[2]), .Z(aes_state_regs_0_mix_columns_1_n200) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U12 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_S20xDP_1_), .ZN(
        aes_state_regs_0_mix_columns_1_n202) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U11 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_S20xDP_4_), .Z(aes_state_regs_0_mix_columns_1_n209) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U10 ( .A(aes_state_regs_0_S30xDP_5_), 
        .B(aes_state_regs_0_S20xDP_5_), .Z(aes_state_regs_0_mix_columns_1_n211) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U9 ( .A(aes_state_regs_0_S30xDP_6_), 
        .B(aes_state_regs_0_S20xDP_6_), .Z(aes_state_regs_0_mix_columns_1_n215) );
  INV_X1 aes_state_regs_0_mix_columns_1_U8 ( .A(aes_state_regs_0_S10xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n213) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U7 ( .A(
        aes_state_regs_0_mix_columns_1_n185), .B(
        aes_state_regs_0_mix_columns_1_n202), .ZN(
        aes_state_regs_0_mix_columns_1_n191) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U6 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_2_), .Z(aes_state_regs_0_mix_columns_1_n192) );
  INV_X1 aes_state_regs_0_mix_columns_1_U5 ( .A(aes_state_regs_0_S20xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n194) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U4 ( .A(aes_state_regs_0_S10xDP_4_), 
        .B(aes_state_regs_0_S00xDP[4]), .Z(aes_state_regs_0_mix_columns_1_n207) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U3 ( .A(aes_state_regs_0_S10xDP_1_), 
        .B(aes_state_regs_0_S00xDP[1]), .Z(aes_state_regs_0_mix_columns_1_n198) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U2 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_0_), .Z(aes_state_regs_0_mix_columns_1_n185) );
  INV_X1 aes_state_regs_0_mix_columns_1_U1 ( .A(aes_state_regs_0_S30xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n206) );
endmodule

