module circuit ( clk, rst, en, enc, p0, p1, r, k, c0, c1, done );
  input [63:0] p0;
  input [63:0] p1;
  input [127:0] r;
  input [127:0] k;
  output [63:0] c0;
  output [63:0] c1;
  input clk, rst, en, enc;
  output done;
  wire   en_sig, start_sig, inv_sig, inv_sig2, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, reg_k0_n340, reg_k0_n339, reg_k0_n338, reg_k0_n337,
         reg_k0_n336, reg_k0_n335, reg_k0_n334, reg_k0_n333, reg_k0_n332,
         reg_k0_n331, reg_k0_n330, reg_k0_n329, reg_k0_n328, reg_k0_n327,
         reg_k0_n326, reg_k0_n325, reg_k0_n324, reg_k0_n323, reg_k0_n322,
         reg_k0_n321, reg_k0_n320, reg_k0_n319, reg_k0_n318, reg_k0_n317,
         reg_k0_n316, reg_k0_n315, reg_k0_n314, reg_k0_n313, reg_k0_n312,
         reg_k0_n311, reg_k0_n310, reg_k0_n309, reg_k0_n308, reg_k0_n307,
         reg_k0_n306, reg_k0_n305, reg_k0_n304, reg_k0_n303, reg_k0_n302,
         reg_k0_n301, reg_k0_n300, reg_k0_n299, reg_k0_n298, reg_k0_n297,
         reg_k0_n296, reg_k0_n295, reg_k0_n294, reg_k0_n293, reg_k0_n292,
         reg_k0_n291, reg_k0_n290, reg_k0_n289, reg_k0_n288, reg_k0_n287,
         reg_k0_n286, reg_k0_n285, reg_k0_n284, reg_k0_n283, reg_k0_n282,
         reg_k0_n281, reg_k0_n280, reg_k0_n279, reg_k0_n278, reg_k0_n277,
         reg_k0_n276, reg_k0_n275, reg_k0_n274, reg_k0_n273, reg_k0_n272,
         reg_k0_n271, reg_k0_n270, reg_k0_n269, reg_k0_n268, reg_k0_n267,
         reg_k0_n266, reg_k0_n265, reg_k0_n264, reg_k0_n263, reg_k0_n262,
         reg_k0_n261, reg_k0_n260, reg_k0_n259, reg_k0_n258, reg_k0_n257,
         reg_k0_n256, reg_k0_n255, reg_k0_n254, reg_k0_n253, reg_k0_n252,
         reg_k0_n251, reg_k0_n250, reg_k0_n249, reg_k0_n248, reg_k0_n247,
         reg_k0_n246, reg_k0_n245, reg_k0_n244, reg_k0_n243, reg_k0_n242,
         reg_k0_n241, reg_k0_n240, reg_k0_n239, reg_k0_n238, reg_k0_n237,
         reg_k0_n236, reg_k0_n235, reg_k0_n234, reg_k0_n233, reg_k0_n232,
         reg_k0_n231, reg_k0_n230, reg_k0_n229, reg_k0_n228, reg_k0_n227,
         reg_k0_n226, reg_k0_n225, reg_k0_n224, reg_k0_n223, reg_k0_n222,
         reg_k0_n221, reg_k0_n220, reg_k0_n219, reg_k0_n218, reg_k0_n217,
         reg_k0_n216, reg_k0_n215, reg_k0_n214, reg_k0_n213, reg_k0_n212,
         reg_k0_n211, reg_k0_n210, reg_k0_n209, reg_k0_n208, reg_k0_n207,
         reg_k0_n206, reg_k0_n205, reg_k0_n204, reg_k0_n203, reg_k0_n202,
         reg_k0_n195, reg_k0_n194, reg_k0_n193, reg_k0_n192, reg_k0_n191,
         reg_k0_n190, reg_k0_n189, reg_k0_n188, reg_k0_n187, reg_k0_n186,
         reg_k0_n185, reg_k0_n184, reg_k0_n183, reg_k0_n182, reg_k0_n181,
         reg_k0_n180, reg_k0_n179, reg_k0_n178, reg_k0_n177, reg_k0_n176,
         reg_k0_n175, reg_k0_n174, reg_k0_n173, reg_k0_n172, reg_k0_n171,
         reg_k0_n170, reg_k0_n169, reg_k0_n168, reg_k0_n167, reg_k0_n166,
         reg_k0_n165, reg_k0_n164, reg_k0_n163, reg_k0_n162, reg_k0_n161,
         reg_k0_n160, reg_k0_n159, reg_k0_n158, reg_k0_n157, reg_k0_n156,
         reg_k0_n155, reg_k0_n154, reg_k0_n153, reg_k0_n152, reg_k0_n151,
         reg_k0_n150, reg_k0_n149, reg_k0_n148, reg_k0_n147, reg_k0_n146,
         reg_k0_n145, reg_k0_n144, reg_k0_n143, reg_k0_n142, reg_k0_n141,
         reg_k0_n140, reg_k0_n139, reg_k0_n138, reg_k0_n137, reg_k0_n136,
         reg_k0_n135, reg_k0_n134, reg_k0_n133, reg_k0_n132, reg_k1_n532,
         reg_k1_n531, reg_k1_n530, reg_k1_n529, reg_k1_n528, reg_k1_n527,
         reg_k1_n526, reg_k1_n525, reg_k1_n524, reg_k1_n523, reg_k1_n522,
         reg_k1_n521, reg_k1_n520, reg_k1_n519, reg_k1_n518, reg_k1_n517,
         reg_k1_n516, reg_k1_n515, reg_k1_n514, reg_k1_n513, reg_k1_n512,
         reg_k1_n511, reg_k1_n510, reg_k1_n509, reg_k1_n508, reg_k1_n507,
         reg_k1_n506, reg_k1_n505, reg_k1_n504, reg_k1_n503, reg_k1_n502,
         reg_k1_n501, reg_k1_n500, reg_k1_n499, reg_k1_n498, reg_k1_n497,
         reg_k1_n496, reg_k1_n495, reg_k1_n494, reg_k1_n493, reg_k1_n492,
         reg_k1_n491, reg_k1_n490, reg_k1_n489, reg_k1_n488, reg_k1_n487,
         reg_k1_n486, reg_k1_n485, reg_k1_n484, reg_k1_n483, reg_k1_n482,
         reg_k1_n481, reg_k1_n480, reg_k1_n479, reg_k1_n478, reg_k1_n477,
         reg_k1_n476, reg_k1_n475, reg_k1_n474, reg_k1_n473, reg_k1_n472,
         reg_k1_n471, reg_k1_n470, reg_k1_n469, reg_k1_n468, reg_k1_n467,
         reg_k1_n466, reg_k1_n465, reg_k1_n464, reg_k1_n463, reg_k1_n462,
         reg_k1_n461, reg_k1_n460, reg_k1_n459, reg_k1_n458, reg_k1_n457,
         reg_k1_n456, reg_k1_n455, reg_k1_n454, reg_k1_n453, reg_k1_n452,
         reg_k1_n451, reg_k1_n450, reg_k1_n449, reg_k1_n448, reg_k1_n447,
         reg_k1_n446, reg_k1_n445, reg_k1_n444, reg_k1_n443, reg_k1_n442,
         reg_k1_n441, reg_k1_n440, reg_k1_n439, reg_k1_n438, reg_k1_n437,
         reg_k1_n436, reg_k1_n435, reg_k1_n434, reg_k1_n433, reg_k1_n432,
         reg_k1_n431, reg_k1_n430, reg_k1_n429, reg_k1_n428, reg_k1_n427,
         reg_k1_n426, reg_k1_n425, reg_k1_n424, reg_k1_n423, reg_k1_n422,
         reg_k1_n421, reg_k1_n420, reg_k1_n419, reg_k1_n418, reg_k1_n417,
         reg_k1_n416, reg_k1_n415, reg_k1_n414, reg_k1_n413, reg_k1_n412,
         reg_k1_n411, reg_k1_n410, reg_k1_n409, reg_k1_n408, reg_k1_n407,
         reg_k1_n406, reg_k1_n405, reg_k1_n404, reg_k1_n403, reg_k1_n402,
         reg_k1_n401, reg_k1_n400, reg_k1_n399, reg_k1_n398, reg_k1_n397,
         reg_k1_n396, reg_k1_n395, reg_k1_n394, reg_k1_n265, reg_k1_n264,
         reg_k1_n263, reg_k1_n262, reg_k1_n261, reg_k1_n260, reg_k1_n259,
         reg_k1_n258, reg_k1_n257, reg_k1_n256, reg_k1_n255, reg_k1_n254,
         reg_k1_n253, reg_k1_n252, reg_k1_n251, reg_k1_n250, reg_k1_n249,
         reg_k1_n248, reg_k1_n247, reg_k1_n246, reg_k1_n245, reg_k1_n244,
         reg_k1_n243, reg_k1_n242, reg_k1_n241, reg_k1_n240, reg_k1_n239,
         reg_k1_n238, reg_k1_n237, reg_k1_n236, reg_k1_n235, reg_k1_n234,
         reg_k1_n233, reg_k1_n232, reg_k1_n231, reg_k1_n230, reg_k1_n229,
         reg_k1_n228, reg_k1_n227, reg_k1_n226, reg_k1_n225, reg_k1_n224,
         reg_k1_n223, reg_k1_n222, reg_k1_n221, reg_k1_n220, reg_k1_n219,
         reg_k1_n218, reg_k1_n217, reg_k1_n216, reg_k1_n215, reg_k1_n214,
         reg_k1_n213, reg_k1_n212, reg_k1_n211, reg_k1_n210, reg_k1_n209,
         reg_k1_n208, reg_k1_n207, reg_k1_n206, reg_k1_n205, reg_k1_n204,
         reg_k1_n203, reg_k1_n202, reg_p0_n531, reg_p0_n530, reg_p0_n529,
         reg_p0_n528, reg_p0_n527, reg_p0_n526, reg_p0_n525, reg_p0_n524,
         reg_p0_n523, reg_p0_n522, reg_p0_n521, reg_p0_n520, reg_p0_n519,
         reg_p0_n518, reg_p0_n517, reg_p0_n516, reg_p0_n515, reg_p0_n514,
         reg_p0_n513, reg_p0_n512, reg_p0_n511, reg_p0_n510, reg_p0_n509,
         reg_p0_n508, reg_p0_n507, reg_p0_n506, reg_p0_n505, reg_p0_n504,
         reg_p0_n503, reg_p0_n502, reg_p0_n501, reg_p0_n500, reg_p0_n499,
         reg_p0_n498, reg_p0_n497, reg_p0_n496, reg_p0_n495, reg_p0_n494,
         reg_p0_n493, reg_p0_n492, reg_p0_n491, reg_p0_n490, reg_p0_n489,
         reg_p0_n488, reg_p0_n487, reg_p0_n486, reg_p0_n485, reg_p0_n484,
         reg_p0_n483, reg_p0_n482, reg_p0_n481, reg_p0_n480, reg_p0_n479,
         reg_p0_n478, reg_p0_n477, reg_p0_n476, reg_p0_n475, reg_p0_n474,
         reg_p0_n473, reg_p0_n472, reg_p0_n471, reg_p0_n470, reg_p0_n469,
         reg_p0_n468, reg_p0_n467, reg_p0_n466, reg_p0_n465, reg_p0_n464,
         reg_p0_n463, reg_p0_n462, reg_p0_n461, reg_p0_n460, reg_p0_n459,
         reg_p0_n458, reg_p0_n457, reg_p0_n456, reg_p0_n455, reg_p0_n454,
         reg_p0_n453, reg_p0_n452, reg_p0_n451, reg_p0_n450, reg_p0_n449,
         reg_p0_n448, reg_p0_n447, reg_p0_n446, reg_p0_n445, reg_p0_n444,
         reg_p0_n443, reg_p0_n442, reg_p0_n441, reg_p0_n440, reg_p0_n439,
         reg_p0_n438, reg_p0_n437, reg_p0_n436, reg_p0_n435, reg_p0_n434,
         reg_p0_n433, reg_p0_n432, reg_p0_n431, reg_p0_n430, reg_p0_n429,
         reg_p0_n428, reg_p0_n427, reg_p0_n426, reg_p0_n425, reg_p0_n424,
         reg_p0_n423, reg_p0_n422, reg_p0_n421, reg_p0_n420, reg_p0_n419,
         reg_p0_n418, reg_p0_n417, reg_p0_n416, reg_p0_n415, reg_p0_n414,
         reg_p0_n413, reg_p0_n412, reg_p0_n411, reg_p0_n410, reg_p0_n409,
         reg_p0_n408, reg_p0_n407, reg_p0_n406, reg_p0_n405, reg_p0_n404,
         reg_p0_n403, reg_p0_n402, reg_p0_n401, reg_p0_n400, reg_p0_n399,
         reg_p0_n398, reg_p0_n397, reg_p0_n396, reg_p0_n395, reg_p0_n394,
         reg_p0_n265, reg_p0_n264, reg_p0_n263, reg_p0_n262, reg_p0_n261,
         reg_p0_n260, reg_p0_n259, reg_p0_n258, reg_p0_n257, reg_p0_n256,
         reg_p0_n255, reg_p0_n254, reg_p0_n253, reg_p0_n252, reg_p0_n251,
         reg_p0_n250, reg_p0_n249, reg_p0_n248, reg_p0_n247, reg_p0_n246,
         reg_p0_n245, reg_p0_n244, reg_p0_n243, reg_p0_n242, reg_p0_n241,
         reg_p0_n240, reg_p0_n239, reg_p0_n238, reg_p0_n237, reg_p0_n236,
         reg_p0_n235, reg_p0_n234, reg_p0_n233, reg_p0_n232, reg_p0_n231,
         reg_p0_n230, reg_p0_n229, reg_p0_n228, reg_p0_n227, reg_p0_n226,
         reg_p0_n225, reg_p0_n224, reg_p0_n223, reg_p0_n222, reg_p0_n221,
         reg_p0_n220, reg_p0_n219, reg_p0_n218, reg_p0_n217, reg_p0_n216,
         reg_p0_n215, reg_p0_n214, reg_p0_n213, reg_p0_n212, reg_p0_n211,
         reg_p0_n210, reg_p0_n209, reg_p0_n208, reg_p0_n207, reg_p0_n206,
         reg_p0_n205, reg_p0_n204, reg_p0_n203, reg_p0_n202, reg_p1_n532,
         reg_p1_n531, reg_p1_n530, reg_p1_n529, reg_p1_n528, reg_p1_n527,
         reg_p1_n526, reg_p1_n525, reg_p1_n524, reg_p1_n523, reg_p1_n522,
         reg_p1_n521, reg_p1_n520, reg_p1_n519, reg_p1_n518, reg_p1_n517,
         reg_p1_n516, reg_p1_n515, reg_p1_n514, reg_p1_n513, reg_p1_n512,
         reg_p1_n511, reg_p1_n510, reg_p1_n509, reg_p1_n508, reg_p1_n507,
         reg_p1_n506, reg_p1_n505, reg_p1_n504, reg_p1_n503, reg_p1_n502,
         reg_p1_n501, reg_p1_n500, reg_p1_n499, reg_p1_n498, reg_p1_n497,
         reg_p1_n496, reg_p1_n495, reg_p1_n494, reg_p1_n493, reg_p1_n492,
         reg_p1_n491, reg_p1_n490, reg_p1_n489, reg_p1_n488, reg_p1_n487,
         reg_p1_n486, reg_p1_n485, reg_p1_n484, reg_p1_n483, reg_p1_n482,
         reg_p1_n481, reg_p1_n480, reg_p1_n479, reg_p1_n478, reg_p1_n477,
         reg_p1_n476, reg_p1_n475, reg_p1_n474, reg_p1_n473, reg_p1_n472,
         reg_p1_n471, reg_p1_n470, reg_p1_n469, reg_p1_n468, reg_p1_n467,
         reg_p1_n466, reg_p1_n465, reg_p1_n464, reg_p1_n463, reg_p1_n462,
         reg_p1_n461, reg_p1_n460, reg_p1_n459, reg_p1_n458, reg_p1_n457,
         reg_p1_n456, reg_p1_n455, reg_p1_n454, reg_p1_n453, reg_p1_n452,
         reg_p1_n451, reg_p1_n450, reg_p1_n449, reg_p1_n448, reg_p1_n447,
         reg_p1_n446, reg_p1_n445, reg_p1_n444, reg_p1_n443, reg_p1_n442,
         reg_p1_n441, reg_p1_n440, reg_p1_n439, reg_p1_n438, reg_p1_n437,
         reg_p1_n436, reg_p1_n435, reg_p1_n434, reg_p1_n433, reg_p1_n432,
         reg_p1_n431, reg_p1_n430, reg_p1_n429, reg_p1_n428, reg_p1_n427,
         reg_p1_n426, reg_p1_n425, reg_p1_n424, reg_p1_n423, reg_p1_n422,
         reg_p1_n421, reg_p1_n420, reg_p1_n419, reg_p1_n418, reg_p1_n417,
         reg_p1_n416, reg_p1_n415, reg_p1_n414, reg_p1_n413, reg_p1_n412,
         reg_p1_n411, reg_p1_n410, reg_p1_n409, reg_p1_n408, reg_p1_n407,
         reg_p1_n406, reg_p1_n405, reg_p1_n404, reg_p1_n403, reg_p1_n402,
         reg_p1_n401, reg_p1_n400, reg_p1_n399, reg_p1_n398, reg_p1_n397,
         reg_p1_n396, reg_p1_n395, reg_p1_n394, reg_p1_n265, reg_p1_n264,
         reg_p1_n263, reg_p1_n262, reg_p1_n261, reg_p1_n260, reg_p1_n259,
         reg_p1_n258, reg_p1_n257, reg_p1_n256, reg_p1_n255, reg_p1_n254,
         reg_p1_n253, reg_p1_n252, reg_p1_n251, reg_p1_n250, reg_p1_n249,
         reg_p1_n248, reg_p1_n247, reg_p1_n246, reg_p1_n245, reg_p1_n244,
         reg_p1_n243, reg_p1_n242, reg_p1_n241, reg_p1_n240, reg_p1_n239,
         reg_p1_n238, reg_p1_n237, reg_p1_n236, reg_p1_n235, reg_p1_n234,
         reg_p1_n233, reg_p1_n232, reg_p1_n231, reg_p1_n230, reg_p1_n229,
         reg_p1_n228, reg_p1_n227, reg_p1_n226, reg_p1_n225, reg_p1_n224,
         reg_p1_n223, reg_p1_n222, reg_p1_n221, reg_p1_n220, reg_p1_n219,
         reg_p1_n218, reg_p1_n217, reg_p1_n216, reg_p1_n215, reg_p1_n214,
         reg_p1_n213, reg_p1_n212, reg_p1_n211, reg_p1_n210, reg_p1_n209,
         reg_p1_n208, reg_p1_n207, reg_p1_n206, reg_p1_n205, reg_p1_n204,
         reg_p1_n203, reg_p1_n202, mux_x_n138, mux_x_n137, mux_x_n136,
         mux_x_n135, mux_y_n267, mux_y_n266, mux_y_n265, mux_y_n264,
         mux_y_n263, cntrl_inst_n168, cntrl_inst_n167, cntrl_inst_n166,
         cntrl_inst_n165, cntrl_inst_n164, cntrl_inst_n163, cntrl_inst_n162,
         cntrl_inst_n161, cntrl_inst_n160, cntrl_inst_n159, cntrl_inst_n158,
         cntrl_inst_n157, cntrl_inst_n156, cntrl_inst_n155, cntrl_inst_n154,
         cntrl_inst_n153, cntrl_inst_n152, cntrl_inst_n151, cntrl_inst_n150,
         cntrl_inst_n149, cntrl_inst_n148, cntrl_inst_n147, cntrl_inst_n146,
         cntrl_inst_n145, cntrl_inst_n144, cntrl_inst_n143, cntrl_inst_n142,
         cntrl_inst_n141, cntrl_inst_n140, cntrl_inst_n139, cntrl_inst_n138,
         cntrl_inst_n137, cntrl_inst_n136, cntrl_inst_n135, cntrl_inst_n134,
         cntrl_inst_n133, cntrl_inst_n132, cntrl_inst_n131, cntrl_inst_n130,
         cntrl_inst_n129, cntrl_inst_n128, cntrl_inst_n127, cntrl_inst_n126,
         cntrl_inst_n125, cntrl_inst_n124, cntrl_inst_n123, cntrl_inst_n122,
         cntrl_inst_n121, cntrl_inst_n120, cntrl_inst_n119, cntrl_inst_n118,
         cntrl_inst_n117, cntrl_inst_n116, cntrl_inst_n115, cntrl_inst_n114,
         cntrl_inst_n113, cntrl_inst_n112, cntrl_inst_n111, cntrl_inst_n110,
         cntrl_inst_n109, cntrl_inst_n108, cntrl_inst_n107, cntrl_inst_n106,
         cntrl_inst_n105, cntrl_inst_n104, cntrl_inst_n103, cntrl_inst_n102,
         cntrl_inst_n101, cntrl_inst_n100, cntrl_inst_n99, cntrl_inst_n98,
         cntrl_inst_n97, cntrl_inst_n96, cntrl_inst_n95, cntrl_inst_n94,
         cntrl_inst_n93, cntrl_inst_n92, cntrl_inst_n91, cntrl_inst_n90,
         cntrl_inst_n89, cntrl_inst_n88, cntrl_inst_n87, cntrl_inst_n86,
         cntrl_inst_n85, cntrl_inst_n84, cntrl_inst_n83, cntrl_inst_n82,
         cntrl_inst_n81, cntrl_inst_n80, cntrl_inst_n79, cntrl_inst_n78,
         cntrl_inst_n77, cntrl_inst_n76, cntrl_inst_n75, cntrl_inst_n74,
         cntrl_inst_n73, cntrl_inst_n72, cntrl_inst_n71, cntrl_inst_n70,
         cntrl_inst_n69, cntrl_inst_n68, cntrl_inst_n67, cntrl_inst_n66,
         cntrl_inst_n65, cntrl_inst_n64, cntrl_inst_n63, cntrl_inst_n62,
         cntrl_inst_n61, cntrl_inst_n60, cntrl_inst_n59, cntrl_inst_n58,
         cntrl_inst_n57, cntrl_inst_n56, cntrl_inst_n55, cntrl_inst_n54,
         cntrl_inst_n53, cntrl_inst_n52, cntrl_inst_n51, cntrl_inst_n50,
         cntrl_inst_n49, cntrl_inst_n48, cntrl_inst_n47, cntrl_inst_n46,
         cntrl_inst_n45, cntrl_inst_n44, cntrl_inst_n43, cntrl_inst_n42,
         cntrl_inst_n41, cntrl_inst_n39, cntrl_inst_n38, cntrl_inst_n37,
         cntrl_inst_n35, cntrl_inst_n34, cntrl_inst_n33, cntrl_inst_n32,
         cntrl_inst_n31, cntrl_inst_n30, cntrl_inst_n29, cntrl_inst_n28,
         cntrl_inst_n27, cntrl_inst_n26, cntrl_inst_n25, cntrl_inst_n24,
         cntrl_inst_n23, cntrl_inst_n22, cntrl_inst_n21, cntrl_inst_n20,
         cntrl_inst_n19, cntrl_inst_n18, cntrl_inst_n17, cntrl_inst_n16,
         cntrl_inst_n15, cntrl_inst_n14, cntrl_inst_n13, cntrl_inst_n12,
         cntrl_inst_n11, cntrl_inst_n10, cntrl_inst_n9, cntrl_inst_n8,
         cntrl_inst_n7, cntrl_inst_n6, cntrl_inst_n5, cntrl_inst_n4,
         cntrl_inst_n3, cntrl_inst_n210, cntrl_inst_n209, cntrl_inst_n208,
         cntrl_inst_n207, cntrl_inst_n40, cntrl_inst_n36,
         cntrl_inst_counter_0_, prince_inst_n34, prince_inst_n33,
         prince_inst_n32, prince_inst_n31, prince_inst_n30, prince_inst_n29,
         prince_inst_n28, prince_inst_n27, prince_inst_n26, prince_inst_n25,
         prince_inst_n24, prince_inst_n23, prince_inst_n22, prince_inst_n21,
         prince_inst_n20, prince_inst_n19, prince_inst_sbox_inst0_n13,
         prince_inst_sbox_inst0_n12, prince_inst_sbox_inst0_n11,
         prince_inst_sbox_inst0_n10, prince_inst_sbox_inst0_n9,
         prince_inst_sbox_inst0_n8, prince_inst_sbox_inst0_n7,
         prince_inst_sbox_inst0_xxxy_inst_n20,
         prince_inst_sbox_inst0_xxxy_inst_n19,
         prince_inst_sbox_inst0_xxxy_inst_n18,
         prince_inst_sbox_inst0_xxxy_inst_n17,
         prince_inst_sbox_inst0_xxxy_inst_n16,
         prince_inst_sbox_inst0_xxxy_inst_n15,
         prince_inst_sbox_inst0_xxxy_inst_n14,
         prince_inst_sbox_inst0_xxxy_inst_n13,
         prince_inst_sbox_inst0_xxxy_inst_n12,
         prince_inst_sbox_inst0_xxxy_inst_n11,
         prince_inst_sbox_inst0_xxxy_inst_n10,
         prince_inst_sbox_inst0_xxxy_inst_n9,
         prince_inst_sbox_inst0_xxxy_inst_n8,
         prince_inst_sbox_inst0_xxxy_inst_n7,
         prince_inst_sbox_inst0_xxxy_inst_n6,
         prince_inst_sbox_inst0_xxxy_inst_n5,
         prince_inst_sbox_inst0_xxxy_inst_n4,
         prince_inst_sbox_inst0_xxxy_inst_n3,
         prince_inst_sbox_inst0_xxxy_inst_n2,
         prince_inst_sbox_inst0_xxxy_inst_n1,
         prince_inst_sbox_inst0_xxyx_inst_n18,
         prince_inst_sbox_inst0_xxyx_inst_n17,
         prince_inst_sbox_inst0_xxyx_inst_n16,
         prince_inst_sbox_inst0_xxyx_inst_n15,
         prince_inst_sbox_inst0_xxyx_inst_n14,
         prince_inst_sbox_inst0_xxyx_inst_n13,
         prince_inst_sbox_inst0_xxyx_inst_n12,
         prince_inst_sbox_inst0_xxyx_inst_n11,
         prince_inst_sbox_inst0_xxyx_inst_n10,
         prince_inst_sbox_inst0_xxyx_inst_n9,
         prince_inst_sbox_inst0_xxyx_inst_n8,
         prince_inst_sbox_inst0_xxyx_inst_n7,
         prince_inst_sbox_inst0_xxyx_inst_n6,
         prince_inst_sbox_inst0_xxyx_inst_n5,
         prince_inst_sbox_inst0_xxyx_inst_n4,
         prince_inst_sbox_inst0_xxyx_inst_n3,
         prince_inst_sbox_inst0_xxyx_inst_n2,
         prince_inst_sbox_inst0_xxyx_inst_n1,
         prince_inst_sbox_inst0_xyxx_inst_n22,
         prince_inst_sbox_inst0_xyxx_inst_n21,
         prince_inst_sbox_inst0_xyxx_inst_n20,
         prince_inst_sbox_inst0_xyxx_inst_n19,
         prince_inst_sbox_inst0_xyxx_inst_n18,
         prince_inst_sbox_inst0_xyxx_inst_n17,
         prince_inst_sbox_inst0_xyxx_inst_n16,
         prince_inst_sbox_inst0_xyxx_inst_n15,
         prince_inst_sbox_inst0_xyxx_inst_n14,
         prince_inst_sbox_inst0_xyxx_inst_n13,
         prince_inst_sbox_inst0_xyxx_inst_n12,
         prince_inst_sbox_inst0_xyxx_inst_n11,
         prince_inst_sbox_inst0_xyxx_inst_n10,
         prince_inst_sbox_inst0_xyxx_inst_n9,
         prince_inst_sbox_inst0_xyxx_inst_n8,
         prince_inst_sbox_inst0_xyxx_inst_n7,
         prince_inst_sbox_inst0_xyxx_inst_n6,
         prince_inst_sbox_inst0_xyxx_inst_n5,
         prince_inst_sbox_inst0_xyxx_inst_n4,
         prince_inst_sbox_inst0_xyxx_inst_n3,
         prince_inst_sbox_inst0_xyxx_inst_n2,
         prince_inst_sbox_inst0_xyxx_inst_n1,
         prince_inst_sbox_inst0_xyyy_inst_n31,
         prince_inst_sbox_inst0_xyyy_inst_n30,
         prince_inst_sbox_inst0_xyyy_inst_n29,
         prince_inst_sbox_inst0_xyyy_inst_n28,
         prince_inst_sbox_inst0_xyyy_inst_n27,
         prince_inst_sbox_inst0_xyyy_inst_n26,
         prince_inst_sbox_inst0_xyyy_inst_n25,
         prince_inst_sbox_inst0_xyyy_inst_n24,
         prince_inst_sbox_inst0_xyyy_inst_n23,
         prince_inst_sbox_inst0_xyyy_inst_n22,
         prince_inst_sbox_inst0_xyyy_inst_n21,
         prince_inst_sbox_inst0_xyyy_inst_n20,
         prince_inst_sbox_inst0_xyyy_inst_n19,
         prince_inst_sbox_inst0_xyyy_inst_n18,
         prince_inst_sbox_inst0_xyyy_inst_n17,
         prince_inst_sbox_inst0_xyyy_inst_n16,
         prince_inst_sbox_inst0_xyyy_inst_n15,
         prince_inst_sbox_inst0_xyyy_inst_n14,
         prince_inst_sbox_inst0_xyyy_inst_n13,
         prince_inst_sbox_inst0_xyyy_inst_n12,
         prince_inst_sbox_inst0_yxxx_inst_n21,
         prince_inst_sbox_inst0_yxxx_inst_n20,
         prince_inst_sbox_inst0_yxxx_inst_n19,
         prince_inst_sbox_inst0_yxxx_inst_n18,
         prince_inst_sbox_inst0_yxxx_inst_n17,
         prince_inst_sbox_inst0_yxxx_inst_n16,
         prince_inst_sbox_inst0_yxxx_inst_n15,
         prince_inst_sbox_inst0_yxxx_inst_n14,
         prince_inst_sbox_inst0_yxxx_inst_n13,
         prince_inst_sbox_inst0_yxxx_inst_n12,
         prince_inst_sbox_inst0_yxxx_inst_n11,
         prince_inst_sbox_inst0_yxxx_inst_n10,
         prince_inst_sbox_inst0_yxxx_inst_n9,
         prince_inst_sbox_inst0_yxxx_inst_n8,
         prince_inst_sbox_inst0_yxxx_inst_n7,
         prince_inst_sbox_inst0_yxxx_inst_n6,
         prince_inst_sbox_inst0_yxxx_inst_n5,
         prince_inst_sbox_inst0_yxxx_inst_n4,
         prince_inst_sbox_inst0_yxxx_inst_n3,
         prince_inst_sbox_inst0_yxxx_inst_n2,
         prince_inst_sbox_inst0_yxyy_inst_n19,
         prince_inst_sbox_inst0_yxyy_inst_n18,
         prince_inst_sbox_inst0_yxyy_inst_n17,
         prince_inst_sbox_inst0_yxyy_inst_n16,
         prince_inst_sbox_inst0_yxyy_inst_n15,
         prince_inst_sbox_inst0_yxyy_inst_n14,
         prince_inst_sbox_inst0_yxyy_inst_n13,
         prince_inst_sbox_inst0_yxyy_inst_n12,
         prince_inst_sbox_inst0_yxyy_inst_n11,
         prince_inst_sbox_inst0_yxyy_inst_n10,
         prince_inst_sbox_inst0_yxyy_inst_n9,
         prince_inst_sbox_inst0_yxyy_inst_n8,
         prince_inst_sbox_inst0_yxyy_inst_n7,
         prince_inst_sbox_inst0_yxyy_inst_n6,
         prince_inst_sbox_inst0_yxyy_inst_n5,
         prince_inst_sbox_inst0_yxyy_inst_n4,
         prince_inst_sbox_inst0_yxyy_inst_n3,
         prince_inst_sbox_inst0_yxyy_inst_n2,
         prince_inst_sbox_inst0_yxyy_inst_n1,
         prince_inst_sbox_inst0_yyxy_inst_n16,
         prince_inst_sbox_inst0_yyxy_inst_n15,
         prince_inst_sbox_inst0_yyxy_inst_n14,
         prince_inst_sbox_inst0_yyxy_inst_n13,
         prince_inst_sbox_inst0_yyxy_inst_n12,
         prince_inst_sbox_inst0_yyxy_inst_n11,
         prince_inst_sbox_inst0_yyxy_inst_n10,
         prince_inst_sbox_inst0_yyxy_inst_n9,
         prince_inst_sbox_inst0_yyxy_inst_n8,
         prince_inst_sbox_inst0_yyxy_inst_n7,
         prince_inst_sbox_inst0_yyxy_inst_n6,
         prince_inst_sbox_inst0_yyxy_inst_n5,
         prince_inst_sbox_inst0_yyxy_inst_n4,
         prince_inst_sbox_inst0_yyxy_inst_n3,
         prince_inst_sbox_inst0_yyxy_inst_n2,
         prince_inst_sbox_inst0_yyxy_inst_n1,
         prince_inst_sbox_inst0_yyyx_inst_n38,
         prince_inst_sbox_inst0_yyyx_inst_n37,
         prince_inst_sbox_inst0_yyyx_inst_n36,
         prince_inst_sbox_inst0_yyyx_inst_n35,
         prince_inst_sbox_inst0_yyyx_inst_n34,
         prince_inst_sbox_inst0_yyyx_inst_n33,
         prince_inst_sbox_inst0_yyyx_inst_n32,
         prince_inst_sbox_inst0_yyyx_inst_n31,
         prince_inst_sbox_inst0_yyyx_inst_n30,
         prince_inst_sbox_inst0_yyyx_inst_n29,
         prince_inst_sbox_inst0_yyyx_inst_n28,
         prince_inst_sbox_inst0_yyyx_inst_n27,
         prince_inst_sbox_inst0_yyyx_inst_n26,
         prince_inst_sbox_inst0_yyyx_inst_n25,
         prince_inst_sbox_inst0_yyyx_inst_n24,
         prince_inst_sbox_inst0_yyyx_inst_n23,
         prince_inst_sbox_inst0_yyyx_inst_n22,
         prince_inst_sbox_inst0_c_inst0_msk0_xr,
         prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n4,
         prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n3,
         prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n2,
         prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n5,
         prince_inst_sbox_inst0_c_inst0_msk1_xr,
         prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst0_msk2_xr,
         prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst0_msk3_xr,
         prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst0_msk4_xr,
         prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst0_msk5_xr,
         prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst0_msk6_xr,
         prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst0_msk7_xr,
         prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst0_ax_n2,
         prince_inst_sbox_inst0_c_inst0_ax_n1,
         prince_inst_sbox_inst0_c_inst0_ay_n6,
         prince_inst_sbox_inst0_c_inst0_ay_n5,
         prince_inst_sbox_inst0_c_inst1_msk0_xr,
         prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_msk1_xr,
         prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_msk2_xr,
         prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_msk3_xr,
         prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_msk4_xr,
         prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_msk5_xr,
         prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_msk6_xr,
         prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_msk7_xr,
         prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst1_ax_n6,
         prince_inst_sbox_inst0_c_inst1_ax_n5,
         prince_inst_sbox_inst0_c_inst1_ay_n6,
         prince_inst_sbox_inst0_c_inst1_ay_n5,
         prince_inst_sbox_inst0_c_inst2_msk0_xr,
         prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_msk1_xr,
         prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_msk2_xr,
         prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_msk3_xr,
         prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_msk4_xr,
         prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_msk5_xr,
         prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_msk6_xr,
         prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_msk7_xr,
         prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst2_ax_n6,
         prince_inst_sbox_inst0_c_inst2_ax_n5,
         prince_inst_sbox_inst0_c_inst2_ay_n6,
         prince_inst_sbox_inst0_c_inst2_ay_n5,
         prince_inst_sbox_inst0_c_inst3_msk0_xr,
         prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_msk1_xr,
         prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_msk2_xr,
         prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_msk3_xr,
         prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_msk4_xr,
         prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_msk5_xr,
         prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_msk6_xr,
         prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_msk7_xr,
         prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst0_c_inst3_ax_n6,
         prince_inst_sbox_inst0_c_inst3_ax_n5,
         prince_inst_sbox_inst0_c_inst3_ay_n6,
         prince_inst_sbox_inst0_c_inst3_ay_n5, prince_inst_sbox_inst1_n13,
         prince_inst_sbox_inst1_n12, prince_inst_sbox_inst1_n11,
         prince_inst_sbox_inst1_n10, prince_inst_sbox_inst1_n9,
         prince_inst_sbox_inst1_n8, prince_inst_sbox_inst1_n7,
         prince_inst_sbox_inst1_xxxy_inst_n70,
         prince_inst_sbox_inst1_xxxy_inst_n69,
         prince_inst_sbox_inst1_xxxy_inst_n68,
         prince_inst_sbox_inst1_xxxy_inst_n67,
         prince_inst_sbox_inst1_xxxy_inst_n66,
         prince_inst_sbox_inst1_xxxy_inst_n65,
         prince_inst_sbox_inst1_xxxy_inst_n64,
         prince_inst_sbox_inst1_xxxy_inst_n63,
         prince_inst_sbox_inst1_xxxy_inst_n62,
         prince_inst_sbox_inst1_xxxy_inst_n61,
         prince_inst_sbox_inst1_xxxy_inst_n60,
         prince_inst_sbox_inst1_xxxy_inst_n59,
         prince_inst_sbox_inst1_xxxy_inst_n58,
         prince_inst_sbox_inst1_xxxy_inst_n57,
         prince_inst_sbox_inst1_xxxy_inst_n56,
         prince_inst_sbox_inst1_xxxy_inst_n55,
         prince_inst_sbox_inst1_xxxy_inst_n54,
         prince_inst_sbox_inst1_xxxy_inst_n53,
         prince_inst_sbox_inst1_xxxy_inst_n52,
         prince_inst_sbox_inst1_xxxy_inst_n51,
         prince_inst_sbox_inst1_xxyx_inst_n55,
         prince_inst_sbox_inst1_xxyx_inst_n54,
         prince_inst_sbox_inst1_xxyx_inst_n53,
         prince_inst_sbox_inst1_xxyx_inst_n52,
         prince_inst_sbox_inst1_xxyx_inst_n51,
         prince_inst_sbox_inst1_xxyx_inst_n50,
         prince_inst_sbox_inst1_xxyx_inst_n49,
         prince_inst_sbox_inst1_xxyx_inst_n48,
         prince_inst_sbox_inst1_xxyx_inst_n47,
         prince_inst_sbox_inst1_xxyx_inst_n46,
         prince_inst_sbox_inst1_xxyx_inst_n45,
         prince_inst_sbox_inst1_xxyx_inst_n44,
         prince_inst_sbox_inst1_xxyx_inst_n43,
         prince_inst_sbox_inst1_xxyx_inst_n42,
         prince_inst_sbox_inst1_xxyx_inst_n41,
         prince_inst_sbox_inst1_xxyx_inst_n40,
         prince_inst_sbox_inst1_xxyx_inst_n39,
         prince_inst_sbox_inst1_xxyx_inst_n38,
         prince_inst_sbox_inst1_xyxx_inst_n74,
         prince_inst_sbox_inst1_xyxx_inst_n73,
         prince_inst_sbox_inst1_xyxx_inst_n72,
         prince_inst_sbox_inst1_xyxx_inst_n71,
         prince_inst_sbox_inst1_xyxx_inst_n70,
         prince_inst_sbox_inst1_xyxx_inst_n69,
         prince_inst_sbox_inst1_xyxx_inst_n68,
         prince_inst_sbox_inst1_xyxx_inst_n67,
         prince_inst_sbox_inst1_xyxx_inst_n66,
         prince_inst_sbox_inst1_xyxx_inst_n65,
         prince_inst_sbox_inst1_xyxx_inst_n64,
         prince_inst_sbox_inst1_xyxx_inst_n63,
         prince_inst_sbox_inst1_xyxx_inst_n62,
         prince_inst_sbox_inst1_xyxx_inst_n61,
         prince_inst_sbox_inst1_xyxx_inst_n60,
         prince_inst_sbox_inst1_xyxx_inst_n59,
         prince_inst_sbox_inst1_xyxx_inst_n58,
         prince_inst_sbox_inst1_xyxx_inst_n57,
         prince_inst_sbox_inst1_xyxx_inst_n56,
         prince_inst_sbox_inst1_xyxx_inst_n55,
         prince_inst_sbox_inst1_xyxx_inst_n54,
         prince_inst_sbox_inst1_xyxx_inst_n53,
         prince_inst_sbox_inst1_xyyy_inst_n61,
         prince_inst_sbox_inst1_xyyy_inst_n60,
         prince_inst_sbox_inst1_xyyy_inst_n59,
         prince_inst_sbox_inst1_xyyy_inst_n58,
         prince_inst_sbox_inst1_xyyy_inst_n57,
         prince_inst_sbox_inst1_xyyy_inst_n56,
         prince_inst_sbox_inst1_xyyy_inst_n55,
         prince_inst_sbox_inst1_xyyy_inst_n54,
         prince_inst_sbox_inst1_xyyy_inst_n53,
         prince_inst_sbox_inst1_xyyy_inst_n52,
         prince_inst_sbox_inst1_xyyy_inst_n51,
         prince_inst_sbox_inst1_xyyy_inst_n50,
         prince_inst_sbox_inst1_xyyy_inst_n49,
         prince_inst_sbox_inst1_xyyy_inst_n48,
         prince_inst_sbox_inst1_xyyy_inst_n47,
         prince_inst_sbox_inst1_xyyy_inst_n46,
         prince_inst_sbox_inst1_xyyy_inst_n45,
         prince_inst_sbox_inst1_xyyy_inst_n44,
         prince_inst_sbox_inst1_xyyy_inst_n43,
         prince_inst_sbox_inst1_xyyy_inst_n42,
         prince_inst_sbox_inst1_yxxx_inst_n64,
         prince_inst_sbox_inst1_yxxx_inst_n63,
         prince_inst_sbox_inst1_yxxx_inst_n62,
         prince_inst_sbox_inst1_yxxx_inst_n61,
         prince_inst_sbox_inst1_yxxx_inst_n60,
         prince_inst_sbox_inst1_yxxx_inst_n59,
         prince_inst_sbox_inst1_yxxx_inst_n58,
         prince_inst_sbox_inst1_yxxx_inst_n57,
         prince_inst_sbox_inst1_yxxx_inst_n56,
         prince_inst_sbox_inst1_yxxx_inst_n55,
         prince_inst_sbox_inst1_yxxx_inst_n54,
         prince_inst_sbox_inst1_yxxx_inst_n53,
         prince_inst_sbox_inst1_yxxx_inst_n52,
         prince_inst_sbox_inst1_yxxx_inst_n51,
         prince_inst_sbox_inst1_yxxx_inst_n50,
         prince_inst_sbox_inst1_yxxx_inst_n49,
         prince_inst_sbox_inst1_yxxx_inst_n48,
         prince_inst_sbox_inst1_yxxx_inst_n47,
         prince_inst_sbox_inst1_yxxx_inst_n46,
         prince_inst_sbox_inst1_yxxx_inst_n45,
         prince_inst_sbox_inst1_yxyy_inst_n67,
         prince_inst_sbox_inst1_yxyy_inst_n66,
         prince_inst_sbox_inst1_yxyy_inst_n65,
         prince_inst_sbox_inst1_yxyy_inst_n64,
         prince_inst_sbox_inst1_yxyy_inst_n63,
         prince_inst_sbox_inst1_yxyy_inst_n62,
         prince_inst_sbox_inst1_yxyy_inst_n61,
         prince_inst_sbox_inst1_yxyy_inst_n60,
         prince_inst_sbox_inst1_yxyy_inst_n59,
         prince_inst_sbox_inst1_yxyy_inst_n58,
         prince_inst_sbox_inst1_yxyy_inst_n57,
         prince_inst_sbox_inst1_yxyy_inst_n56,
         prince_inst_sbox_inst1_yxyy_inst_n55,
         prince_inst_sbox_inst1_yxyy_inst_n54,
         prince_inst_sbox_inst1_yxyy_inst_n53,
         prince_inst_sbox_inst1_yxyy_inst_n52,
         prince_inst_sbox_inst1_yxyy_inst_n51,
         prince_inst_sbox_inst1_yxyy_inst_n50,
         prince_inst_sbox_inst1_yxyy_inst_n49,
         prince_inst_sbox_inst1_yyxy_inst_n75,
         prince_inst_sbox_inst1_yyxy_inst_n74,
         prince_inst_sbox_inst1_yyxy_inst_n73,
         prince_inst_sbox_inst1_yyxy_inst_n72,
         prince_inst_sbox_inst1_yyxy_inst_n71,
         prince_inst_sbox_inst1_yyxy_inst_n70,
         prince_inst_sbox_inst1_yyxy_inst_n69,
         prince_inst_sbox_inst1_yyxy_inst_n68,
         prince_inst_sbox_inst1_yyxy_inst_n67,
         prince_inst_sbox_inst1_yyxy_inst_n66,
         prince_inst_sbox_inst1_yyxy_inst_n65,
         prince_inst_sbox_inst1_yyxy_inst_n64,
         prince_inst_sbox_inst1_yyxy_inst_n63,
         prince_inst_sbox_inst1_yyxy_inst_n62,
         prince_inst_sbox_inst1_yyxy_inst_n61,
         prince_inst_sbox_inst1_yyxy_inst_n60,
         prince_inst_sbox_inst1_yyxy_inst_n59,
         prince_inst_sbox_inst1_yyxy_inst_n58,
         prince_inst_sbox_inst1_yyxy_inst_n57,
         prince_inst_sbox_inst1_yyxy_inst_n56,
         prince_inst_sbox_inst1_yyxy_inst_n55,
         prince_inst_sbox_inst1_yyxy_inst_n54,
         prince_inst_sbox_inst1_yyxy_inst_n53,
         prince_inst_sbox_inst1_yyyx_inst_n58,
         prince_inst_sbox_inst1_yyyx_inst_n57,
         prince_inst_sbox_inst1_yyyx_inst_n56,
         prince_inst_sbox_inst1_yyyx_inst_n55,
         prince_inst_sbox_inst1_yyyx_inst_n54,
         prince_inst_sbox_inst1_yyyx_inst_n53,
         prince_inst_sbox_inst1_yyyx_inst_n52,
         prince_inst_sbox_inst1_yyyx_inst_n51,
         prince_inst_sbox_inst1_yyyx_inst_n50,
         prince_inst_sbox_inst1_yyyx_inst_n49,
         prince_inst_sbox_inst1_yyyx_inst_n48,
         prince_inst_sbox_inst1_yyyx_inst_n47,
         prince_inst_sbox_inst1_yyyx_inst_n46,
         prince_inst_sbox_inst1_yyyx_inst_n45,
         prince_inst_sbox_inst1_yyyx_inst_n44,
         prince_inst_sbox_inst1_yyyx_inst_n43,
         prince_inst_sbox_inst1_yyyx_inst_n42,
         prince_inst_sbox_inst1_c_inst0_msk0_xr,
         prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_msk1_xr,
         prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_msk2_xr,
         prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_msk3_xr,
         prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_msk4_xr,
         prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_msk5_xr,
         prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_msk6_xr,
         prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_msk7_xr,
         prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst0_ax_n6,
         prince_inst_sbox_inst1_c_inst0_ax_n5,
         prince_inst_sbox_inst1_c_inst0_ay_n6,
         prince_inst_sbox_inst1_c_inst0_ay_n5,
         prince_inst_sbox_inst1_c_inst1_msk0_xr,
         prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_msk1_xr,
         prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_msk2_xr,
         prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_msk3_xr,
         prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_msk4_xr,
         prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_msk5_xr,
         prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_msk6_xr,
         prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_msk7_xr,
         prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst1_ax_n6,
         prince_inst_sbox_inst1_c_inst1_ax_n5,
         prince_inst_sbox_inst1_c_inst1_ay_n6,
         prince_inst_sbox_inst1_c_inst1_ay_n5,
         prince_inst_sbox_inst1_c_inst2_msk0_xr,
         prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_msk1_xr,
         prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_msk2_xr,
         prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_msk3_xr,
         prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_msk4_xr,
         prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_msk5_xr,
         prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_msk6_xr,
         prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_msk7_xr,
         prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst2_ax_n6,
         prince_inst_sbox_inst1_c_inst2_ax_n5,
         prince_inst_sbox_inst1_c_inst2_ay_n6,
         prince_inst_sbox_inst1_c_inst2_ay_n5,
         prince_inst_sbox_inst1_c_inst3_msk0_xr,
         prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_msk1_xr,
         prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_msk2_xr,
         prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_msk3_xr,
         prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_msk4_xr,
         prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_msk5_xr,
         prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_msk6_xr,
         prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_msk7_xr,
         prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst1_c_inst3_ax_n6,
         prince_inst_sbox_inst1_c_inst3_ax_n5,
         prince_inst_sbox_inst1_c_inst3_ay_n6,
         prince_inst_sbox_inst1_c_inst3_ay_n5, prince_inst_sbox_inst2_n12,
         prince_inst_sbox_inst2_n11, prince_inst_sbox_inst2_n10,
         prince_inst_sbox_inst2_n9, prince_inst_sbox_inst2_n8,
         prince_inst_sbox_inst2_n7, prince_inst_sbox_inst2_n6,
         prince_inst_sbox_inst2_xxxy_inst_n70,
         prince_inst_sbox_inst2_xxxy_inst_n69,
         prince_inst_sbox_inst2_xxxy_inst_n68,
         prince_inst_sbox_inst2_xxxy_inst_n67,
         prince_inst_sbox_inst2_xxxy_inst_n66,
         prince_inst_sbox_inst2_xxxy_inst_n65,
         prince_inst_sbox_inst2_xxxy_inst_n64,
         prince_inst_sbox_inst2_xxxy_inst_n63,
         prince_inst_sbox_inst2_xxxy_inst_n62,
         prince_inst_sbox_inst2_xxxy_inst_n61,
         prince_inst_sbox_inst2_xxxy_inst_n60,
         prince_inst_sbox_inst2_xxxy_inst_n59,
         prince_inst_sbox_inst2_xxxy_inst_n58,
         prince_inst_sbox_inst2_xxxy_inst_n57,
         prince_inst_sbox_inst2_xxxy_inst_n56,
         prince_inst_sbox_inst2_xxxy_inst_n55,
         prince_inst_sbox_inst2_xxxy_inst_n54,
         prince_inst_sbox_inst2_xxxy_inst_n53,
         prince_inst_sbox_inst2_xxxy_inst_n52,
         prince_inst_sbox_inst2_xxxy_inst_n51,
         prince_inst_sbox_inst2_xxyx_inst_n55,
         prince_inst_sbox_inst2_xxyx_inst_n54,
         prince_inst_sbox_inst2_xxyx_inst_n53,
         prince_inst_sbox_inst2_xxyx_inst_n52,
         prince_inst_sbox_inst2_xxyx_inst_n51,
         prince_inst_sbox_inst2_xxyx_inst_n50,
         prince_inst_sbox_inst2_xxyx_inst_n49,
         prince_inst_sbox_inst2_xxyx_inst_n48,
         prince_inst_sbox_inst2_xxyx_inst_n47,
         prince_inst_sbox_inst2_xxyx_inst_n46,
         prince_inst_sbox_inst2_xxyx_inst_n45,
         prince_inst_sbox_inst2_xxyx_inst_n44,
         prince_inst_sbox_inst2_xxyx_inst_n43,
         prince_inst_sbox_inst2_xxyx_inst_n42,
         prince_inst_sbox_inst2_xxyx_inst_n41,
         prince_inst_sbox_inst2_xxyx_inst_n40,
         prince_inst_sbox_inst2_xxyx_inst_n39,
         prince_inst_sbox_inst2_xxyx_inst_n38,
         prince_inst_sbox_inst2_xyxx_inst_n74,
         prince_inst_sbox_inst2_xyxx_inst_n73,
         prince_inst_sbox_inst2_xyxx_inst_n72,
         prince_inst_sbox_inst2_xyxx_inst_n71,
         prince_inst_sbox_inst2_xyxx_inst_n70,
         prince_inst_sbox_inst2_xyxx_inst_n69,
         prince_inst_sbox_inst2_xyxx_inst_n68,
         prince_inst_sbox_inst2_xyxx_inst_n67,
         prince_inst_sbox_inst2_xyxx_inst_n66,
         prince_inst_sbox_inst2_xyxx_inst_n65,
         prince_inst_sbox_inst2_xyxx_inst_n64,
         prince_inst_sbox_inst2_xyxx_inst_n63,
         prince_inst_sbox_inst2_xyxx_inst_n62,
         prince_inst_sbox_inst2_xyxx_inst_n61,
         prince_inst_sbox_inst2_xyxx_inst_n60,
         prince_inst_sbox_inst2_xyxx_inst_n59,
         prince_inst_sbox_inst2_xyxx_inst_n58,
         prince_inst_sbox_inst2_xyxx_inst_n57,
         prince_inst_sbox_inst2_xyxx_inst_n56,
         prince_inst_sbox_inst2_xyxx_inst_n55,
         prince_inst_sbox_inst2_xyxx_inst_n54,
         prince_inst_sbox_inst2_xyxx_inst_n53,
         prince_inst_sbox_inst2_xyyy_inst_n61,
         prince_inst_sbox_inst2_xyyy_inst_n60,
         prince_inst_sbox_inst2_xyyy_inst_n59,
         prince_inst_sbox_inst2_xyyy_inst_n58,
         prince_inst_sbox_inst2_xyyy_inst_n57,
         prince_inst_sbox_inst2_xyyy_inst_n56,
         prince_inst_sbox_inst2_xyyy_inst_n55,
         prince_inst_sbox_inst2_xyyy_inst_n54,
         prince_inst_sbox_inst2_xyyy_inst_n53,
         prince_inst_sbox_inst2_xyyy_inst_n52,
         prince_inst_sbox_inst2_xyyy_inst_n51,
         prince_inst_sbox_inst2_xyyy_inst_n50,
         prince_inst_sbox_inst2_xyyy_inst_n49,
         prince_inst_sbox_inst2_xyyy_inst_n48,
         prince_inst_sbox_inst2_xyyy_inst_n47,
         prince_inst_sbox_inst2_xyyy_inst_n46,
         prince_inst_sbox_inst2_xyyy_inst_n45,
         prince_inst_sbox_inst2_xyyy_inst_n44,
         prince_inst_sbox_inst2_xyyy_inst_n43,
         prince_inst_sbox_inst2_xyyy_inst_n42,
         prince_inst_sbox_inst2_yxxx_inst_n64,
         prince_inst_sbox_inst2_yxxx_inst_n63,
         prince_inst_sbox_inst2_yxxx_inst_n62,
         prince_inst_sbox_inst2_yxxx_inst_n61,
         prince_inst_sbox_inst2_yxxx_inst_n60,
         prince_inst_sbox_inst2_yxxx_inst_n59,
         prince_inst_sbox_inst2_yxxx_inst_n58,
         prince_inst_sbox_inst2_yxxx_inst_n57,
         prince_inst_sbox_inst2_yxxx_inst_n56,
         prince_inst_sbox_inst2_yxxx_inst_n55,
         prince_inst_sbox_inst2_yxxx_inst_n54,
         prince_inst_sbox_inst2_yxxx_inst_n53,
         prince_inst_sbox_inst2_yxxx_inst_n52,
         prince_inst_sbox_inst2_yxxx_inst_n51,
         prince_inst_sbox_inst2_yxxx_inst_n50,
         prince_inst_sbox_inst2_yxxx_inst_n49,
         prince_inst_sbox_inst2_yxxx_inst_n48,
         prince_inst_sbox_inst2_yxxx_inst_n47,
         prince_inst_sbox_inst2_yxxx_inst_n46,
         prince_inst_sbox_inst2_yxxx_inst_n45,
         prince_inst_sbox_inst2_yxyy_inst_n67,
         prince_inst_sbox_inst2_yxyy_inst_n66,
         prince_inst_sbox_inst2_yxyy_inst_n65,
         prince_inst_sbox_inst2_yxyy_inst_n64,
         prince_inst_sbox_inst2_yxyy_inst_n63,
         prince_inst_sbox_inst2_yxyy_inst_n62,
         prince_inst_sbox_inst2_yxyy_inst_n61,
         prince_inst_sbox_inst2_yxyy_inst_n60,
         prince_inst_sbox_inst2_yxyy_inst_n59,
         prince_inst_sbox_inst2_yxyy_inst_n58,
         prince_inst_sbox_inst2_yxyy_inst_n57,
         prince_inst_sbox_inst2_yxyy_inst_n56,
         prince_inst_sbox_inst2_yxyy_inst_n55,
         prince_inst_sbox_inst2_yxyy_inst_n54,
         prince_inst_sbox_inst2_yxyy_inst_n53,
         prince_inst_sbox_inst2_yxyy_inst_n52,
         prince_inst_sbox_inst2_yxyy_inst_n51,
         prince_inst_sbox_inst2_yxyy_inst_n50,
         prince_inst_sbox_inst2_yxyy_inst_n49,
         prince_inst_sbox_inst2_yyxy_inst_n75,
         prince_inst_sbox_inst2_yyxy_inst_n74,
         prince_inst_sbox_inst2_yyxy_inst_n73,
         prince_inst_sbox_inst2_yyxy_inst_n72,
         prince_inst_sbox_inst2_yyxy_inst_n71,
         prince_inst_sbox_inst2_yyxy_inst_n70,
         prince_inst_sbox_inst2_yyxy_inst_n69,
         prince_inst_sbox_inst2_yyxy_inst_n68,
         prince_inst_sbox_inst2_yyxy_inst_n67,
         prince_inst_sbox_inst2_yyxy_inst_n66,
         prince_inst_sbox_inst2_yyxy_inst_n65,
         prince_inst_sbox_inst2_yyxy_inst_n64,
         prince_inst_sbox_inst2_yyxy_inst_n63,
         prince_inst_sbox_inst2_yyxy_inst_n62,
         prince_inst_sbox_inst2_yyxy_inst_n61,
         prince_inst_sbox_inst2_yyxy_inst_n60,
         prince_inst_sbox_inst2_yyxy_inst_n59,
         prince_inst_sbox_inst2_yyxy_inst_n58,
         prince_inst_sbox_inst2_yyxy_inst_n57,
         prince_inst_sbox_inst2_yyxy_inst_n56,
         prince_inst_sbox_inst2_yyxy_inst_n55,
         prince_inst_sbox_inst2_yyxy_inst_n54,
         prince_inst_sbox_inst2_yyxy_inst_n53,
         prince_inst_sbox_inst2_yyyx_inst_n58,
         prince_inst_sbox_inst2_yyyx_inst_n57,
         prince_inst_sbox_inst2_yyyx_inst_n56,
         prince_inst_sbox_inst2_yyyx_inst_n55,
         prince_inst_sbox_inst2_yyyx_inst_n54,
         prince_inst_sbox_inst2_yyyx_inst_n53,
         prince_inst_sbox_inst2_yyyx_inst_n52,
         prince_inst_sbox_inst2_yyyx_inst_n51,
         prince_inst_sbox_inst2_yyyx_inst_n50,
         prince_inst_sbox_inst2_yyyx_inst_n49,
         prince_inst_sbox_inst2_yyyx_inst_n48,
         prince_inst_sbox_inst2_yyyx_inst_n47,
         prince_inst_sbox_inst2_yyyx_inst_n46,
         prince_inst_sbox_inst2_yyyx_inst_n45,
         prince_inst_sbox_inst2_yyyx_inst_n44,
         prince_inst_sbox_inst2_yyyx_inst_n43,
         prince_inst_sbox_inst2_yyyx_inst_n42,
         prince_inst_sbox_inst2_c_inst0_msk0_xr,
         prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_msk1_xr,
         prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_msk2_xr,
         prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_msk3_xr,
         prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_msk4_xr,
         prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_msk5_xr,
         prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_msk6_xr,
         prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_msk7_xr,
         prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst0_ax_n6,
         prince_inst_sbox_inst2_c_inst0_ax_n5,
         prince_inst_sbox_inst2_c_inst0_ay_n6,
         prince_inst_sbox_inst2_c_inst0_ay_n5,
         prince_inst_sbox_inst2_c_inst1_msk0_xr,
         prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_msk1_xr,
         prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_msk2_xr,
         prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_msk3_xr,
         prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_msk4_xr,
         prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_msk5_xr,
         prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_msk6_xr,
         prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_msk7_xr,
         prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst1_ax_n6,
         prince_inst_sbox_inst2_c_inst1_ax_n5,
         prince_inst_sbox_inst2_c_inst1_ay_n6,
         prince_inst_sbox_inst2_c_inst1_ay_n5,
         prince_inst_sbox_inst2_c_inst2_msk0_xr,
         prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_msk1_xr,
         prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_msk2_xr,
         prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_msk3_xr,
         prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_msk4_xr,
         prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_msk5_xr,
         prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_msk6_xr,
         prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_msk7_xr,
         prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst2_ax_n6,
         prince_inst_sbox_inst2_c_inst2_ax_n5,
         prince_inst_sbox_inst2_c_inst2_ay_n6,
         prince_inst_sbox_inst2_c_inst2_ay_n5,
         prince_inst_sbox_inst2_c_inst3_msk0_xr,
         prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_msk1_xr,
         prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_msk2_xr,
         prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_msk3_xr,
         prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_msk4_xr,
         prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_msk5_xr,
         prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_msk6_xr,
         prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_msk7_xr,
         prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst2_c_inst3_ax_n6,
         prince_inst_sbox_inst2_c_inst3_ax_n5,
         prince_inst_sbox_inst2_c_inst3_ay_n6,
         prince_inst_sbox_inst2_c_inst3_ay_n5, prince_inst_sbox_inst3_n12,
         prince_inst_sbox_inst3_n11, prince_inst_sbox_inst3_n10,
         prince_inst_sbox_inst3_n9, prince_inst_sbox_inst3_n8,
         prince_inst_sbox_inst3_n7, prince_inst_sbox_inst3_n6,
         prince_inst_sbox_inst3_xxxy_inst_n70,
         prince_inst_sbox_inst3_xxxy_inst_n69,
         prince_inst_sbox_inst3_xxxy_inst_n68,
         prince_inst_sbox_inst3_xxxy_inst_n67,
         prince_inst_sbox_inst3_xxxy_inst_n66,
         prince_inst_sbox_inst3_xxxy_inst_n65,
         prince_inst_sbox_inst3_xxxy_inst_n64,
         prince_inst_sbox_inst3_xxxy_inst_n63,
         prince_inst_sbox_inst3_xxxy_inst_n62,
         prince_inst_sbox_inst3_xxxy_inst_n61,
         prince_inst_sbox_inst3_xxxy_inst_n60,
         prince_inst_sbox_inst3_xxxy_inst_n59,
         prince_inst_sbox_inst3_xxxy_inst_n58,
         prince_inst_sbox_inst3_xxxy_inst_n57,
         prince_inst_sbox_inst3_xxxy_inst_n56,
         prince_inst_sbox_inst3_xxxy_inst_n55,
         prince_inst_sbox_inst3_xxxy_inst_n54,
         prince_inst_sbox_inst3_xxxy_inst_n53,
         prince_inst_sbox_inst3_xxxy_inst_n52,
         prince_inst_sbox_inst3_xxxy_inst_n51,
         prince_inst_sbox_inst3_xxyx_inst_n55,
         prince_inst_sbox_inst3_xxyx_inst_n54,
         prince_inst_sbox_inst3_xxyx_inst_n53,
         prince_inst_sbox_inst3_xxyx_inst_n52,
         prince_inst_sbox_inst3_xxyx_inst_n51,
         prince_inst_sbox_inst3_xxyx_inst_n50,
         prince_inst_sbox_inst3_xxyx_inst_n49,
         prince_inst_sbox_inst3_xxyx_inst_n48,
         prince_inst_sbox_inst3_xxyx_inst_n47,
         prince_inst_sbox_inst3_xxyx_inst_n46,
         prince_inst_sbox_inst3_xxyx_inst_n45,
         prince_inst_sbox_inst3_xxyx_inst_n44,
         prince_inst_sbox_inst3_xxyx_inst_n43,
         prince_inst_sbox_inst3_xxyx_inst_n42,
         prince_inst_sbox_inst3_xxyx_inst_n41,
         prince_inst_sbox_inst3_xxyx_inst_n40,
         prince_inst_sbox_inst3_xxyx_inst_n39,
         prince_inst_sbox_inst3_xxyx_inst_n38,
         prince_inst_sbox_inst3_xyxx_inst_n74,
         prince_inst_sbox_inst3_xyxx_inst_n73,
         prince_inst_sbox_inst3_xyxx_inst_n72,
         prince_inst_sbox_inst3_xyxx_inst_n71,
         prince_inst_sbox_inst3_xyxx_inst_n70,
         prince_inst_sbox_inst3_xyxx_inst_n69,
         prince_inst_sbox_inst3_xyxx_inst_n68,
         prince_inst_sbox_inst3_xyxx_inst_n67,
         prince_inst_sbox_inst3_xyxx_inst_n66,
         prince_inst_sbox_inst3_xyxx_inst_n65,
         prince_inst_sbox_inst3_xyxx_inst_n64,
         prince_inst_sbox_inst3_xyxx_inst_n63,
         prince_inst_sbox_inst3_xyxx_inst_n62,
         prince_inst_sbox_inst3_xyxx_inst_n61,
         prince_inst_sbox_inst3_xyxx_inst_n60,
         prince_inst_sbox_inst3_xyxx_inst_n59,
         prince_inst_sbox_inst3_xyxx_inst_n58,
         prince_inst_sbox_inst3_xyxx_inst_n57,
         prince_inst_sbox_inst3_xyxx_inst_n56,
         prince_inst_sbox_inst3_xyxx_inst_n55,
         prince_inst_sbox_inst3_xyxx_inst_n54,
         prince_inst_sbox_inst3_xyxx_inst_n53,
         prince_inst_sbox_inst3_xyyy_inst_n61,
         prince_inst_sbox_inst3_xyyy_inst_n60,
         prince_inst_sbox_inst3_xyyy_inst_n59,
         prince_inst_sbox_inst3_xyyy_inst_n58,
         prince_inst_sbox_inst3_xyyy_inst_n57,
         prince_inst_sbox_inst3_xyyy_inst_n56,
         prince_inst_sbox_inst3_xyyy_inst_n55,
         prince_inst_sbox_inst3_xyyy_inst_n54,
         prince_inst_sbox_inst3_xyyy_inst_n53,
         prince_inst_sbox_inst3_xyyy_inst_n52,
         prince_inst_sbox_inst3_xyyy_inst_n51,
         prince_inst_sbox_inst3_xyyy_inst_n50,
         prince_inst_sbox_inst3_xyyy_inst_n49,
         prince_inst_sbox_inst3_xyyy_inst_n48,
         prince_inst_sbox_inst3_xyyy_inst_n47,
         prince_inst_sbox_inst3_xyyy_inst_n46,
         prince_inst_sbox_inst3_xyyy_inst_n45,
         prince_inst_sbox_inst3_xyyy_inst_n44,
         prince_inst_sbox_inst3_xyyy_inst_n43,
         prince_inst_sbox_inst3_xyyy_inst_n42,
         prince_inst_sbox_inst3_yxxx_inst_n64,
         prince_inst_sbox_inst3_yxxx_inst_n63,
         prince_inst_sbox_inst3_yxxx_inst_n62,
         prince_inst_sbox_inst3_yxxx_inst_n61,
         prince_inst_sbox_inst3_yxxx_inst_n60,
         prince_inst_sbox_inst3_yxxx_inst_n59,
         prince_inst_sbox_inst3_yxxx_inst_n58,
         prince_inst_sbox_inst3_yxxx_inst_n57,
         prince_inst_sbox_inst3_yxxx_inst_n56,
         prince_inst_sbox_inst3_yxxx_inst_n55,
         prince_inst_sbox_inst3_yxxx_inst_n54,
         prince_inst_sbox_inst3_yxxx_inst_n53,
         prince_inst_sbox_inst3_yxxx_inst_n52,
         prince_inst_sbox_inst3_yxxx_inst_n51,
         prince_inst_sbox_inst3_yxxx_inst_n50,
         prince_inst_sbox_inst3_yxxx_inst_n49,
         prince_inst_sbox_inst3_yxxx_inst_n48,
         prince_inst_sbox_inst3_yxxx_inst_n47,
         prince_inst_sbox_inst3_yxxx_inst_n46,
         prince_inst_sbox_inst3_yxxx_inst_n45,
         prince_inst_sbox_inst3_yxyy_inst_n67,
         prince_inst_sbox_inst3_yxyy_inst_n66,
         prince_inst_sbox_inst3_yxyy_inst_n65,
         prince_inst_sbox_inst3_yxyy_inst_n64,
         prince_inst_sbox_inst3_yxyy_inst_n63,
         prince_inst_sbox_inst3_yxyy_inst_n62,
         prince_inst_sbox_inst3_yxyy_inst_n61,
         prince_inst_sbox_inst3_yxyy_inst_n60,
         prince_inst_sbox_inst3_yxyy_inst_n59,
         prince_inst_sbox_inst3_yxyy_inst_n58,
         prince_inst_sbox_inst3_yxyy_inst_n57,
         prince_inst_sbox_inst3_yxyy_inst_n56,
         prince_inst_sbox_inst3_yxyy_inst_n55,
         prince_inst_sbox_inst3_yxyy_inst_n54,
         prince_inst_sbox_inst3_yxyy_inst_n53,
         prince_inst_sbox_inst3_yxyy_inst_n52,
         prince_inst_sbox_inst3_yxyy_inst_n51,
         prince_inst_sbox_inst3_yxyy_inst_n50,
         prince_inst_sbox_inst3_yxyy_inst_n49,
         prince_inst_sbox_inst3_yyxy_inst_n75,
         prince_inst_sbox_inst3_yyxy_inst_n74,
         prince_inst_sbox_inst3_yyxy_inst_n73,
         prince_inst_sbox_inst3_yyxy_inst_n72,
         prince_inst_sbox_inst3_yyxy_inst_n71,
         prince_inst_sbox_inst3_yyxy_inst_n70,
         prince_inst_sbox_inst3_yyxy_inst_n69,
         prince_inst_sbox_inst3_yyxy_inst_n68,
         prince_inst_sbox_inst3_yyxy_inst_n67,
         prince_inst_sbox_inst3_yyxy_inst_n66,
         prince_inst_sbox_inst3_yyxy_inst_n65,
         prince_inst_sbox_inst3_yyxy_inst_n64,
         prince_inst_sbox_inst3_yyxy_inst_n63,
         prince_inst_sbox_inst3_yyxy_inst_n62,
         prince_inst_sbox_inst3_yyxy_inst_n61,
         prince_inst_sbox_inst3_yyxy_inst_n60,
         prince_inst_sbox_inst3_yyxy_inst_n59,
         prince_inst_sbox_inst3_yyxy_inst_n58,
         prince_inst_sbox_inst3_yyxy_inst_n57,
         prince_inst_sbox_inst3_yyxy_inst_n56,
         prince_inst_sbox_inst3_yyxy_inst_n55,
         prince_inst_sbox_inst3_yyxy_inst_n54,
         prince_inst_sbox_inst3_yyxy_inst_n53,
         prince_inst_sbox_inst3_yyyx_inst_n58,
         prince_inst_sbox_inst3_yyyx_inst_n57,
         prince_inst_sbox_inst3_yyyx_inst_n56,
         prince_inst_sbox_inst3_yyyx_inst_n55,
         prince_inst_sbox_inst3_yyyx_inst_n54,
         prince_inst_sbox_inst3_yyyx_inst_n53,
         prince_inst_sbox_inst3_yyyx_inst_n52,
         prince_inst_sbox_inst3_yyyx_inst_n51,
         prince_inst_sbox_inst3_yyyx_inst_n50,
         prince_inst_sbox_inst3_yyyx_inst_n49,
         prince_inst_sbox_inst3_yyyx_inst_n48,
         prince_inst_sbox_inst3_yyyx_inst_n47,
         prince_inst_sbox_inst3_yyyx_inst_n46,
         prince_inst_sbox_inst3_yyyx_inst_n45,
         prince_inst_sbox_inst3_yyyx_inst_n44,
         prince_inst_sbox_inst3_yyyx_inst_n43,
         prince_inst_sbox_inst3_yyyx_inst_n42,
         prince_inst_sbox_inst3_c_inst0_msk0_xr,
         prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_msk1_xr,
         prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_msk2_xr,
         prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_msk3_xr,
         prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_msk4_xr,
         prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_msk5_xr,
         prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_msk6_xr,
         prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_msk7_xr,
         prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst0_ax_n6,
         prince_inst_sbox_inst3_c_inst0_ax_n5,
         prince_inst_sbox_inst3_c_inst0_ay_n6,
         prince_inst_sbox_inst3_c_inst0_ay_n5,
         prince_inst_sbox_inst3_c_inst1_msk0_xr,
         prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_msk1_xr,
         prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_msk2_xr,
         prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_msk3_xr,
         prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_msk4_xr,
         prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_msk5_xr,
         prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_msk6_xr,
         prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_msk7_xr,
         prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst1_ax_n6,
         prince_inst_sbox_inst3_c_inst1_ax_n5,
         prince_inst_sbox_inst3_c_inst1_ay_n6,
         prince_inst_sbox_inst3_c_inst1_ay_n5,
         prince_inst_sbox_inst3_c_inst2_msk0_xr,
         prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_msk1_xr,
         prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_msk2_xr,
         prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_msk3_xr,
         prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_msk4_xr,
         prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_msk5_xr,
         prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_msk6_xr,
         prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_msk7_xr,
         prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst2_ax_n6,
         prince_inst_sbox_inst3_c_inst2_ax_n5,
         prince_inst_sbox_inst3_c_inst2_ay_n6,
         prince_inst_sbox_inst3_c_inst2_ay_n5,
         prince_inst_sbox_inst3_c_inst3_msk0_xr,
         prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_msk1_xr,
         prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_msk2_xr,
         prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_msk3_xr,
         prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_msk4_xr,
         prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_msk5_xr,
         prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_msk6_xr,
         prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_msk7_xr,
         prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst3_c_inst3_ax_n6,
         prince_inst_sbox_inst3_c_inst3_ax_n5,
         prince_inst_sbox_inst3_c_inst3_ay_n6,
         prince_inst_sbox_inst3_c_inst3_ay_n5, prince_inst_sbox_inst4_n12,
         prince_inst_sbox_inst4_n11, prince_inst_sbox_inst4_n10,
         prince_inst_sbox_inst4_n9, prince_inst_sbox_inst4_n8,
         prince_inst_sbox_inst4_n7, prince_inst_sbox_inst4_n6,
         prince_inst_sbox_inst4_xxxy_inst_n69,
         prince_inst_sbox_inst4_xxxy_inst_n68,
         prince_inst_sbox_inst4_xxxy_inst_n67,
         prince_inst_sbox_inst4_xxxy_inst_n66,
         prince_inst_sbox_inst4_xxxy_inst_n65,
         prince_inst_sbox_inst4_xxxy_inst_n64,
         prince_inst_sbox_inst4_xxxy_inst_n63,
         prince_inst_sbox_inst4_xxxy_inst_n62,
         prince_inst_sbox_inst4_xxxy_inst_n61,
         prince_inst_sbox_inst4_xxxy_inst_n60,
         prince_inst_sbox_inst4_xxxy_inst_n59,
         prince_inst_sbox_inst4_xxxy_inst_n58,
         prince_inst_sbox_inst4_xxxy_inst_n57,
         prince_inst_sbox_inst4_xxxy_inst_n56,
         prince_inst_sbox_inst4_xxxy_inst_n55,
         prince_inst_sbox_inst4_xxxy_inst_n54,
         prince_inst_sbox_inst4_xxxy_inst_n53,
         prince_inst_sbox_inst4_xxxy_inst_n52,
         prince_inst_sbox_inst4_xxxy_inst_n51,
         prince_inst_sbox_inst4_xxyx_inst_n55,
         prince_inst_sbox_inst4_xxyx_inst_n54,
         prince_inst_sbox_inst4_xxyx_inst_n53,
         prince_inst_sbox_inst4_xxyx_inst_n52,
         prince_inst_sbox_inst4_xxyx_inst_n51,
         prince_inst_sbox_inst4_xxyx_inst_n50,
         prince_inst_sbox_inst4_xxyx_inst_n49,
         prince_inst_sbox_inst4_xxyx_inst_n48,
         prince_inst_sbox_inst4_xxyx_inst_n47,
         prince_inst_sbox_inst4_xxyx_inst_n46,
         prince_inst_sbox_inst4_xxyx_inst_n45,
         prince_inst_sbox_inst4_xxyx_inst_n44,
         prince_inst_sbox_inst4_xxyx_inst_n43,
         prince_inst_sbox_inst4_xxyx_inst_n42,
         prince_inst_sbox_inst4_xxyx_inst_n41,
         prince_inst_sbox_inst4_xxyx_inst_n40,
         prince_inst_sbox_inst4_xxyx_inst_n39,
         prince_inst_sbox_inst4_xxyx_inst_n38,
         prince_inst_sbox_inst4_xyxx_inst_n74,
         prince_inst_sbox_inst4_xyxx_inst_n73,
         prince_inst_sbox_inst4_xyxx_inst_n72,
         prince_inst_sbox_inst4_xyxx_inst_n71,
         prince_inst_sbox_inst4_xyxx_inst_n70,
         prince_inst_sbox_inst4_xyxx_inst_n69,
         prince_inst_sbox_inst4_xyxx_inst_n68,
         prince_inst_sbox_inst4_xyxx_inst_n67,
         prince_inst_sbox_inst4_xyxx_inst_n66,
         prince_inst_sbox_inst4_xyxx_inst_n65,
         prince_inst_sbox_inst4_xyxx_inst_n64,
         prince_inst_sbox_inst4_xyxx_inst_n63,
         prince_inst_sbox_inst4_xyxx_inst_n62,
         prince_inst_sbox_inst4_xyxx_inst_n61,
         prince_inst_sbox_inst4_xyxx_inst_n60,
         prince_inst_sbox_inst4_xyxx_inst_n59,
         prince_inst_sbox_inst4_xyxx_inst_n58,
         prince_inst_sbox_inst4_xyxx_inst_n57,
         prince_inst_sbox_inst4_xyxx_inst_n56,
         prince_inst_sbox_inst4_xyxx_inst_n55,
         prince_inst_sbox_inst4_xyxx_inst_n54,
         prince_inst_sbox_inst4_xyxx_inst_n53,
         prince_inst_sbox_inst4_xyyy_inst_n61,
         prince_inst_sbox_inst4_xyyy_inst_n60,
         prince_inst_sbox_inst4_xyyy_inst_n59,
         prince_inst_sbox_inst4_xyyy_inst_n58,
         prince_inst_sbox_inst4_xyyy_inst_n57,
         prince_inst_sbox_inst4_xyyy_inst_n56,
         prince_inst_sbox_inst4_xyyy_inst_n55,
         prince_inst_sbox_inst4_xyyy_inst_n54,
         prince_inst_sbox_inst4_xyyy_inst_n53,
         prince_inst_sbox_inst4_xyyy_inst_n52,
         prince_inst_sbox_inst4_xyyy_inst_n51,
         prince_inst_sbox_inst4_xyyy_inst_n50,
         prince_inst_sbox_inst4_xyyy_inst_n49,
         prince_inst_sbox_inst4_xyyy_inst_n48,
         prince_inst_sbox_inst4_xyyy_inst_n47,
         prince_inst_sbox_inst4_xyyy_inst_n46,
         prince_inst_sbox_inst4_xyyy_inst_n45,
         prince_inst_sbox_inst4_xyyy_inst_n44,
         prince_inst_sbox_inst4_xyyy_inst_n43,
         prince_inst_sbox_inst4_xyyy_inst_n42,
         prince_inst_sbox_inst4_yxxx_inst_n64,
         prince_inst_sbox_inst4_yxxx_inst_n63,
         prince_inst_sbox_inst4_yxxx_inst_n62,
         prince_inst_sbox_inst4_yxxx_inst_n61,
         prince_inst_sbox_inst4_yxxx_inst_n60,
         prince_inst_sbox_inst4_yxxx_inst_n59,
         prince_inst_sbox_inst4_yxxx_inst_n58,
         prince_inst_sbox_inst4_yxxx_inst_n57,
         prince_inst_sbox_inst4_yxxx_inst_n56,
         prince_inst_sbox_inst4_yxxx_inst_n55,
         prince_inst_sbox_inst4_yxxx_inst_n54,
         prince_inst_sbox_inst4_yxxx_inst_n53,
         prince_inst_sbox_inst4_yxxx_inst_n52,
         prince_inst_sbox_inst4_yxxx_inst_n51,
         prince_inst_sbox_inst4_yxxx_inst_n50,
         prince_inst_sbox_inst4_yxxx_inst_n49,
         prince_inst_sbox_inst4_yxxx_inst_n48,
         prince_inst_sbox_inst4_yxxx_inst_n47,
         prince_inst_sbox_inst4_yxxx_inst_n46,
         prince_inst_sbox_inst4_yxxx_inst_n45,
         prince_inst_sbox_inst4_yxyy_inst_n68,
         prince_inst_sbox_inst4_yxyy_inst_n67,
         prince_inst_sbox_inst4_yxyy_inst_n66,
         prince_inst_sbox_inst4_yxyy_inst_n65,
         prince_inst_sbox_inst4_yxyy_inst_n64,
         prince_inst_sbox_inst4_yxyy_inst_n63,
         prince_inst_sbox_inst4_yxyy_inst_n62,
         prince_inst_sbox_inst4_yxyy_inst_n61,
         prince_inst_sbox_inst4_yxyy_inst_n60,
         prince_inst_sbox_inst4_yxyy_inst_n59,
         prince_inst_sbox_inst4_yxyy_inst_n58,
         prince_inst_sbox_inst4_yxyy_inst_n57,
         prince_inst_sbox_inst4_yxyy_inst_n56,
         prince_inst_sbox_inst4_yxyy_inst_n55,
         prince_inst_sbox_inst4_yxyy_inst_n54,
         prince_inst_sbox_inst4_yxyy_inst_n53,
         prince_inst_sbox_inst4_yxyy_inst_n52,
         prince_inst_sbox_inst4_yxyy_inst_n51,
         prince_inst_sbox_inst4_yxyy_inst_n50,
         prince_inst_sbox_inst4_yxyy_inst_n49,
         prince_inst_sbox_inst4_yyxy_inst_n75,
         prince_inst_sbox_inst4_yyxy_inst_n74,
         prince_inst_sbox_inst4_yyxy_inst_n73,
         prince_inst_sbox_inst4_yyxy_inst_n72,
         prince_inst_sbox_inst4_yyxy_inst_n71,
         prince_inst_sbox_inst4_yyxy_inst_n70,
         prince_inst_sbox_inst4_yyxy_inst_n69,
         prince_inst_sbox_inst4_yyxy_inst_n68,
         prince_inst_sbox_inst4_yyxy_inst_n67,
         prince_inst_sbox_inst4_yyxy_inst_n66,
         prince_inst_sbox_inst4_yyxy_inst_n65,
         prince_inst_sbox_inst4_yyxy_inst_n64,
         prince_inst_sbox_inst4_yyxy_inst_n63,
         prince_inst_sbox_inst4_yyxy_inst_n62,
         prince_inst_sbox_inst4_yyxy_inst_n61,
         prince_inst_sbox_inst4_yyxy_inst_n60,
         prince_inst_sbox_inst4_yyxy_inst_n59,
         prince_inst_sbox_inst4_yyxy_inst_n58,
         prince_inst_sbox_inst4_yyxy_inst_n57,
         prince_inst_sbox_inst4_yyxy_inst_n56,
         prince_inst_sbox_inst4_yyxy_inst_n55,
         prince_inst_sbox_inst4_yyxy_inst_n54,
         prince_inst_sbox_inst4_yyxy_inst_n53,
         prince_inst_sbox_inst4_yyyx_inst_n58,
         prince_inst_sbox_inst4_yyyx_inst_n57,
         prince_inst_sbox_inst4_yyyx_inst_n56,
         prince_inst_sbox_inst4_yyyx_inst_n55,
         prince_inst_sbox_inst4_yyyx_inst_n54,
         prince_inst_sbox_inst4_yyyx_inst_n53,
         prince_inst_sbox_inst4_yyyx_inst_n52,
         prince_inst_sbox_inst4_yyyx_inst_n51,
         prince_inst_sbox_inst4_yyyx_inst_n50,
         prince_inst_sbox_inst4_yyyx_inst_n49,
         prince_inst_sbox_inst4_yyyx_inst_n48,
         prince_inst_sbox_inst4_yyyx_inst_n47,
         prince_inst_sbox_inst4_yyyx_inst_n46,
         prince_inst_sbox_inst4_yyyx_inst_n45,
         prince_inst_sbox_inst4_yyyx_inst_n44,
         prince_inst_sbox_inst4_yyyx_inst_n43,
         prince_inst_sbox_inst4_yyyx_inst_n42,
         prince_inst_sbox_inst4_c_inst0_msk0_xr,
         prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_msk1_xr,
         prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_msk2_xr,
         prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_msk3_xr,
         prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_msk4_xr,
         prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_msk5_xr,
         prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_msk6_xr,
         prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_msk7_xr,
         prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst0_ax_n6,
         prince_inst_sbox_inst4_c_inst0_ax_n5,
         prince_inst_sbox_inst4_c_inst0_ay_n6,
         prince_inst_sbox_inst4_c_inst0_ay_n5,
         prince_inst_sbox_inst4_c_inst1_msk0_xr,
         prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_msk1_xr,
         prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_msk2_xr,
         prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_msk3_xr,
         prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_msk4_xr,
         prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_msk5_xr,
         prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_msk6_xr,
         prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_msk7_xr,
         prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst1_ax_n6,
         prince_inst_sbox_inst4_c_inst1_ax_n5,
         prince_inst_sbox_inst4_c_inst1_ay_n6,
         prince_inst_sbox_inst4_c_inst1_ay_n5,
         prince_inst_sbox_inst4_c_inst2_msk0_xr,
         prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_msk1_xr,
         prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_msk2_xr,
         prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_msk3_xr,
         prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_msk4_xr,
         prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_msk5_xr,
         prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_msk6_xr,
         prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_msk7_xr,
         prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst2_ax_n6,
         prince_inst_sbox_inst4_c_inst2_ax_n5,
         prince_inst_sbox_inst4_c_inst2_ay_n6,
         prince_inst_sbox_inst4_c_inst2_ay_n5,
         prince_inst_sbox_inst4_c_inst3_msk0_xr,
         prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_msk1_xr,
         prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_msk2_xr,
         prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_msk3_xr,
         prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_msk4_xr,
         prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_msk5_xr,
         prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_msk6_xr,
         prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_msk7_xr,
         prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst4_c_inst3_ax_n6,
         prince_inst_sbox_inst4_c_inst3_ax_n5,
         prince_inst_sbox_inst4_c_inst3_ay_n6,
         prince_inst_sbox_inst4_c_inst3_ay_n5, prince_inst_sbox_inst5_n12,
         prince_inst_sbox_inst5_n11, prince_inst_sbox_inst5_n10,
         prince_inst_sbox_inst5_n9, prince_inst_sbox_inst5_n8,
         prince_inst_sbox_inst5_n7, prince_inst_sbox_inst5_n6,
         prince_inst_sbox_inst5_xxxy_inst_n69,
         prince_inst_sbox_inst5_xxxy_inst_n68,
         prince_inst_sbox_inst5_xxxy_inst_n67,
         prince_inst_sbox_inst5_xxxy_inst_n66,
         prince_inst_sbox_inst5_xxxy_inst_n65,
         prince_inst_sbox_inst5_xxxy_inst_n64,
         prince_inst_sbox_inst5_xxxy_inst_n63,
         prince_inst_sbox_inst5_xxxy_inst_n62,
         prince_inst_sbox_inst5_xxxy_inst_n61,
         prince_inst_sbox_inst5_xxxy_inst_n60,
         prince_inst_sbox_inst5_xxxy_inst_n59,
         prince_inst_sbox_inst5_xxxy_inst_n58,
         prince_inst_sbox_inst5_xxxy_inst_n57,
         prince_inst_sbox_inst5_xxxy_inst_n56,
         prince_inst_sbox_inst5_xxxy_inst_n55,
         prince_inst_sbox_inst5_xxxy_inst_n54,
         prince_inst_sbox_inst5_xxxy_inst_n53,
         prince_inst_sbox_inst5_xxxy_inst_n52,
         prince_inst_sbox_inst5_xxxy_inst_n51,
         prince_inst_sbox_inst5_xxyx_inst_n55,
         prince_inst_sbox_inst5_xxyx_inst_n54,
         prince_inst_sbox_inst5_xxyx_inst_n53,
         prince_inst_sbox_inst5_xxyx_inst_n52,
         prince_inst_sbox_inst5_xxyx_inst_n51,
         prince_inst_sbox_inst5_xxyx_inst_n50,
         prince_inst_sbox_inst5_xxyx_inst_n49,
         prince_inst_sbox_inst5_xxyx_inst_n48,
         prince_inst_sbox_inst5_xxyx_inst_n47,
         prince_inst_sbox_inst5_xxyx_inst_n46,
         prince_inst_sbox_inst5_xxyx_inst_n45,
         prince_inst_sbox_inst5_xxyx_inst_n44,
         prince_inst_sbox_inst5_xxyx_inst_n43,
         prince_inst_sbox_inst5_xxyx_inst_n42,
         prince_inst_sbox_inst5_xxyx_inst_n41,
         prince_inst_sbox_inst5_xxyx_inst_n40,
         prince_inst_sbox_inst5_xxyx_inst_n39,
         prince_inst_sbox_inst5_xxyx_inst_n38,
         prince_inst_sbox_inst5_xyxx_inst_n74,
         prince_inst_sbox_inst5_xyxx_inst_n73,
         prince_inst_sbox_inst5_xyxx_inst_n72,
         prince_inst_sbox_inst5_xyxx_inst_n71,
         prince_inst_sbox_inst5_xyxx_inst_n70,
         prince_inst_sbox_inst5_xyxx_inst_n69,
         prince_inst_sbox_inst5_xyxx_inst_n68,
         prince_inst_sbox_inst5_xyxx_inst_n67,
         prince_inst_sbox_inst5_xyxx_inst_n66,
         prince_inst_sbox_inst5_xyxx_inst_n65,
         prince_inst_sbox_inst5_xyxx_inst_n64,
         prince_inst_sbox_inst5_xyxx_inst_n63,
         prince_inst_sbox_inst5_xyxx_inst_n62,
         prince_inst_sbox_inst5_xyxx_inst_n61,
         prince_inst_sbox_inst5_xyxx_inst_n60,
         prince_inst_sbox_inst5_xyxx_inst_n59,
         prince_inst_sbox_inst5_xyxx_inst_n58,
         prince_inst_sbox_inst5_xyxx_inst_n57,
         prince_inst_sbox_inst5_xyxx_inst_n56,
         prince_inst_sbox_inst5_xyxx_inst_n55,
         prince_inst_sbox_inst5_xyxx_inst_n54,
         prince_inst_sbox_inst5_xyxx_inst_n53,
         prince_inst_sbox_inst5_xyyy_inst_n61,
         prince_inst_sbox_inst5_xyyy_inst_n60,
         prince_inst_sbox_inst5_xyyy_inst_n59,
         prince_inst_sbox_inst5_xyyy_inst_n58,
         prince_inst_sbox_inst5_xyyy_inst_n57,
         prince_inst_sbox_inst5_xyyy_inst_n56,
         prince_inst_sbox_inst5_xyyy_inst_n55,
         prince_inst_sbox_inst5_xyyy_inst_n54,
         prince_inst_sbox_inst5_xyyy_inst_n53,
         prince_inst_sbox_inst5_xyyy_inst_n52,
         prince_inst_sbox_inst5_xyyy_inst_n51,
         prince_inst_sbox_inst5_xyyy_inst_n50,
         prince_inst_sbox_inst5_xyyy_inst_n49,
         prince_inst_sbox_inst5_xyyy_inst_n48,
         prince_inst_sbox_inst5_xyyy_inst_n47,
         prince_inst_sbox_inst5_xyyy_inst_n46,
         prince_inst_sbox_inst5_xyyy_inst_n45,
         prince_inst_sbox_inst5_xyyy_inst_n44,
         prince_inst_sbox_inst5_xyyy_inst_n43,
         prince_inst_sbox_inst5_xyyy_inst_n42,
         prince_inst_sbox_inst5_yxxx_inst_n64,
         prince_inst_sbox_inst5_yxxx_inst_n63,
         prince_inst_sbox_inst5_yxxx_inst_n62,
         prince_inst_sbox_inst5_yxxx_inst_n61,
         prince_inst_sbox_inst5_yxxx_inst_n60,
         prince_inst_sbox_inst5_yxxx_inst_n59,
         prince_inst_sbox_inst5_yxxx_inst_n58,
         prince_inst_sbox_inst5_yxxx_inst_n57,
         prince_inst_sbox_inst5_yxxx_inst_n56,
         prince_inst_sbox_inst5_yxxx_inst_n55,
         prince_inst_sbox_inst5_yxxx_inst_n54,
         prince_inst_sbox_inst5_yxxx_inst_n53,
         prince_inst_sbox_inst5_yxxx_inst_n52,
         prince_inst_sbox_inst5_yxxx_inst_n51,
         prince_inst_sbox_inst5_yxxx_inst_n50,
         prince_inst_sbox_inst5_yxxx_inst_n49,
         prince_inst_sbox_inst5_yxxx_inst_n48,
         prince_inst_sbox_inst5_yxxx_inst_n47,
         prince_inst_sbox_inst5_yxxx_inst_n46,
         prince_inst_sbox_inst5_yxxx_inst_n45,
         prince_inst_sbox_inst5_yxyy_inst_n68,
         prince_inst_sbox_inst5_yxyy_inst_n67,
         prince_inst_sbox_inst5_yxyy_inst_n66,
         prince_inst_sbox_inst5_yxyy_inst_n65,
         prince_inst_sbox_inst5_yxyy_inst_n64,
         prince_inst_sbox_inst5_yxyy_inst_n63,
         prince_inst_sbox_inst5_yxyy_inst_n62,
         prince_inst_sbox_inst5_yxyy_inst_n61,
         prince_inst_sbox_inst5_yxyy_inst_n60,
         prince_inst_sbox_inst5_yxyy_inst_n59,
         prince_inst_sbox_inst5_yxyy_inst_n58,
         prince_inst_sbox_inst5_yxyy_inst_n57,
         prince_inst_sbox_inst5_yxyy_inst_n56,
         prince_inst_sbox_inst5_yxyy_inst_n55,
         prince_inst_sbox_inst5_yxyy_inst_n54,
         prince_inst_sbox_inst5_yxyy_inst_n53,
         prince_inst_sbox_inst5_yxyy_inst_n52,
         prince_inst_sbox_inst5_yxyy_inst_n51,
         prince_inst_sbox_inst5_yxyy_inst_n50,
         prince_inst_sbox_inst5_yxyy_inst_n49,
         prince_inst_sbox_inst5_yyxy_inst_n75,
         prince_inst_sbox_inst5_yyxy_inst_n74,
         prince_inst_sbox_inst5_yyxy_inst_n73,
         prince_inst_sbox_inst5_yyxy_inst_n72,
         prince_inst_sbox_inst5_yyxy_inst_n71,
         prince_inst_sbox_inst5_yyxy_inst_n70,
         prince_inst_sbox_inst5_yyxy_inst_n69,
         prince_inst_sbox_inst5_yyxy_inst_n68,
         prince_inst_sbox_inst5_yyxy_inst_n67,
         prince_inst_sbox_inst5_yyxy_inst_n66,
         prince_inst_sbox_inst5_yyxy_inst_n65,
         prince_inst_sbox_inst5_yyxy_inst_n64,
         prince_inst_sbox_inst5_yyxy_inst_n63,
         prince_inst_sbox_inst5_yyxy_inst_n62,
         prince_inst_sbox_inst5_yyxy_inst_n61,
         prince_inst_sbox_inst5_yyxy_inst_n60,
         prince_inst_sbox_inst5_yyxy_inst_n59,
         prince_inst_sbox_inst5_yyxy_inst_n58,
         prince_inst_sbox_inst5_yyxy_inst_n57,
         prince_inst_sbox_inst5_yyxy_inst_n56,
         prince_inst_sbox_inst5_yyxy_inst_n55,
         prince_inst_sbox_inst5_yyxy_inst_n54,
         prince_inst_sbox_inst5_yyxy_inst_n53,
         prince_inst_sbox_inst5_yyyx_inst_n58,
         prince_inst_sbox_inst5_yyyx_inst_n57,
         prince_inst_sbox_inst5_yyyx_inst_n56,
         prince_inst_sbox_inst5_yyyx_inst_n55,
         prince_inst_sbox_inst5_yyyx_inst_n54,
         prince_inst_sbox_inst5_yyyx_inst_n53,
         prince_inst_sbox_inst5_yyyx_inst_n52,
         prince_inst_sbox_inst5_yyyx_inst_n51,
         prince_inst_sbox_inst5_yyyx_inst_n50,
         prince_inst_sbox_inst5_yyyx_inst_n49,
         prince_inst_sbox_inst5_yyyx_inst_n48,
         prince_inst_sbox_inst5_yyyx_inst_n47,
         prince_inst_sbox_inst5_yyyx_inst_n46,
         prince_inst_sbox_inst5_yyyx_inst_n45,
         prince_inst_sbox_inst5_yyyx_inst_n44,
         prince_inst_sbox_inst5_yyyx_inst_n43,
         prince_inst_sbox_inst5_yyyx_inst_n42,
         prince_inst_sbox_inst5_c_inst0_msk0_xr,
         prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_msk1_xr,
         prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_msk2_xr,
         prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_msk3_xr,
         prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_msk4_xr,
         prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_msk5_xr,
         prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_msk6_xr,
         prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_msk7_xr,
         prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst0_ax_n6,
         prince_inst_sbox_inst5_c_inst0_ax_n5,
         prince_inst_sbox_inst5_c_inst0_ay_n6,
         prince_inst_sbox_inst5_c_inst0_ay_n5,
         prince_inst_sbox_inst5_c_inst1_msk0_xr,
         prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_msk1_xr,
         prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_msk2_xr,
         prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_msk3_xr,
         prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_msk4_xr,
         prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_msk5_xr,
         prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_msk6_xr,
         prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_msk7_xr,
         prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst1_ax_n6,
         prince_inst_sbox_inst5_c_inst1_ax_n5,
         prince_inst_sbox_inst5_c_inst1_ay_n6,
         prince_inst_sbox_inst5_c_inst1_ay_n5,
         prince_inst_sbox_inst5_c_inst2_msk0_xr,
         prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_msk1_xr,
         prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_msk2_xr,
         prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_msk3_xr,
         prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_msk4_xr,
         prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_msk5_xr,
         prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_msk6_xr,
         prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_msk7_xr,
         prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst2_ax_n6,
         prince_inst_sbox_inst5_c_inst2_ax_n5,
         prince_inst_sbox_inst5_c_inst2_ay_n6,
         prince_inst_sbox_inst5_c_inst2_ay_n5,
         prince_inst_sbox_inst5_c_inst3_msk0_xr,
         prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_msk1_xr,
         prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_msk2_xr,
         prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_msk3_xr,
         prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_msk4_xr,
         prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_msk5_xr,
         prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_msk6_xr,
         prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_msk7_xr,
         prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst5_c_inst3_ax_n6,
         prince_inst_sbox_inst5_c_inst3_ax_n5,
         prince_inst_sbox_inst5_c_inst3_ay_n6,
         prince_inst_sbox_inst5_c_inst3_ay_n5, prince_inst_sbox_inst6_n12,
         prince_inst_sbox_inst6_n11, prince_inst_sbox_inst6_n10,
         prince_inst_sbox_inst6_n9, prince_inst_sbox_inst6_n8,
         prince_inst_sbox_inst6_n7, prince_inst_sbox_inst6_n6,
         prince_inst_sbox_inst6_xxxy_inst_n69,
         prince_inst_sbox_inst6_xxxy_inst_n68,
         prince_inst_sbox_inst6_xxxy_inst_n67,
         prince_inst_sbox_inst6_xxxy_inst_n66,
         prince_inst_sbox_inst6_xxxy_inst_n65,
         prince_inst_sbox_inst6_xxxy_inst_n64,
         prince_inst_sbox_inst6_xxxy_inst_n63,
         prince_inst_sbox_inst6_xxxy_inst_n62,
         prince_inst_sbox_inst6_xxxy_inst_n61,
         prince_inst_sbox_inst6_xxxy_inst_n60,
         prince_inst_sbox_inst6_xxxy_inst_n59,
         prince_inst_sbox_inst6_xxxy_inst_n58,
         prince_inst_sbox_inst6_xxxy_inst_n57,
         prince_inst_sbox_inst6_xxxy_inst_n56,
         prince_inst_sbox_inst6_xxxy_inst_n55,
         prince_inst_sbox_inst6_xxxy_inst_n54,
         prince_inst_sbox_inst6_xxxy_inst_n53,
         prince_inst_sbox_inst6_xxxy_inst_n52,
         prince_inst_sbox_inst6_xxxy_inst_n51,
         prince_inst_sbox_inst6_xxyx_inst_n55,
         prince_inst_sbox_inst6_xxyx_inst_n54,
         prince_inst_sbox_inst6_xxyx_inst_n53,
         prince_inst_sbox_inst6_xxyx_inst_n52,
         prince_inst_sbox_inst6_xxyx_inst_n51,
         prince_inst_sbox_inst6_xxyx_inst_n50,
         prince_inst_sbox_inst6_xxyx_inst_n49,
         prince_inst_sbox_inst6_xxyx_inst_n48,
         prince_inst_sbox_inst6_xxyx_inst_n47,
         prince_inst_sbox_inst6_xxyx_inst_n46,
         prince_inst_sbox_inst6_xxyx_inst_n45,
         prince_inst_sbox_inst6_xxyx_inst_n44,
         prince_inst_sbox_inst6_xxyx_inst_n43,
         prince_inst_sbox_inst6_xxyx_inst_n42,
         prince_inst_sbox_inst6_xxyx_inst_n41,
         prince_inst_sbox_inst6_xxyx_inst_n40,
         prince_inst_sbox_inst6_xxyx_inst_n39,
         prince_inst_sbox_inst6_xxyx_inst_n38,
         prince_inst_sbox_inst6_xyxx_inst_n74,
         prince_inst_sbox_inst6_xyxx_inst_n73,
         prince_inst_sbox_inst6_xyxx_inst_n72,
         prince_inst_sbox_inst6_xyxx_inst_n71,
         prince_inst_sbox_inst6_xyxx_inst_n70,
         prince_inst_sbox_inst6_xyxx_inst_n69,
         prince_inst_sbox_inst6_xyxx_inst_n68,
         prince_inst_sbox_inst6_xyxx_inst_n67,
         prince_inst_sbox_inst6_xyxx_inst_n66,
         prince_inst_sbox_inst6_xyxx_inst_n65,
         prince_inst_sbox_inst6_xyxx_inst_n64,
         prince_inst_sbox_inst6_xyxx_inst_n63,
         prince_inst_sbox_inst6_xyxx_inst_n62,
         prince_inst_sbox_inst6_xyxx_inst_n61,
         prince_inst_sbox_inst6_xyxx_inst_n60,
         prince_inst_sbox_inst6_xyxx_inst_n59,
         prince_inst_sbox_inst6_xyxx_inst_n58,
         prince_inst_sbox_inst6_xyxx_inst_n57,
         prince_inst_sbox_inst6_xyxx_inst_n56,
         prince_inst_sbox_inst6_xyxx_inst_n55,
         prince_inst_sbox_inst6_xyxx_inst_n54,
         prince_inst_sbox_inst6_xyxx_inst_n53,
         prince_inst_sbox_inst6_xyyy_inst_n61,
         prince_inst_sbox_inst6_xyyy_inst_n60,
         prince_inst_sbox_inst6_xyyy_inst_n59,
         prince_inst_sbox_inst6_xyyy_inst_n58,
         prince_inst_sbox_inst6_xyyy_inst_n57,
         prince_inst_sbox_inst6_xyyy_inst_n56,
         prince_inst_sbox_inst6_xyyy_inst_n55,
         prince_inst_sbox_inst6_xyyy_inst_n54,
         prince_inst_sbox_inst6_xyyy_inst_n53,
         prince_inst_sbox_inst6_xyyy_inst_n52,
         prince_inst_sbox_inst6_xyyy_inst_n51,
         prince_inst_sbox_inst6_xyyy_inst_n50,
         prince_inst_sbox_inst6_xyyy_inst_n49,
         prince_inst_sbox_inst6_xyyy_inst_n48,
         prince_inst_sbox_inst6_xyyy_inst_n47,
         prince_inst_sbox_inst6_xyyy_inst_n46,
         prince_inst_sbox_inst6_xyyy_inst_n45,
         prince_inst_sbox_inst6_xyyy_inst_n44,
         prince_inst_sbox_inst6_xyyy_inst_n43,
         prince_inst_sbox_inst6_xyyy_inst_n42,
         prince_inst_sbox_inst6_yxxx_inst_n64,
         prince_inst_sbox_inst6_yxxx_inst_n63,
         prince_inst_sbox_inst6_yxxx_inst_n62,
         prince_inst_sbox_inst6_yxxx_inst_n61,
         prince_inst_sbox_inst6_yxxx_inst_n60,
         prince_inst_sbox_inst6_yxxx_inst_n59,
         prince_inst_sbox_inst6_yxxx_inst_n58,
         prince_inst_sbox_inst6_yxxx_inst_n57,
         prince_inst_sbox_inst6_yxxx_inst_n56,
         prince_inst_sbox_inst6_yxxx_inst_n55,
         prince_inst_sbox_inst6_yxxx_inst_n54,
         prince_inst_sbox_inst6_yxxx_inst_n53,
         prince_inst_sbox_inst6_yxxx_inst_n52,
         prince_inst_sbox_inst6_yxxx_inst_n51,
         prince_inst_sbox_inst6_yxxx_inst_n50,
         prince_inst_sbox_inst6_yxxx_inst_n49,
         prince_inst_sbox_inst6_yxxx_inst_n48,
         prince_inst_sbox_inst6_yxxx_inst_n47,
         prince_inst_sbox_inst6_yxxx_inst_n46,
         prince_inst_sbox_inst6_yxxx_inst_n45,
         prince_inst_sbox_inst6_yxyy_inst_n68,
         prince_inst_sbox_inst6_yxyy_inst_n67,
         prince_inst_sbox_inst6_yxyy_inst_n66,
         prince_inst_sbox_inst6_yxyy_inst_n65,
         prince_inst_sbox_inst6_yxyy_inst_n64,
         prince_inst_sbox_inst6_yxyy_inst_n63,
         prince_inst_sbox_inst6_yxyy_inst_n62,
         prince_inst_sbox_inst6_yxyy_inst_n61,
         prince_inst_sbox_inst6_yxyy_inst_n60,
         prince_inst_sbox_inst6_yxyy_inst_n59,
         prince_inst_sbox_inst6_yxyy_inst_n58,
         prince_inst_sbox_inst6_yxyy_inst_n57,
         prince_inst_sbox_inst6_yxyy_inst_n56,
         prince_inst_sbox_inst6_yxyy_inst_n55,
         prince_inst_sbox_inst6_yxyy_inst_n54,
         prince_inst_sbox_inst6_yxyy_inst_n53,
         prince_inst_sbox_inst6_yxyy_inst_n52,
         prince_inst_sbox_inst6_yxyy_inst_n51,
         prince_inst_sbox_inst6_yxyy_inst_n50,
         prince_inst_sbox_inst6_yxyy_inst_n49,
         prince_inst_sbox_inst6_yyxy_inst_n75,
         prince_inst_sbox_inst6_yyxy_inst_n74,
         prince_inst_sbox_inst6_yyxy_inst_n73,
         prince_inst_sbox_inst6_yyxy_inst_n72,
         prince_inst_sbox_inst6_yyxy_inst_n71,
         prince_inst_sbox_inst6_yyxy_inst_n70,
         prince_inst_sbox_inst6_yyxy_inst_n69,
         prince_inst_sbox_inst6_yyxy_inst_n68,
         prince_inst_sbox_inst6_yyxy_inst_n67,
         prince_inst_sbox_inst6_yyxy_inst_n66,
         prince_inst_sbox_inst6_yyxy_inst_n65,
         prince_inst_sbox_inst6_yyxy_inst_n64,
         prince_inst_sbox_inst6_yyxy_inst_n63,
         prince_inst_sbox_inst6_yyxy_inst_n62,
         prince_inst_sbox_inst6_yyxy_inst_n61,
         prince_inst_sbox_inst6_yyxy_inst_n60,
         prince_inst_sbox_inst6_yyxy_inst_n59,
         prince_inst_sbox_inst6_yyxy_inst_n58,
         prince_inst_sbox_inst6_yyxy_inst_n57,
         prince_inst_sbox_inst6_yyxy_inst_n56,
         prince_inst_sbox_inst6_yyxy_inst_n55,
         prince_inst_sbox_inst6_yyxy_inst_n54,
         prince_inst_sbox_inst6_yyxy_inst_n53,
         prince_inst_sbox_inst6_yyyx_inst_n58,
         prince_inst_sbox_inst6_yyyx_inst_n57,
         prince_inst_sbox_inst6_yyyx_inst_n56,
         prince_inst_sbox_inst6_yyyx_inst_n55,
         prince_inst_sbox_inst6_yyyx_inst_n54,
         prince_inst_sbox_inst6_yyyx_inst_n53,
         prince_inst_sbox_inst6_yyyx_inst_n52,
         prince_inst_sbox_inst6_yyyx_inst_n51,
         prince_inst_sbox_inst6_yyyx_inst_n50,
         prince_inst_sbox_inst6_yyyx_inst_n49,
         prince_inst_sbox_inst6_yyyx_inst_n48,
         prince_inst_sbox_inst6_yyyx_inst_n47,
         prince_inst_sbox_inst6_yyyx_inst_n46,
         prince_inst_sbox_inst6_yyyx_inst_n45,
         prince_inst_sbox_inst6_yyyx_inst_n44,
         prince_inst_sbox_inst6_yyyx_inst_n43,
         prince_inst_sbox_inst6_yyyx_inst_n42,
         prince_inst_sbox_inst6_c_inst0_msk0_xr,
         prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_msk1_xr,
         prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_msk2_xr,
         prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_msk3_xr,
         prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_msk4_xr,
         prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_msk5_xr,
         prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_msk6_xr,
         prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_msk7_xr,
         prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst0_ax_n6,
         prince_inst_sbox_inst6_c_inst0_ax_n5,
         prince_inst_sbox_inst6_c_inst0_ay_n6,
         prince_inst_sbox_inst6_c_inst0_ay_n5,
         prince_inst_sbox_inst6_c_inst1_msk0_xr,
         prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_msk1_xr,
         prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_msk2_xr,
         prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_msk3_xr,
         prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_msk4_xr,
         prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_msk5_xr,
         prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_msk6_xr,
         prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_msk7_xr,
         prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst1_ax_n6,
         prince_inst_sbox_inst6_c_inst1_ax_n5,
         prince_inst_sbox_inst6_c_inst1_ay_n6,
         prince_inst_sbox_inst6_c_inst1_ay_n5,
         prince_inst_sbox_inst6_c_inst2_msk0_xr,
         prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_msk1_xr,
         prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_msk2_xr,
         prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_msk3_xr,
         prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_msk4_xr,
         prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_msk5_xr,
         prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_msk6_xr,
         prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_msk7_xr,
         prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst2_ax_n6,
         prince_inst_sbox_inst6_c_inst2_ax_n5,
         prince_inst_sbox_inst6_c_inst2_ay_n6,
         prince_inst_sbox_inst6_c_inst2_ay_n5,
         prince_inst_sbox_inst6_c_inst3_msk0_xr,
         prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_msk1_xr,
         prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_msk2_xr,
         prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_msk3_xr,
         prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_msk4_xr,
         prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_msk5_xr,
         prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_msk6_xr,
         prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_msk7_xr,
         prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst6_c_inst3_ax_n6,
         prince_inst_sbox_inst6_c_inst3_ax_n5,
         prince_inst_sbox_inst6_c_inst3_ay_n6,
         prince_inst_sbox_inst6_c_inst3_ay_n5, prince_inst_sbox_inst7_n10,
         prince_inst_sbox_inst7_n9, prince_inst_sbox_inst7_n8,
         prince_inst_sbox_inst7_n7, prince_inst_sbox_inst7_n6,
         prince_inst_sbox_inst7_xxxy_inst_n70,
         prince_inst_sbox_inst7_xxxy_inst_n69,
         prince_inst_sbox_inst7_xxxy_inst_n68,
         prince_inst_sbox_inst7_xxxy_inst_n67,
         prince_inst_sbox_inst7_xxxy_inst_n66,
         prince_inst_sbox_inst7_xxxy_inst_n65,
         prince_inst_sbox_inst7_xxxy_inst_n64,
         prince_inst_sbox_inst7_xxxy_inst_n63,
         prince_inst_sbox_inst7_xxxy_inst_n62,
         prince_inst_sbox_inst7_xxxy_inst_n61,
         prince_inst_sbox_inst7_xxxy_inst_n60,
         prince_inst_sbox_inst7_xxxy_inst_n59,
         prince_inst_sbox_inst7_xxxy_inst_n58,
         prince_inst_sbox_inst7_xxxy_inst_n57,
         prince_inst_sbox_inst7_xxxy_inst_n56,
         prince_inst_sbox_inst7_xxxy_inst_n55,
         prince_inst_sbox_inst7_xxxy_inst_n54,
         prince_inst_sbox_inst7_xxxy_inst_n53,
         prince_inst_sbox_inst7_xxxy_inst_n52,
         prince_inst_sbox_inst7_xxxy_inst_n51,
         prince_inst_sbox_inst7_xxyx_inst_n55,
         prince_inst_sbox_inst7_xxyx_inst_n54,
         prince_inst_sbox_inst7_xxyx_inst_n53,
         prince_inst_sbox_inst7_xxyx_inst_n52,
         prince_inst_sbox_inst7_xxyx_inst_n51,
         prince_inst_sbox_inst7_xxyx_inst_n50,
         prince_inst_sbox_inst7_xxyx_inst_n49,
         prince_inst_sbox_inst7_xxyx_inst_n48,
         prince_inst_sbox_inst7_xxyx_inst_n47,
         prince_inst_sbox_inst7_xxyx_inst_n46,
         prince_inst_sbox_inst7_xxyx_inst_n45,
         prince_inst_sbox_inst7_xxyx_inst_n44,
         prince_inst_sbox_inst7_xxyx_inst_n43,
         prince_inst_sbox_inst7_xxyx_inst_n42,
         prince_inst_sbox_inst7_xxyx_inst_n41,
         prince_inst_sbox_inst7_xxyx_inst_n40,
         prince_inst_sbox_inst7_xxyx_inst_n39,
         prince_inst_sbox_inst7_xxyx_inst_n38,
         prince_inst_sbox_inst7_xyxx_inst_n74,
         prince_inst_sbox_inst7_xyxx_inst_n73,
         prince_inst_sbox_inst7_xyxx_inst_n72,
         prince_inst_sbox_inst7_xyxx_inst_n71,
         prince_inst_sbox_inst7_xyxx_inst_n70,
         prince_inst_sbox_inst7_xyxx_inst_n69,
         prince_inst_sbox_inst7_xyxx_inst_n68,
         prince_inst_sbox_inst7_xyxx_inst_n67,
         prince_inst_sbox_inst7_xyxx_inst_n66,
         prince_inst_sbox_inst7_xyxx_inst_n65,
         prince_inst_sbox_inst7_xyxx_inst_n64,
         prince_inst_sbox_inst7_xyxx_inst_n63,
         prince_inst_sbox_inst7_xyxx_inst_n62,
         prince_inst_sbox_inst7_xyxx_inst_n61,
         prince_inst_sbox_inst7_xyxx_inst_n60,
         prince_inst_sbox_inst7_xyxx_inst_n59,
         prince_inst_sbox_inst7_xyxx_inst_n58,
         prince_inst_sbox_inst7_xyxx_inst_n57,
         prince_inst_sbox_inst7_xyxx_inst_n56,
         prince_inst_sbox_inst7_xyxx_inst_n55,
         prince_inst_sbox_inst7_xyxx_inst_n54,
         prince_inst_sbox_inst7_xyxx_inst_n53,
         prince_inst_sbox_inst7_xyyy_inst_n61,
         prince_inst_sbox_inst7_xyyy_inst_n60,
         prince_inst_sbox_inst7_xyyy_inst_n59,
         prince_inst_sbox_inst7_xyyy_inst_n58,
         prince_inst_sbox_inst7_xyyy_inst_n57,
         prince_inst_sbox_inst7_xyyy_inst_n56,
         prince_inst_sbox_inst7_xyyy_inst_n55,
         prince_inst_sbox_inst7_xyyy_inst_n54,
         prince_inst_sbox_inst7_xyyy_inst_n53,
         prince_inst_sbox_inst7_xyyy_inst_n52,
         prince_inst_sbox_inst7_xyyy_inst_n51,
         prince_inst_sbox_inst7_xyyy_inst_n50,
         prince_inst_sbox_inst7_xyyy_inst_n49,
         prince_inst_sbox_inst7_xyyy_inst_n48,
         prince_inst_sbox_inst7_xyyy_inst_n47,
         prince_inst_sbox_inst7_xyyy_inst_n46,
         prince_inst_sbox_inst7_xyyy_inst_n45,
         prince_inst_sbox_inst7_xyyy_inst_n44,
         prince_inst_sbox_inst7_xyyy_inst_n43,
         prince_inst_sbox_inst7_xyyy_inst_n42,
         prince_inst_sbox_inst7_yxxx_inst_n64,
         prince_inst_sbox_inst7_yxxx_inst_n63,
         prince_inst_sbox_inst7_yxxx_inst_n62,
         prince_inst_sbox_inst7_yxxx_inst_n61,
         prince_inst_sbox_inst7_yxxx_inst_n60,
         prince_inst_sbox_inst7_yxxx_inst_n59,
         prince_inst_sbox_inst7_yxxx_inst_n58,
         prince_inst_sbox_inst7_yxxx_inst_n57,
         prince_inst_sbox_inst7_yxxx_inst_n56,
         prince_inst_sbox_inst7_yxxx_inst_n55,
         prince_inst_sbox_inst7_yxxx_inst_n54,
         prince_inst_sbox_inst7_yxxx_inst_n53,
         prince_inst_sbox_inst7_yxxx_inst_n52,
         prince_inst_sbox_inst7_yxxx_inst_n51,
         prince_inst_sbox_inst7_yxxx_inst_n50,
         prince_inst_sbox_inst7_yxxx_inst_n49,
         prince_inst_sbox_inst7_yxxx_inst_n48,
         prince_inst_sbox_inst7_yxxx_inst_n47,
         prince_inst_sbox_inst7_yxxx_inst_n46,
         prince_inst_sbox_inst7_yxxx_inst_n45,
         prince_inst_sbox_inst7_yxyy_inst_n67,
         prince_inst_sbox_inst7_yxyy_inst_n66,
         prince_inst_sbox_inst7_yxyy_inst_n65,
         prince_inst_sbox_inst7_yxyy_inst_n64,
         prince_inst_sbox_inst7_yxyy_inst_n63,
         prince_inst_sbox_inst7_yxyy_inst_n62,
         prince_inst_sbox_inst7_yxyy_inst_n61,
         prince_inst_sbox_inst7_yxyy_inst_n60,
         prince_inst_sbox_inst7_yxyy_inst_n59,
         prince_inst_sbox_inst7_yxyy_inst_n58,
         prince_inst_sbox_inst7_yxyy_inst_n57,
         prince_inst_sbox_inst7_yxyy_inst_n56,
         prince_inst_sbox_inst7_yxyy_inst_n55,
         prince_inst_sbox_inst7_yxyy_inst_n54,
         prince_inst_sbox_inst7_yxyy_inst_n53,
         prince_inst_sbox_inst7_yxyy_inst_n52,
         prince_inst_sbox_inst7_yxyy_inst_n51,
         prince_inst_sbox_inst7_yxyy_inst_n50,
         prince_inst_sbox_inst7_yxyy_inst_n49,
         prince_inst_sbox_inst7_yyxy_inst_n75,
         prince_inst_sbox_inst7_yyxy_inst_n74,
         prince_inst_sbox_inst7_yyxy_inst_n73,
         prince_inst_sbox_inst7_yyxy_inst_n72,
         prince_inst_sbox_inst7_yyxy_inst_n71,
         prince_inst_sbox_inst7_yyxy_inst_n70,
         prince_inst_sbox_inst7_yyxy_inst_n69,
         prince_inst_sbox_inst7_yyxy_inst_n68,
         prince_inst_sbox_inst7_yyxy_inst_n67,
         prince_inst_sbox_inst7_yyxy_inst_n66,
         prince_inst_sbox_inst7_yyxy_inst_n65,
         prince_inst_sbox_inst7_yyxy_inst_n64,
         prince_inst_sbox_inst7_yyxy_inst_n63,
         prince_inst_sbox_inst7_yyxy_inst_n62,
         prince_inst_sbox_inst7_yyxy_inst_n61,
         prince_inst_sbox_inst7_yyxy_inst_n60,
         prince_inst_sbox_inst7_yyxy_inst_n59,
         prince_inst_sbox_inst7_yyxy_inst_n58,
         prince_inst_sbox_inst7_yyxy_inst_n57,
         prince_inst_sbox_inst7_yyxy_inst_n56,
         prince_inst_sbox_inst7_yyxy_inst_n55,
         prince_inst_sbox_inst7_yyxy_inst_n54,
         prince_inst_sbox_inst7_yyxy_inst_n53,
         prince_inst_sbox_inst7_yyyx_inst_n58,
         prince_inst_sbox_inst7_yyyx_inst_n57,
         prince_inst_sbox_inst7_yyyx_inst_n56,
         prince_inst_sbox_inst7_yyyx_inst_n55,
         prince_inst_sbox_inst7_yyyx_inst_n54,
         prince_inst_sbox_inst7_yyyx_inst_n53,
         prince_inst_sbox_inst7_yyyx_inst_n52,
         prince_inst_sbox_inst7_yyyx_inst_n51,
         prince_inst_sbox_inst7_yyyx_inst_n50,
         prince_inst_sbox_inst7_yyyx_inst_n49,
         prince_inst_sbox_inst7_yyyx_inst_n48,
         prince_inst_sbox_inst7_yyyx_inst_n47,
         prince_inst_sbox_inst7_yyyx_inst_n46,
         prince_inst_sbox_inst7_yyyx_inst_n45,
         prince_inst_sbox_inst7_yyyx_inst_n44,
         prince_inst_sbox_inst7_yyyx_inst_n43,
         prince_inst_sbox_inst7_yyyx_inst_n42,
         prince_inst_sbox_inst7_c_inst0_msk0_xr,
         prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_msk1_xr,
         prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_msk2_xr,
         prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_msk3_xr,
         prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_msk4_xr,
         prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_msk5_xr,
         prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_msk6_xr,
         prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_msk7_xr,
         prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst0_ax_n6,
         prince_inst_sbox_inst7_c_inst0_ax_n5,
         prince_inst_sbox_inst7_c_inst0_ay_n6,
         prince_inst_sbox_inst7_c_inst0_ay_n5,
         prince_inst_sbox_inst7_c_inst1_msk0_xr,
         prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_msk1_xr,
         prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_msk2_xr,
         prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_msk3_xr,
         prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_msk4_xr,
         prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_msk5_xr,
         prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_msk6_xr,
         prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_msk7_xr,
         prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst1_ax_n6,
         prince_inst_sbox_inst7_c_inst1_ax_n5,
         prince_inst_sbox_inst7_c_inst1_ay_n6,
         prince_inst_sbox_inst7_c_inst1_ay_n5,
         prince_inst_sbox_inst7_c_inst2_msk0_xr,
         prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_msk1_xr,
         prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_msk2_xr,
         prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_msk3_xr,
         prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_msk4_xr,
         prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_msk5_xr,
         prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_msk6_xr,
         prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_msk7_xr,
         prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst2_ax_n6,
         prince_inst_sbox_inst7_c_inst2_ax_n5,
         prince_inst_sbox_inst7_c_inst2_ay_n6,
         prince_inst_sbox_inst7_c_inst2_ay_n5,
         prince_inst_sbox_inst7_c_inst3_msk0_xr,
         prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_msk1_xr,
         prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_msk2_xr,
         prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_msk3_xr,
         prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_msk4_xr,
         prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_msk5_xr,
         prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_msk6_xr,
         prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_msk7_xr,
         prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst7_c_inst3_ax_n6,
         prince_inst_sbox_inst7_c_inst3_ax_n5,
         prince_inst_sbox_inst7_c_inst3_ay_n6,
         prince_inst_sbox_inst7_c_inst3_ay_n5, prince_inst_sbox_inst8_n10,
         prince_inst_sbox_inst8_n9, prince_inst_sbox_inst8_n8,
         prince_inst_sbox_inst8_n7, prince_inst_sbox_inst8_n6,
         prince_inst_sbox_inst8_xxxy_inst_n69,
         prince_inst_sbox_inst8_xxxy_inst_n68,
         prince_inst_sbox_inst8_xxxy_inst_n67,
         prince_inst_sbox_inst8_xxxy_inst_n66,
         prince_inst_sbox_inst8_xxxy_inst_n65,
         prince_inst_sbox_inst8_xxxy_inst_n64,
         prince_inst_sbox_inst8_xxxy_inst_n63,
         prince_inst_sbox_inst8_xxxy_inst_n62,
         prince_inst_sbox_inst8_xxxy_inst_n61,
         prince_inst_sbox_inst8_xxxy_inst_n60,
         prince_inst_sbox_inst8_xxxy_inst_n59,
         prince_inst_sbox_inst8_xxxy_inst_n58,
         prince_inst_sbox_inst8_xxxy_inst_n57,
         prince_inst_sbox_inst8_xxxy_inst_n56,
         prince_inst_sbox_inst8_xxxy_inst_n55,
         prince_inst_sbox_inst8_xxxy_inst_n54,
         prince_inst_sbox_inst8_xxxy_inst_n53,
         prince_inst_sbox_inst8_xxxy_inst_n52,
         prince_inst_sbox_inst8_xxxy_inst_n51,
         prince_inst_sbox_inst8_xxyx_inst_n55,
         prince_inst_sbox_inst8_xxyx_inst_n54,
         prince_inst_sbox_inst8_xxyx_inst_n53,
         prince_inst_sbox_inst8_xxyx_inst_n52,
         prince_inst_sbox_inst8_xxyx_inst_n51,
         prince_inst_sbox_inst8_xxyx_inst_n50,
         prince_inst_sbox_inst8_xxyx_inst_n49,
         prince_inst_sbox_inst8_xxyx_inst_n48,
         prince_inst_sbox_inst8_xxyx_inst_n47,
         prince_inst_sbox_inst8_xxyx_inst_n46,
         prince_inst_sbox_inst8_xxyx_inst_n45,
         prince_inst_sbox_inst8_xxyx_inst_n44,
         prince_inst_sbox_inst8_xxyx_inst_n43,
         prince_inst_sbox_inst8_xxyx_inst_n42,
         prince_inst_sbox_inst8_xxyx_inst_n41,
         prince_inst_sbox_inst8_xxyx_inst_n40,
         prince_inst_sbox_inst8_xxyx_inst_n39,
         prince_inst_sbox_inst8_xxyx_inst_n38,
         prince_inst_sbox_inst8_xyxx_inst_n74,
         prince_inst_sbox_inst8_xyxx_inst_n73,
         prince_inst_sbox_inst8_xyxx_inst_n72,
         prince_inst_sbox_inst8_xyxx_inst_n71,
         prince_inst_sbox_inst8_xyxx_inst_n70,
         prince_inst_sbox_inst8_xyxx_inst_n69,
         prince_inst_sbox_inst8_xyxx_inst_n68,
         prince_inst_sbox_inst8_xyxx_inst_n67,
         prince_inst_sbox_inst8_xyxx_inst_n66,
         prince_inst_sbox_inst8_xyxx_inst_n65,
         prince_inst_sbox_inst8_xyxx_inst_n64,
         prince_inst_sbox_inst8_xyxx_inst_n63,
         prince_inst_sbox_inst8_xyxx_inst_n62,
         prince_inst_sbox_inst8_xyxx_inst_n61,
         prince_inst_sbox_inst8_xyxx_inst_n60,
         prince_inst_sbox_inst8_xyxx_inst_n59,
         prince_inst_sbox_inst8_xyxx_inst_n58,
         prince_inst_sbox_inst8_xyxx_inst_n57,
         prince_inst_sbox_inst8_xyxx_inst_n56,
         prince_inst_sbox_inst8_xyxx_inst_n55,
         prince_inst_sbox_inst8_xyxx_inst_n54,
         prince_inst_sbox_inst8_xyxx_inst_n53,
         prince_inst_sbox_inst8_xyyy_inst_n61,
         prince_inst_sbox_inst8_xyyy_inst_n60,
         prince_inst_sbox_inst8_xyyy_inst_n59,
         prince_inst_sbox_inst8_xyyy_inst_n58,
         prince_inst_sbox_inst8_xyyy_inst_n57,
         prince_inst_sbox_inst8_xyyy_inst_n56,
         prince_inst_sbox_inst8_xyyy_inst_n55,
         prince_inst_sbox_inst8_xyyy_inst_n54,
         prince_inst_sbox_inst8_xyyy_inst_n53,
         prince_inst_sbox_inst8_xyyy_inst_n52,
         prince_inst_sbox_inst8_xyyy_inst_n51,
         prince_inst_sbox_inst8_xyyy_inst_n50,
         prince_inst_sbox_inst8_xyyy_inst_n49,
         prince_inst_sbox_inst8_xyyy_inst_n48,
         prince_inst_sbox_inst8_xyyy_inst_n47,
         prince_inst_sbox_inst8_xyyy_inst_n46,
         prince_inst_sbox_inst8_xyyy_inst_n45,
         prince_inst_sbox_inst8_xyyy_inst_n44,
         prince_inst_sbox_inst8_xyyy_inst_n43,
         prince_inst_sbox_inst8_xyyy_inst_n42,
         prince_inst_sbox_inst8_yxxx_inst_n64,
         prince_inst_sbox_inst8_yxxx_inst_n63,
         prince_inst_sbox_inst8_yxxx_inst_n62,
         prince_inst_sbox_inst8_yxxx_inst_n61,
         prince_inst_sbox_inst8_yxxx_inst_n60,
         prince_inst_sbox_inst8_yxxx_inst_n59,
         prince_inst_sbox_inst8_yxxx_inst_n58,
         prince_inst_sbox_inst8_yxxx_inst_n57,
         prince_inst_sbox_inst8_yxxx_inst_n56,
         prince_inst_sbox_inst8_yxxx_inst_n55,
         prince_inst_sbox_inst8_yxxx_inst_n54,
         prince_inst_sbox_inst8_yxxx_inst_n53,
         prince_inst_sbox_inst8_yxxx_inst_n52,
         prince_inst_sbox_inst8_yxxx_inst_n51,
         prince_inst_sbox_inst8_yxxx_inst_n50,
         prince_inst_sbox_inst8_yxxx_inst_n49,
         prince_inst_sbox_inst8_yxxx_inst_n48,
         prince_inst_sbox_inst8_yxxx_inst_n47,
         prince_inst_sbox_inst8_yxxx_inst_n46,
         prince_inst_sbox_inst8_yxxx_inst_n45,
         prince_inst_sbox_inst8_yxyy_inst_n68,
         prince_inst_sbox_inst8_yxyy_inst_n67,
         prince_inst_sbox_inst8_yxyy_inst_n66,
         prince_inst_sbox_inst8_yxyy_inst_n65,
         prince_inst_sbox_inst8_yxyy_inst_n64,
         prince_inst_sbox_inst8_yxyy_inst_n63,
         prince_inst_sbox_inst8_yxyy_inst_n62,
         prince_inst_sbox_inst8_yxyy_inst_n61,
         prince_inst_sbox_inst8_yxyy_inst_n60,
         prince_inst_sbox_inst8_yxyy_inst_n59,
         prince_inst_sbox_inst8_yxyy_inst_n58,
         prince_inst_sbox_inst8_yxyy_inst_n57,
         prince_inst_sbox_inst8_yxyy_inst_n56,
         prince_inst_sbox_inst8_yxyy_inst_n55,
         prince_inst_sbox_inst8_yxyy_inst_n54,
         prince_inst_sbox_inst8_yxyy_inst_n53,
         prince_inst_sbox_inst8_yxyy_inst_n52,
         prince_inst_sbox_inst8_yxyy_inst_n51,
         prince_inst_sbox_inst8_yxyy_inst_n50,
         prince_inst_sbox_inst8_yxyy_inst_n49,
         prince_inst_sbox_inst8_yyxy_inst_n75,
         prince_inst_sbox_inst8_yyxy_inst_n74,
         prince_inst_sbox_inst8_yyxy_inst_n73,
         prince_inst_sbox_inst8_yyxy_inst_n72,
         prince_inst_sbox_inst8_yyxy_inst_n71,
         prince_inst_sbox_inst8_yyxy_inst_n70,
         prince_inst_sbox_inst8_yyxy_inst_n69,
         prince_inst_sbox_inst8_yyxy_inst_n68,
         prince_inst_sbox_inst8_yyxy_inst_n67,
         prince_inst_sbox_inst8_yyxy_inst_n66,
         prince_inst_sbox_inst8_yyxy_inst_n65,
         prince_inst_sbox_inst8_yyxy_inst_n64,
         prince_inst_sbox_inst8_yyxy_inst_n63,
         prince_inst_sbox_inst8_yyxy_inst_n62,
         prince_inst_sbox_inst8_yyxy_inst_n61,
         prince_inst_sbox_inst8_yyxy_inst_n60,
         prince_inst_sbox_inst8_yyxy_inst_n59,
         prince_inst_sbox_inst8_yyxy_inst_n58,
         prince_inst_sbox_inst8_yyxy_inst_n57,
         prince_inst_sbox_inst8_yyxy_inst_n56,
         prince_inst_sbox_inst8_yyxy_inst_n55,
         prince_inst_sbox_inst8_yyxy_inst_n54,
         prince_inst_sbox_inst8_yyxy_inst_n53,
         prince_inst_sbox_inst8_yyyx_inst_n58,
         prince_inst_sbox_inst8_yyyx_inst_n57,
         prince_inst_sbox_inst8_yyyx_inst_n56,
         prince_inst_sbox_inst8_yyyx_inst_n55,
         prince_inst_sbox_inst8_yyyx_inst_n54,
         prince_inst_sbox_inst8_yyyx_inst_n53,
         prince_inst_sbox_inst8_yyyx_inst_n52,
         prince_inst_sbox_inst8_yyyx_inst_n51,
         prince_inst_sbox_inst8_yyyx_inst_n50,
         prince_inst_sbox_inst8_yyyx_inst_n49,
         prince_inst_sbox_inst8_yyyx_inst_n48,
         prince_inst_sbox_inst8_yyyx_inst_n47,
         prince_inst_sbox_inst8_yyyx_inst_n46,
         prince_inst_sbox_inst8_yyyx_inst_n45,
         prince_inst_sbox_inst8_yyyx_inst_n44,
         prince_inst_sbox_inst8_yyyx_inst_n43,
         prince_inst_sbox_inst8_yyyx_inst_n42,
         prince_inst_sbox_inst8_c_inst0_msk0_xr,
         prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_msk1_xr,
         prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_msk2_xr,
         prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_msk3_xr,
         prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_msk4_xr,
         prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_msk5_xr,
         prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_msk6_xr,
         prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_msk7_xr,
         prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst0_ax_n6,
         prince_inst_sbox_inst8_c_inst0_ax_n5,
         prince_inst_sbox_inst8_c_inst0_ay_n6,
         prince_inst_sbox_inst8_c_inst0_ay_n5,
         prince_inst_sbox_inst8_c_inst1_msk0_xr,
         prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_msk1_xr,
         prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_msk2_xr,
         prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_msk3_xr,
         prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_msk4_xr,
         prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_msk5_xr,
         prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_msk6_xr,
         prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_msk7_xr,
         prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst1_ax_n6,
         prince_inst_sbox_inst8_c_inst1_ax_n5,
         prince_inst_sbox_inst8_c_inst1_ay_n6,
         prince_inst_sbox_inst8_c_inst1_ay_n5,
         prince_inst_sbox_inst8_c_inst2_msk0_xr,
         prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_msk1_xr,
         prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_msk2_xr,
         prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_msk3_xr,
         prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_msk4_xr,
         prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_msk5_xr,
         prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_msk6_xr,
         prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_msk7_xr,
         prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst2_ax_n6,
         prince_inst_sbox_inst8_c_inst2_ax_n5,
         prince_inst_sbox_inst8_c_inst2_ay_n6,
         prince_inst_sbox_inst8_c_inst2_ay_n5,
         prince_inst_sbox_inst8_c_inst3_msk0_xr,
         prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_msk1_xr,
         prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_msk2_xr,
         prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_msk3_xr,
         prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_msk4_xr,
         prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_msk5_xr,
         prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_msk6_xr,
         prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_msk7_xr,
         prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst8_c_inst3_ax_n6,
         prince_inst_sbox_inst8_c_inst3_ax_n5,
         prince_inst_sbox_inst8_c_inst3_ay_n6,
         prince_inst_sbox_inst8_c_inst3_ay_n5, prince_inst_sbox_inst9_n10,
         prince_inst_sbox_inst9_n9, prince_inst_sbox_inst9_n8,
         prince_inst_sbox_inst9_n7, prince_inst_sbox_inst9_n6,
         prince_inst_sbox_inst9_xxxy_inst_n69,
         prince_inst_sbox_inst9_xxxy_inst_n68,
         prince_inst_sbox_inst9_xxxy_inst_n67,
         prince_inst_sbox_inst9_xxxy_inst_n66,
         prince_inst_sbox_inst9_xxxy_inst_n65,
         prince_inst_sbox_inst9_xxxy_inst_n64,
         prince_inst_sbox_inst9_xxxy_inst_n63,
         prince_inst_sbox_inst9_xxxy_inst_n62,
         prince_inst_sbox_inst9_xxxy_inst_n61,
         prince_inst_sbox_inst9_xxxy_inst_n60,
         prince_inst_sbox_inst9_xxxy_inst_n59,
         prince_inst_sbox_inst9_xxxy_inst_n58,
         prince_inst_sbox_inst9_xxxy_inst_n57,
         prince_inst_sbox_inst9_xxxy_inst_n56,
         prince_inst_sbox_inst9_xxxy_inst_n55,
         prince_inst_sbox_inst9_xxxy_inst_n54,
         prince_inst_sbox_inst9_xxxy_inst_n53,
         prince_inst_sbox_inst9_xxxy_inst_n52,
         prince_inst_sbox_inst9_xxxy_inst_n51,
         prince_inst_sbox_inst9_xxyx_inst_n55,
         prince_inst_sbox_inst9_xxyx_inst_n54,
         prince_inst_sbox_inst9_xxyx_inst_n53,
         prince_inst_sbox_inst9_xxyx_inst_n52,
         prince_inst_sbox_inst9_xxyx_inst_n51,
         prince_inst_sbox_inst9_xxyx_inst_n50,
         prince_inst_sbox_inst9_xxyx_inst_n49,
         prince_inst_sbox_inst9_xxyx_inst_n48,
         prince_inst_sbox_inst9_xxyx_inst_n47,
         prince_inst_sbox_inst9_xxyx_inst_n46,
         prince_inst_sbox_inst9_xxyx_inst_n45,
         prince_inst_sbox_inst9_xxyx_inst_n44,
         prince_inst_sbox_inst9_xxyx_inst_n43,
         prince_inst_sbox_inst9_xxyx_inst_n42,
         prince_inst_sbox_inst9_xxyx_inst_n41,
         prince_inst_sbox_inst9_xxyx_inst_n40,
         prince_inst_sbox_inst9_xxyx_inst_n39,
         prince_inst_sbox_inst9_xxyx_inst_n38,
         prince_inst_sbox_inst9_xyxx_inst_n74,
         prince_inst_sbox_inst9_xyxx_inst_n73,
         prince_inst_sbox_inst9_xyxx_inst_n72,
         prince_inst_sbox_inst9_xyxx_inst_n71,
         prince_inst_sbox_inst9_xyxx_inst_n70,
         prince_inst_sbox_inst9_xyxx_inst_n69,
         prince_inst_sbox_inst9_xyxx_inst_n68,
         prince_inst_sbox_inst9_xyxx_inst_n67,
         prince_inst_sbox_inst9_xyxx_inst_n66,
         prince_inst_sbox_inst9_xyxx_inst_n65,
         prince_inst_sbox_inst9_xyxx_inst_n64,
         prince_inst_sbox_inst9_xyxx_inst_n63,
         prince_inst_sbox_inst9_xyxx_inst_n62,
         prince_inst_sbox_inst9_xyxx_inst_n61,
         prince_inst_sbox_inst9_xyxx_inst_n60,
         prince_inst_sbox_inst9_xyxx_inst_n59,
         prince_inst_sbox_inst9_xyxx_inst_n58,
         prince_inst_sbox_inst9_xyxx_inst_n57,
         prince_inst_sbox_inst9_xyxx_inst_n56,
         prince_inst_sbox_inst9_xyxx_inst_n55,
         prince_inst_sbox_inst9_xyxx_inst_n54,
         prince_inst_sbox_inst9_xyxx_inst_n53,
         prince_inst_sbox_inst9_xyyy_inst_n61,
         prince_inst_sbox_inst9_xyyy_inst_n60,
         prince_inst_sbox_inst9_xyyy_inst_n59,
         prince_inst_sbox_inst9_xyyy_inst_n58,
         prince_inst_sbox_inst9_xyyy_inst_n57,
         prince_inst_sbox_inst9_xyyy_inst_n56,
         prince_inst_sbox_inst9_xyyy_inst_n55,
         prince_inst_sbox_inst9_xyyy_inst_n54,
         prince_inst_sbox_inst9_xyyy_inst_n53,
         prince_inst_sbox_inst9_xyyy_inst_n52,
         prince_inst_sbox_inst9_xyyy_inst_n51,
         prince_inst_sbox_inst9_xyyy_inst_n50,
         prince_inst_sbox_inst9_xyyy_inst_n49,
         prince_inst_sbox_inst9_xyyy_inst_n48,
         prince_inst_sbox_inst9_xyyy_inst_n47,
         prince_inst_sbox_inst9_xyyy_inst_n46,
         prince_inst_sbox_inst9_xyyy_inst_n45,
         prince_inst_sbox_inst9_xyyy_inst_n44,
         prince_inst_sbox_inst9_xyyy_inst_n43,
         prince_inst_sbox_inst9_xyyy_inst_n42,
         prince_inst_sbox_inst9_yxxx_inst_n64,
         prince_inst_sbox_inst9_yxxx_inst_n63,
         prince_inst_sbox_inst9_yxxx_inst_n62,
         prince_inst_sbox_inst9_yxxx_inst_n61,
         prince_inst_sbox_inst9_yxxx_inst_n60,
         prince_inst_sbox_inst9_yxxx_inst_n59,
         prince_inst_sbox_inst9_yxxx_inst_n58,
         prince_inst_sbox_inst9_yxxx_inst_n57,
         prince_inst_sbox_inst9_yxxx_inst_n56,
         prince_inst_sbox_inst9_yxxx_inst_n55,
         prince_inst_sbox_inst9_yxxx_inst_n54,
         prince_inst_sbox_inst9_yxxx_inst_n53,
         prince_inst_sbox_inst9_yxxx_inst_n52,
         prince_inst_sbox_inst9_yxxx_inst_n51,
         prince_inst_sbox_inst9_yxxx_inst_n50,
         prince_inst_sbox_inst9_yxxx_inst_n49,
         prince_inst_sbox_inst9_yxxx_inst_n48,
         prince_inst_sbox_inst9_yxxx_inst_n47,
         prince_inst_sbox_inst9_yxxx_inst_n46,
         prince_inst_sbox_inst9_yxxx_inst_n45,
         prince_inst_sbox_inst9_yxyy_inst_n68,
         prince_inst_sbox_inst9_yxyy_inst_n67,
         prince_inst_sbox_inst9_yxyy_inst_n66,
         prince_inst_sbox_inst9_yxyy_inst_n65,
         prince_inst_sbox_inst9_yxyy_inst_n64,
         prince_inst_sbox_inst9_yxyy_inst_n63,
         prince_inst_sbox_inst9_yxyy_inst_n62,
         prince_inst_sbox_inst9_yxyy_inst_n61,
         prince_inst_sbox_inst9_yxyy_inst_n60,
         prince_inst_sbox_inst9_yxyy_inst_n59,
         prince_inst_sbox_inst9_yxyy_inst_n58,
         prince_inst_sbox_inst9_yxyy_inst_n57,
         prince_inst_sbox_inst9_yxyy_inst_n56,
         prince_inst_sbox_inst9_yxyy_inst_n55,
         prince_inst_sbox_inst9_yxyy_inst_n54,
         prince_inst_sbox_inst9_yxyy_inst_n53,
         prince_inst_sbox_inst9_yxyy_inst_n52,
         prince_inst_sbox_inst9_yxyy_inst_n51,
         prince_inst_sbox_inst9_yxyy_inst_n50,
         prince_inst_sbox_inst9_yxyy_inst_n49,
         prince_inst_sbox_inst9_yyxy_inst_n75,
         prince_inst_sbox_inst9_yyxy_inst_n74,
         prince_inst_sbox_inst9_yyxy_inst_n73,
         prince_inst_sbox_inst9_yyxy_inst_n72,
         prince_inst_sbox_inst9_yyxy_inst_n71,
         prince_inst_sbox_inst9_yyxy_inst_n70,
         prince_inst_sbox_inst9_yyxy_inst_n69,
         prince_inst_sbox_inst9_yyxy_inst_n68,
         prince_inst_sbox_inst9_yyxy_inst_n67,
         prince_inst_sbox_inst9_yyxy_inst_n66,
         prince_inst_sbox_inst9_yyxy_inst_n65,
         prince_inst_sbox_inst9_yyxy_inst_n64,
         prince_inst_sbox_inst9_yyxy_inst_n63,
         prince_inst_sbox_inst9_yyxy_inst_n62,
         prince_inst_sbox_inst9_yyxy_inst_n61,
         prince_inst_sbox_inst9_yyxy_inst_n60,
         prince_inst_sbox_inst9_yyxy_inst_n59,
         prince_inst_sbox_inst9_yyxy_inst_n58,
         prince_inst_sbox_inst9_yyxy_inst_n57,
         prince_inst_sbox_inst9_yyxy_inst_n56,
         prince_inst_sbox_inst9_yyxy_inst_n55,
         prince_inst_sbox_inst9_yyxy_inst_n54,
         prince_inst_sbox_inst9_yyxy_inst_n53,
         prince_inst_sbox_inst9_yyyx_inst_n58,
         prince_inst_sbox_inst9_yyyx_inst_n57,
         prince_inst_sbox_inst9_yyyx_inst_n56,
         prince_inst_sbox_inst9_yyyx_inst_n55,
         prince_inst_sbox_inst9_yyyx_inst_n54,
         prince_inst_sbox_inst9_yyyx_inst_n53,
         prince_inst_sbox_inst9_yyyx_inst_n52,
         prince_inst_sbox_inst9_yyyx_inst_n51,
         prince_inst_sbox_inst9_yyyx_inst_n50,
         prince_inst_sbox_inst9_yyyx_inst_n49,
         prince_inst_sbox_inst9_yyyx_inst_n48,
         prince_inst_sbox_inst9_yyyx_inst_n47,
         prince_inst_sbox_inst9_yyyx_inst_n46,
         prince_inst_sbox_inst9_yyyx_inst_n45,
         prince_inst_sbox_inst9_yyyx_inst_n44,
         prince_inst_sbox_inst9_yyyx_inst_n43,
         prince_inst_sbox_inst9_yyyx_inst_n42,
         prince_inst_sbox_inst9_c_inst0_msk0_xr,
         prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_msk1_xr,
         prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_msk2_xr,
         prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_msk3_xr,
         prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_msk4_xr,
         prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_msk5_xr,
         prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_msk6_xr,
         prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_msk7_xr,
         prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst0_ax_n6,
         prince_inst_sbox_inst9_c_inst0_ax_n5,
         prince_inst_sbox_inst9_c_inst0_ay_n6,
         prince_inst_sbox_inst9_c_inst0_ay_n5,
         prince_inst_sbox_inst9_c_inst1_msk0_xr,
         prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_msk1_xr,
         prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_msk2_xr,
         prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_msk3_xr,
         prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_msk4_xr,
         prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_msk5_xr,
         prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_msk6_xr,
         prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_msk7_xr,
         prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst1_ax_n6,
         prince_inst_sbox_inst9_c_inst1_ax_n5,
         prince_inst_sbox_inst9_c_inst1_ay_n6,
         prince_inst_sbox_inst9_c_inst1_ay_n5,
         prince_inst_sbox_inst9_c_inst2_msk0_xr,
         prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_msk1_xr,
         prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_msk2_xr,
         prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_msk3_xr,
         prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_msk4_xr,
         prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_msk5_xr,
         prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_msk6_xr,
         prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_msk7_xr,
         prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst2_ax_n6,
         prince_inst_sbox_inst9_c_inst2_ax_n5,
         prince_inst_sbox_inst9_c_inst2_ay_n6,
         prince_inst_sbox_inst9_c_inst2_ay_n5,
         prince_inst_sbox_inst9_c_inst3_msk0_xr,
         prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_msk1_xr,
         prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_msk2_xr,
         prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_msk3_xr,
         prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_msk4_xr,
         prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_msk5_xr,
         prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_msk6_xr,
         prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_msk7_xr,
         prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst9_c_inst3_ax_n6,
         prince_inst_sbox_inst9_c_inst3_ax_n5,
         prince_inst_sbox_inst9_c_inst3_ay_n6,
         prince_inst_sbox_inst9_c_inst3_ay_n5, prince_inst_sbox_inst10_n11,
         prince_inst_sbox_inst10_n10, prince_inst_sbox_inst10_n9,
         prince_inst_sbox_inst10_n8, prince_inst_sbox_inst10_n7,
         prince_inst_sbox_inst10_xxxy_inst_n69,
         prince_inst_sbox_inst10_xxxy_inst_n68,
         prince_inst_sbox_inst10_xxxy_inst_n67,
         prince_inst_sbox_inst10_xxxy_inst_n66,
         prince_inst_sbox_inst10_xxxy_inst_n65,
         prince_inst_sbox_inst10_xxxy_inst_n64,
         prince_inst_sbox_inst10_xxxy_inst_n63,
         prince_inst_sbox_inst10_xxxy_inst_n62,
         prince_inst_sbox_inst10_xxxy_inst_n61,
         prince_inst_sbox_inst10_xxxy_inst_n60,
         prince_inst_sbox_inst10_xxxy_inst_n59,
         prince_inst_sbox_inst10_xxxy_inst_n58,
         prince_inst_sbox_inst10_xxxy_inst_n57,
         prince_inst_sbox_inst10_xxxy_inst_n56,
         prince_inst_sbox_inst10_xxxy_inst_n55,
         prince_inst_sbox_inst10_xxxy_inst_n54,
         prince_inst_sbox_inst10_xxxy_inst_n53,
         prince_inst_sbox_inst10_xxxy_inst_n52,
         prince_inst_sbox_inst10_xxxy_inst_n51,
         prince_inst_sbox_inst10_xxyx_inst_n55,
         prince_inst_sbox_inst10_xxyx_inst_n54,
         prince_inst_sbox_inst10_xxyx_inst_n53,
         prince_inst_sbox_inst10_xxyx_inst_n52,
         prince_inst_sbox_inst10_xxyx_inst_n51,
         prince_inst_sbox_inst10_xxyx_inst_n50,
         prince_inst_sbox_inst10_xxyx_inst_n49,
         prince_inst_sbox_inst10_xxyx_inst_n48,
         prince_inst_sbox_inst10_xxyx_inst_n47,
         prince_inst_sbox_inst10_xxyx_inst_n46,
         prince_inst_sbox_inst10_xxyx_inst_n45,
         prince_inst_sbox_inst10_xxyx_inst_n44,
         prince_inst_sbox_inst10_xxyx_inst_n43,
         prince_inst_sbox_inst10_xxyx_inst_n42,
         prince_inst_sbox_inst10_xxyx_inst_n41,
         prince_inst_sbox_inst10_xxyx_inst_n40,
         prince_inst_sbox_inst10_xxyx_inst_n39,
         prince_inst_sbox_inst10_xxyx_inst_n38,
         prince_inst_sbox_inst10_xyxx_inst_n74,
         prince_inst_sbox_inst10_xyxx_inst_n73,
         prince_inst_sbox_inst10_xyxx_inst_n72,
         prince_inst_sbox_inst10_xyxx_inst_n71,
         prince_inst_sbox_inst10_xyxx_inst_n70,
         prince_inst_sbox_inst10_xyxx_inst_n69,
         prince_inst_sbox_inst10_xyxx_inst_n68,
         prince_inst_sbox_inst10_xyxx_inst_n67,
         prince_inst_sbox_inst10_xyxx_inst_n66,
         prince_inst_sbox_inst10_xyxx_inst_n65,
         prince_inst_sbox_inst10_xyxx_inst_n64,
         prince_inst_sbox_inst10_xyxx_inst_n63,
         prince_inst_sbox_inst10_xyxx_inst_n62,
         prince_inst_sbox_inst10_xyxx_inst_n61,
         prince_inst_sbox_inst10_xyxx_inst_n60,
         prince_inst_sbox_inst10_xyxx_inst_n59,
         prince_inst_sbox_inst10_xyxx_inst_n58,
         prince_inst_sbox_inst10_xyxx_inst_n57,
         prince_inst_sbox_inst10_xyxx_inst_n56,
         prince_inst_sbox_inst10_xyxx_inst_n55,
         prince_inst_sbox_inst10_xyxx_inst_n54,
         prince_inst_sbox_inst10_xyxx_inst_n53,
         prince_inst_sbox_inst10_xyyy_inst_n61,
         prince_inst_sbox_inst10_xyyy_inst_n60,
         prince_inst_sbox_inst10_xyyy_inst_n59,
         prince_inst_sbox_inst10_xyyy_inst_n58,
         prince_inst_sbox_inst10_xyyy_inst_n57,
         prince_inst_sbox_inst10_xyyy_inst_n56,
         prince_inst_sbox_inst10_xyyy_inst_n55,
         prince_inst_sbox_inst10_xyyy_inst_n54,
         prince_inst_sbox_inst10_xyyy_inst_n53,
         prince_inst_sbox_inst10_xyyy_inst_n52,
         prince_inst_sbox_inst10_xyyy_inst_n51,
         prince_inst_sbox_inst10_xyyy_inst_n50,
         prince_inst_sbox_inst10_xyyy_inst_n49,
         prince_inst_sbox_inst10_xyyy_inst_n48,
         prince_inst_sbox_inst10_xyyy_inst_n47,
         prince_inst_sbox_inst10_xyyy_inst_n46,
         prince_inst_sbox_inst10_xyyy_inst_n45,
         prince_inst_sbox_inst10_xyyy_inst_n44,
         prince_inst_sbox_inst10_xyyy_inst_n43,
         prince_inst_sbox_inst10_xyyy_inst_n42,
         prince_inst_sbox_inst10_yxxx_inst_n64,
         prince_inst_sbox_inst10_yxxx_inst_n63,
         prince_inst_sbox_inst10_yxxx_inst_n62,
         prince_inst_sbox_inst10_yxxx_inst_n61,
         prince_inst_sbox_inst10_yxxx_inst_n60,
         prince_inst_sbox_inst10_yxxx_inst_n59,
         prince_inst_sbox_inst10_yxxx_inst_n58,
         prince_inst_sbox_inst10_yxxx_inst_n57,
         prince_inst_sbox_inst10_yxxx_inst_n56,
         prince_inst_sbox_inst10_yxxx_inst_n55,
         prince_inst_sbox_inst10_yxxx_inst_n54,
         prince_inst_sbox_inst10_yxxx_inst_n53,
         prince_inst_sbox_inst10_yxxx_inst_n52,
         prince_inst_sbox_inst10_yxxx_inst_n51,
         prince_inst_sbox_inst10_yxxx_inst_n50,
         prince_inst_sbox_inst10_yxxx_inst_n49,
         prince_inst_sbox_inst10_yxxx_inst_n48,
         prince_inst_sbox_inst10_yxxx_inst_n47,
         prince_inst_sbox_inst10_yxxx_inst_n46,
         prince_inst_sbox_inst10_yxxx_inst_n45,
         prince_inst_sbox_inst10_yxyy_inst_n68,
         prince_inst_sbox_inst10_yxyy_inst_n67,
         prince_inst_sbox_inst10_yxyy_inst_n66,
         prince_inst_sbox_inst10_yxyy_inst_n65,
         prince_inst_sbox_inst10_yxyy_inst_n64,
         prince_inst_sbox_inst10_yxyy_inst_n63,
         prince_inst_sbox_inst10_yxyy_inst_n62,
         prince_inst_sbox_inst10_yxyy_inst_n61,
         prince_inst_sbox_inst10_yxyy_inst_n60,
         prince_inst_sbox_inst10_yxyy_inst_n59,
         prince_inst_sbox_inst10_yxyy_inst_n58,
         prince_inst_sbox_inst10_yxyy_inst_n57,
         prince_inst_sbox_inst10_yxyy_inst_n56,
         prince_inst_sbox_inst10_yxyy_inst_n55,
         prince_inst_sbox_inst10_yxyy_inst_n54,
         prince_inst_sbox_inst10_yxyy_inst_n53,
         prince_inst_sbox_inst10_yxyy_inst_n52,
         prince_inst_sbox_inst10_yxyy_inst_n51,
         prince_inst_sbox_inst10_yxyy_inst_n50,
         prince_inst_sbox_inst10_yxyy_inst_n49,
         prince_inst_sbox_inst10_yyxy_inst_n75,
         prince_inst_sbox_inst10_yyxy_inst_n74,
         prince_inst_sbox_inst10_yyxy_inst_n73,
         prince_inst_sbox_inst10_yyxy_inst_n72,
         prince_inst_sbox_inst10_yyxy_inst_n71,
         prince_inst_sbox_inst10_yyxy_inst_n70,
         prince_inst_sbox_inst10_yyxy_inst_n69,
         prince_inst_sbox_inst10_yyxy_inst_n68,
         prince_inst_sbox_inst10_yyxy_inst_n67,
         prince_inst_sbox_inst10_yyxy_inst_n66,
         prince_inst_sbox_inst10_yyxy_inst_n65,
         prince_inst_sbox_inst10_yyxy_inst_n64,
         prince_inst_sbox_inst10_yyxy_inst_n63,
         prince_inst_sbox_inst10_yyxy_inst_n62,
         prince_inst_sbox_inst10_yyxy_inst_n61,
         prince_inst_sbox_inst10_yyxy_inst_n60,
         prince_inst_sbox_inst10_yyxy_inst_n59,
         prince_inst_sbox_inst10_yyxy_inst_n58,
         prince_inst_sbox_inst10_yyxy_inst_n57,
         prince_inst_sbox_inst10_yyxy_inst_n56,
         prince_inst_sbox_inst10_yyxy_inst_n55,
         prince_inst_sbox_inst10_yyxy_inst_n54,
         prince_inst_sbox_inst10_yyxy_inst_n53,
         prince_inst_sbox_inst10_yyyx_inst_n58,
         prince_inst_sbox_inst10_yyyx_inst_n57,
         prince_inst_sbox_inst10_yyyx_inst_n56,
         prince_inst_sbox_inst10_yyyx_inst_n55,
         prince_inst_sbox_inst10_yyyx_inst_n54,
         prince_inst_sbox_inst10_yyyx_inst_n53,
         prince_inst_sbox_inst10_yyyx_inst_n52,
         prince_inst_sbox_inst10_yyyx_inst_n51,
         prince_inst_sbox_inst10_yyyx_inst_n50,
         prince_inst_sbox_inst10_yyyx_inst_n49,
         prince_inst_sbox_inst10_yyyx_inst_n48,
         prince_inst_sbox_inst10_yyyx_inst_n47,
         prince_inst_sbox_inst10_yyyx_inst_n46,
         prince_inst_sbox_inst10_yyyx_inst_n45,
         prince_inst_sbox_inst10_yyyx_inst_n44,
         prince_inst_sbox_inst10_yyyx_inst_n43,
         prince_inst_sbox_inst10_yyyx_inst_n42,
         prince_inst_sbox_inst10_c_inst0_msk0_xr,
         prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_msk1_xr,
         prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_msk2_xr,
         prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_msk3_xr,
         prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_msk4_xr,
         prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_msk5_xr,
         prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_msk6_xr,
         prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_msk7_xr,
         prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst0_ax_n6,
         prince_inst_sbox_inst10_c_inst0_ax_n5,
         prince_inst_sbox_inst10_c_inst0_ay_n6,
         prince_inst_sbox_inst10_c_inst0_ay_n5,
         prince_inst_sbox_inst10_c_inst1_msk0_xr,
         prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_msk1_xr,
         prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_msk2_xr,
         prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_msk3_xr,
         prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_msk4_xr,
         prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_msk5_xr,
         prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_msk6_xr,
         prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_msk7_xr,
         prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst1_ax_n6,
         prince_inst_sbox_inst10_c_inst1_ax_n5,
         prince_inst_sbox_inst10_c_inst1_ay_n6,
         prince_inst_sbox_inst10_c_inst1_ay_n5,
         prince_inst_sbox_inst10_c_inst2_msk0_xr,
         prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_msk1_xr,
         prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_msk2_xr,
         prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_msk3_xr,
         prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_msk4_xr,
         prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_msk5_xr,
         prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_msk6_xr,
         prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_msk7_xr,
         prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst2_ax_n6,
         prince_inst_sbox_inst10_c_inst2_ax_n5,
         prince_inst_sbox_inst10_c_inst2_ay_n6,
         prince_inst_sbox_inst10_c_inst2_ay_n5,
         prince_inst_sbox_inst10_c_inst3_msk0_xr,
         prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_msk1_xr,
         prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_msk2_xr,
         prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_msk3_xr,
         prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_msk4_xr,
         prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_msk5_xr,
         prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_msk6_xr,
         prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_msk7_xr,
         prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst10_c_inst3_ax_n6,
         prince_inst_sbox_inst10_c_inst3_ax_n5,
         prince_inst_sbox_inst10_c_inst3_ay_n6,
         prince_inst_sbox_inst10_c_inst3_ay_n5, prince_inst_sbox_inst11_n13,
         prince_inst_sbox_inst11_n12, prince_inst_sbox_inst11_n11,
         prince_inst_sbox_inst11_n10, prince_inst_sbox_inst11_n9,
         prince_inst_sbox_inst11_n8, prince_inst_sbox_inst11_n7,
         prince_inst_sbox_inst11_xxxy_inst_n69,
         prince_inst_sbox_inst11_xxxy_inst_n68,
         prince_inst_sbox_inst11_xxxy_inst_n67,
         prince_inst_sbox_inst11_xxxy_inst_n66,
         prince_inst_sbox_inst11_xxxy_inst_n65,
         prince_inst_sbox_inst11_xxxy_inst_n64,
         prince_inst_sbox_inst11_xxxy_inst_n63,
         prince_inst_sbox_inst11_xxxy_inst_n62,
         prince_inst_sbox_inst11_xxxy_inst_n61,
         prince_inst_sbox_inst11_xxxy_inst_n60,
         prince_inst_sbox_inst11_xxxy_inst_n59,
         prince_inst_sbox_inst11_xxxy_inst_n58,
         prince_inst_sbox_inst11_xxxy_inst_n57,
         prince_inst_sbox_inst11_xxxy_inst_n56,
         prince_inst_sbox_inst11_xxxy_inst_n55,
         prince_inst_sbox_inst11_xxxy_inst_n54,
         prince_inst_sbox_inst11_xxxy_inst_n53,
         prince_inst_sbox_inst11_xxxy_inst_n52,
         prince_inst_sbox_inst11_xxxy_inst_n51,
         prince_inst_sbox_inst11_xxyx_inst_n55,
         prince_inst_sbox_inst11_xxyx_inst_n54,
         prince_inst_sbox_inst11_xxyx_inst_n53,
         prince_inst_sbox_inst11_xxyx_inst_n52,
         prince_inst_sbox_inst11_xxyx_inst_n51,
         prince_inst_sbox_inst11_xxyx_inst_n50,
         prince_inst_sbox_inst11_xxyx_inst_n49,
         prince_inst_sbox_inst11_xxyx_inst_n48,
         prince_inst_sbox_inst11_xxyx_inst_n47,
         prince_inst_sbox_inst11_xxyx_inst_n46,
         prince_inst_sbox_inst11_xxyx_inst_n45,
         prince_inst_sbox_inst11_xxyx_inst_n44,
         prince_inst_sbox_inst11_xxyx_inst_n43,
         prince_inst_sbox_inst11_xxyx_inst_n42,
         prince_inst_sbox_inst11_xxyx_inst_n41,
         prince_inst_sbox_inst11_xxyx_inst_n40,
         prince_inst_sbox_inst11_xxyx_inst_n39,
         prince_inst_sbox_inst11_xxyx_inst_n38,
         prince_inst_sbox_inst11_xyxx_inst_n74,
         prince_inst_sbox_inst11_xyxx_inst_n73,
         prince_inst_sbox_inst11_xyxx_inst_n72,
         prince_inst_sbox_inst11_xyxx_inst_n71,
         prince_inst_sbox_inst11_xyxx_inst_n70,
         prince_inst_sbox_inst11_xyxx_inst_n69,
         prince_inst_sbox_inst11_xyxx_inst_n68,
         prince_inst_sbox_inst11_xyxx_inst_n67,
         prince_inst_sbox_inst11_xyxx_inst_n66,
         prince_inst_sbox_inst11_xyxx_inst_n65,
         prince_inst_sbox_inst11_xyxx_inst_n64,
         prince_inst_sbox_inst11_xyxx_inst_n63,
         prince_inst_sbox_inst11_xyxx_inst_n62,
         prince_inst_sbox_inst11_xyxx_inst_n61,
         prince_inst_sbox_inst11_xyxx_inst_n60,
         prince_inst_sbox_inst11_xyxx_inst_n59,
         prince_inst_sbox_inst11_xyxx_inst_n58,
         prince_inst_sbox_inst11_xyxx_inst_n57,
         prince_inst_sbox_inst11_xyxx_inst_n56,
         prince_inst_sbox_inst11_xyxx_inst_n55,
         prince_inst_sbox_inst11_xyxx_inst_n54,
         prince_inst_sbox_inst11_xyxx_inst_n53,
         prince_inst_sbox_inst11_xyyy_inst_n61,
         prince_inst_sbox_inst11_xyyy_inst_n60,
         prince_inst_sbox_inst11_xyyy_inst_n59,
         prince_inst_sbox_inst11_xyyy_inst_n58,
         prince_inst_sbox_inst11_xyyy_inst_n57,
         prince_inst_sbox_inst11_xyyy_inst_n56,
         prince_inst_sbox_inst11_xyyy_inst_n55,
         prince_inst_sbox_inst11_xyyy_inst_n54,
         prince_inst_sbox_inst11_xyyy_inst_n53,
         prince_inst_sbox_inst11_xyyy_inst_n52,
         prince_inst_sbox_inst11_xyyy_inst_n51,
         prince_inst_sbox_inst11_xyyy_inst_n50,
         prince_inst_sbox_inst11_xyyy_inst_n49,
         prince_inst_sbox_inst11_xyyy_inst_n48,
         prince_inst_sbox_inst11_xyyy_inst_n47,
         prince_inst_sbox_inst11_xyyy_inst_n46,
         prince_inst_sbox_inst11_xyyy_inst_n45,
         prince_inst_sbox_inst11_xyyy_inst_n44,
         prince_inst_sbox_inst11_xyyy_inst_n43,
         prince_inst_sbox_inst11_xyyy_inst_n42,
         prince_inst_sbox_inst11_yxxx_inst_n64,
         prince_inst_sbox_inst11_yxxx_inst_n63,
         prince_inst_sbox_inst11_yxxx_inst_n62,
         prince_inst_sbox_inst11_yxxx_inst_n61,
         prince_inst_sbox_inst11_yxxx_inst_n60,
         prince_inst_sbox_inst11_yxxx_inst_n59,
         prince_inst_sbox_inst11_yxxx_inst_n58,
         prince_inst_sbox_inst11_yxxx_inst_n57,
         prince_inst_sbox_inst11_yxxx_inst_n56,
         prince_inst_sbox_inst11_yxxx_inst_n55,
         prince_inst_sbox_inst11_yxxx_inst_n54,
         prince_inst_sbox_inst11_yxxx_inst_n53,
         prince_inst_sbox_inst11_yxxx_inst_n52,
         prince_inst_sbox_inst11_yxxx_inst_n51,
         prince_inst_sbox_inst11_yxxx_inst_n50,
         prince_inst_sbox_inst11_yxxx_inst_n49,
         prince_inst_sbox_inst11_yxxx_inst_n48,
         prince_inst_sbox_inst11_yxxx_inst_n47,
         prince_inst_sbox_inst11_yxxx_inst_n46,
         prince_inst_sbox_inst11_yxxx_inst_n45,
         prince_inst_sbox_inst11_yxyy_inst_n68,
         prince_inst_sbox_inst11_yxyy_inst_n67,
         prince_inst_sbox_inst11_yxyy_inst_n66,
         prince_inst_sbox_inst11_yxyy_inst_n65,
         prince_inst_sbox_inst11_yxyy_inst_n64,
         prince_inst_sbox_inst11_yxyy_inst_n63,
         prince_inst_sbox_inst11_yxyy_inst_n62,
         prince_inst_sbox_inst11_yxyy_inst_n61,
         prince_inst_sbox_inst11_yxyy_inst_n60,
         prince_inst_sbox_inst11_yxyy_inst_n59,
         prince_inst_sbox_inst11_yxyy_inst_n58,
         prince_inst_sbox_inst11_yxyy_inst_n57,
         prince_inst_sbox_inst11_yxyy_inst_n56,
         prince_inst_sbox_inst11_yxyy_inst_n55,
         prince_inst_sbox_inst11_yxyy_inst_n54,
         prince_inst_sbox_inst11_yxyy_inst_n53,
         prince_inst_sbox_inst11_yxyy_inst_n52,
         prince_inst_sbox_inst11_yxyy_inst_n51,
         prince_inst_sbox_inst11_yxyy_inst_n50,
         prince_inst_sbox_inst11_yxyy_inst_n49,
         prince_inst_sbox_inst11_yyxy_inst_n75,
         prince_inst_sbox_inst11_yyxy_inst_n74,
         prince_inst_sbox_inst11_yyxy_inst_n73,
         prince_inst_sbox_inst11_yyxy_inst_n72,
         prince_inst_sbox_inst11_yyxy_inst_n71,
         prince_inst_sbox_inst11_yyxy_inst_n70,
         prince_inst_sbox_inst11_yyxy_inst_n69,
         prince_inst_sbox_inst11_yyxy_inst_n68,
         prince_inst_sbox_inst11_yyxy_inst_n67,
         prince_inst_sbox_inst11_yyxy_inst_n66,
         prince_inst_sbox_inst11_yyxy_inst_n65,
         prince_inst_sbox_inst11_yyxy_inst_n64,
         prince_inst_sbox_inst11_yyxy_inst_n63,
         prince_inst_sbox_inst11_yyxy_inst_n62,
         prince_inst_sbox_inst11_yyxy_inst_n61,
         prince_inst_sbox_inst11_yyxy_inst_n60,
         prince_inst_sbox_inst11_yyxy_inst_n59,
         prince_inst_sbox_inst11_yyxy_inst_n58,
         prince_inst_sbox_inst11_yyxy_inst_n57,
         prince_inst_sbox_inst11_yyxy_inst_n56,
         prince_inst_sbox_inst11_yyxy_inst_n55,
         prince_inst_sbox_inst11_yyxy_inst_n54,
         prince_inst_sbox_inst11_yyxy_inst_n53,
         prince_inst_sbox_inst11_yyyx_inst_n58,
         prince_inst_sbox_inst11_yyyx_inst_n57,
         prince_inst_sbox_inst11_yyyx_inst_n56,
         prince_inst_sbox_inst11_yyyx_inst_n55,
         prince_inst_sbox_inst11_yyyx_inst_n54,
         prince_inst_sbox_inst11_yyyx_inst_n53,
         prince_inst_sbox_inst11_yyyx_inst_n52,
         prince_inst_sbox_inst11_yyyx_inst_n51,
         prince_inst_sbox_inst11_yyyx_inst_n50,
         prince_inst_sbox_inst11_yyyx_inst_n49,
         prince_inst_sbox_inst11_yyyx_inst_n48,
         prince_inst_sbox_inst11_yyyx_inst_n47,
         prince_inst_sbox_inst11_yyyx_inst_n46,
         prince_inst_sbox_inst11_yyyx_inst_n45,
         prince_inst_sbox_inst11_yyyx_inst_n44,
         prince_inst_sbox_inst11_yyyx_inst_n43,
         prince_inst_sbox_inst11_yyyx_inst_n42,
         prince_inst_sbox_inst11_c_inst0_msk0_xr,
         prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_msk1_xr,
         prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_msk2_xr,
         prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_msk3_xr,
         prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_msk4_xr,
         prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_msk5_xr,
         prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_msk6_xr,
         prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_msk7_xr,
         prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst0_ax_n6,
         prince_inst_sbox_inst11_c_inst0_ax_n5,
         prince_inst_sbox_inst11_c_inst0_ay_n6,
         prince_inst_sbox_inst11_c_inst0_ay_n5,
         prince_inst_sbox_inst11_c_inst1_msk0_xr,
         prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_msk1_xr,
         prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_msk2_xr,
         prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_msk3_xr,
         prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_msk4_xr,
         prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_msk5_xr,
         prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_msk6_xr,
         prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_msk7_xr,
         prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst1_ax_n6,
         prince_inst_sbox_inst11_c_inst1_ax_n5,
         prince_inst_sbox_inst11_c_inst1_ay_n6,
         prince_inst_sbox_inst11_c_inst1_ay_n5,
         prince_inst_sbox_inst11_c_inst2_msk0_xr,
         prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_msk1_xr,
         prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_msk2_xr,
         prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_msk3_xr,
         prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_msk4_xr,
         prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_msk5_xr,
         prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_msk6_xr,
         prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_msk7_xr,
         prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst2_ax_n6,
         prince_inst_sbox_inst11_c_inst2_ax_n5,
         prince_inst_sbox_inst11_c_inst2_ay_n6,
         prince_inst_sbox_inst11_c_inst2_ay_n5,
         prince_inst_sbox_inst11_c_inst3_msk0_xr,
         prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_msk1_xr,
         prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_msk2_xr,
         prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_msk3_xr,
         prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_msk4_xr,
         prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_msk5_xr,
         prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_msk6_xr,
         prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_msk7_xr,
         prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst11_c_inst3_ax_n6,
         prince_inst_sbox_inst11_c_inst3_ax_n5,
         prince_inst_sbox_inst11_c_inst3_ay_n6,
         prince_inst_sbox_inst11_c_inst3_ay_n5, prince_inst_sbox_inst12_n13,
         prince_inst_sbox_inst12_n12, prince_inst_sbox_inst12_n11,
         prince_inst_sbox_inst12_n10, prince_inst_sbox_inst12_n9,
         prince_inst_sbox_inst12_n8, prince_inst_sbox_inst12_n7,
         prince_inst_sbox_inst12_xxxy_inst_n69,
         prince_inst_sbox_inst12_xxxy_inst_n68,
         prince_inst_sbox_inst12_xxxy_inst_n67,
         prince_inst_sbox_inst12_xxxy_inst_n66,
         prince_inst_sbox_inst12_xxxy_inst_n65,
         prince_inst_sbox_inst12_xxxy_inst_n64,
         prince_inst_sbox_inst12_xxxy_inst_n63,
         prince_inst_sbox_inst12_xxxy_inst_n62,
         prince_inst_sbox_inst12_xxxy_inst_n61,
         prince_inst_sbox_inst12_xxxy_inst_n60,
         prince_inst_sbox_inst12_xxxy_inst_n59,
         prince_inst_sbox_inst12_xxxy_inst_n58,
         prince_inst_sbox_inst12_xxxy_inst_n57,
         prince_inst_sbox_inst12_xxxy_inst_n56,
         prince_inst_sbox_inst12_xxxy_inst_n55,
         prince_inst_sbox_inst12_xxxy_inst_n54,
         prince_inst_sbox_inst12_xxxy_inst_n53,
         prince_inst_sbox_inst12_xxxy_inst_n52,
         prince_inst_sbox_inst12_xxxy_inst_n51,
         prince_inst_sbox_inst12_xxyx_inst_n55,
         prince_inst_sbox_inst12_xxyx_inst_n54,
         prince_inst_sbox_inst12_xxyx_inst_n53,
         prince_inst_sbox_inst12_xxyx_inst_n52,
         prince_inst_sbox_inst12_xxyx_inst_n51,
         prince_inst_sbox_inst12_xxyx_inst_n50,
         prince_inst_sbox_inst12_xxyx_inst_n49,
         prince_inst_sbox_inst12_xxyx_inst_n48,
         prince_inst_sbox_inst12_xxyx_inst_n47,
         prince_inst_sbox_inst12_xxyx_inst_n46,
         prince_inst_sbox_inst12_xxyx_inst_n45,
         prince_inst_sbox_inst12_xxyx_inst_n44,
         prince_inst_sbox_inst12_xxyx_inst_n43,
         prince_inst_sbox_inst12_xxyx_inst_n42,
         prince_inst_sbox_inst12_xxyx_inst_n41,
         prince_inst_sbox_inst12_xxyx_inst_n40,
         prince_inst_sbox_inst12_xxyx_inst_n39,
         prince_inst_sbox_inst12_xxyx_inst_n38,
         prince_inst_sbox_inst12_xyxx_inst_n74,
         prince_inst_sbox_inst12_xyxx_inst_n73,
         prince_inst_sbox_inst12_xyxx_inst_n72,
         prince_inst_sbox_inst12_xyxx_inst_n71,
         prince_inst_sbox_inst12_xyxx_inst_n70,
         prince_inst_sbox_inst12_xyxx_inst_n69,
         prince_inst_sbox_inst12_xyxx_inst_n68,
         prince_inst_sbox_inst12_xyxx_inst_n67,
         prince_inst_sbox_inst12_xyxx_inst_n66,
         prince_inst_sbox_inst12_xyxx_inst_n65,
         prince_inst_sbox_inst12_xyxx_inst_n64,
         prince_inst_sbox_inst12_xyxx_inst_n63,
         prince_inst_sbox_inst12_xyxx_inst_n62,
         prince_inst_sbox_inst12_xyxx_inst_n61,
         prince_inst_sbox_inst12_xyxx_inst_n60,
         prince_inst_sbox_inst12_xyxx_inst_n59,
         prince_inst_sbox_inst12_xyxx_inst_n58,
         prince_inst_sbox_inst12_xyxx_inst_n57,
         prince_inst_sbox_inst12_xyxx_inst_n56,
         prince_inst_sbox_inst12_xyxx_inst_n55,
         prince_inst_sbox_inst12_xyxx_inst_n54,
         prince_inst_sbox_inst12_xyxx_inst_n53,
         prince_inst_sbox_inst12_xyyy_inst_n61,
         prince_inst_sbox_inst12_xyyy_inst_n60,
         prince_inst_sbox_inst12_xyyy_inst_n59,
         prince_inst_sbox_inst12_xyyy_inst_n58,
         prince_inst_sbox_inst12_xyyy_inst_n57,
         prince_inst_sbox_inst12_xyyy_inst_n56,
         prince_inst_sbox_inst12_xyyy_inst_n55,
         prince_inst_sbox_inst12_xyyy_inst_n54,
         prince_inst_sbox_inst12_xyyy_inst_n53,
         prince_inst_sbox_inst12_xyyy_inst_n52,
         prince_inst_sbox_inst12_xyyy_inst_n51,
         prince_inst_sbox_inst12_xyyy_inst_n50,
         prince_inst_sbox_inst12_xyyy_inst_n49,
         prince_inst_sbox_inst12_xyyy_inst_n48,
         prince_inst_sbox_inst12_xyyy_inst_n47,
         prince_inst_sbox_inst12_xyyy_inst_n46,
         prince_inst_sbox_inst12_xyyy_inst_n45,
         prince_inst_sbox_inst12_xyyy_inst_n44,
         prince_inst_sbox_inst12_xyyy_inst_n43,
         prince_inst_sbox_inst12_xyyy_inst_n42,
         prince_inst_sbox_inst12_yxxx_inst_n64,
         prince_inst_sbox_inst12_yxxx_inst_n63,
         prince_inst_sbox_inst12_yxxx_inst_n62,
         prince_inst_sbox_inst12_yxxx_inst_n61,
         prince_inst_sbox_inst12_yxxx_inst_n60,
         prince_inst_sbox_inst12_yxxx_inst_n59,
         prince_inst_sbox_inst12_yxxx_inst_n58,
         prince_inst_sbox_inst12_yxxx_inst_n57,
         prince_inst_sbox_inst12_yxxx_inst_n56,
         prince_inst_sbox_inst12_yxxx_inst_n55,
         prince_inst_sbox_inst12_yxxx_inst_n54,
         prince_inst_sbox_inst12_yxxx_inst_n53,
         prince_inst_sbox_inst12_yxxx_inst_n52,
         prince_inst_sbox_inst12_yxxx_inst_n51,
         prince_inst_sbox_inst12_yxxx_inst_n50,
         prince_inst_sbox_inst12_yxxx_inst_n49,
         prince_inst_sbox_inst12_yxxx_inst_n48,
         prince_inst_sbox_inst12_yxxx_inst_n47,
         prince_inst_sbox_inst12_yxxx_inst_n46,
         prince_inst_sbox_inst12_yxxx_inst_n45,
         prince_inst_sbox_inst12_yxyy_inst_n68,
         prince_inst_sbox_inst12_yxyy_inst_n67,
         prince_inst_sbox_inst12_yxyy_inst_n66,
         prince_inst_sbox_inst12_yxyy_inst_n65,
         prince_inst_sbox_inst12_yxyy_inst_n64,
         prince_inst_sbox_inst12_yxyy_inst_n63,
         prince_inst_sbox_inst12_yxyy_inst_n62,
         prince_inst_sbox_inst12_yxyy_inst_n61,
         prince_inst_sbox_inst12_yxyy_inst_n60,
         prince_inst_sbox_inst12_yxyy_inst_n59,
         prince_inst_sbox_inst12_yxyy_inst_n58,
         prince_inst_sbox_inst12_yxyy_inst_n57,
         prince_inst_sbox_inst12_yxyy_inst_n56,
         prince_inst_sbox_inst12_yxyy_inst_n55,
         prince_inst_sbox_inst12_yxyy_inst_n54,
         prince_inst_sbox_inst12_yxyy_inst_n53,
         prince_inst_sbox_inst12_yxyy_inst_n52,
         prince_inst_sbox_inst12_yxyy_inst_n51,
         prince_inst_sbox_inst12_yxyy_inst_n50,
         prince_inst_sbox_inst12_yxyy_inst_n49,
         prince_inst_sbox_inst12_yyxy_inst_n75,
         prince_inst_sbox_inst12_yyxy_inst_n74,
         prince_inst_sbox_inst12_yyxy_inst_n73,
         prince_inst_sbox_inst12_yyxy_inst_n72,
         prince_inst_sbox_inst12_yyxy_inst_n71,
         prince_inst_sbox_inst12_yyxy_inst_n70,
         prince_inst_sbox_inst12_yyxy_inst_n69,
         prince_inst_sbox_inst12_yyxy_inst_n68,
         prince_inst_sbox_inst12_yyxy_inst_n67,
         prince_inst_sbox_inst12_yyxy_inst_n66,
         prince_inst_sbox_inst12_yyxy_inst_n65,
         prince_inst_sbox_inst12_yyxy_inst_n64,
         prince_inst_sbox_inst12_yyxy_inst_n63,
         prince_inst_sbox_inst12_yyxy_inst_n62,
         prince_inst_sbox_inst12_yyxy_inst_n61,
         prince_inst_sbox_inst12_yyxy_inst_n60,
         prince_inst_sbox_inst12_yyxy_inst_n59,
         prince_inst_sbox_inst12_yyxy_inst_n58,
         prince_inst_sbox_inst12_yyxy_inst_n57,
         prince_inst_sbox_inst12_yyxy_inst_n56,
         prince_inst_sbox_inst12_yyxy_inst_n55,
         prince_inst_sbox_inst12_yyxy_inst_n54,
         prince_inst_sbox_inst12_yyxy_inst_n53,
         prince_inst_sbox_inst12_yyyx_inst_n58,
         prince_inst_sbox_inst12_yyyx_inst_n57,
         prince_inst_sbox_inst12_yyyx_inst_n56,
         prince_inst_sbox_inst12_yyyx_inst_n55,
         prince_inst_sbox_inst12_yyyx_inst_n54,
         prince_inst_sbox_inst12_yyyx_inst_n53,
         prince_inst_sbox_inst12_yyyx_inst_n52,
         prince_inst_sbox_inst12_yyyx_inst_n51,
         prince_inst_sbox_inst12_yyyx_inst_n50,
         prince_inst_sbox_inst12_yyyx_inst_n49,
         prince_inst_sbox_inst12_yyyx_inst_n48,
         prince_inst_sbox_inst12_yyyx_inst_n47,
         prince_inst_sbox_inst12_yyyx_inst_n46,
         prince_inst_sbox_inst12_yyyx_inst_n45,
         prince_inst_sbox_inst12_yyyx_inst_n44,
         prince_inst_sbox_inst12_yyyx_inst_n43,
         prince_inst_sbox_inst12_yyyx_inst_n42,
         prince_inst_sbox_inst12_c_inst0_msk0_xr,
         prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_msk1_xr,
         prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_msk2_xr,
         prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_msk3_xr,
         prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_msk4_xr,
         prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_msk5_xr,
         prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_msk6_xr,
         prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_msk7_xr,
         prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst0_ax_n6,
         prince_inst_sbox_inst12_c_inst0_ax_n5,
         prince_inst_sbox_inst12_c_inst0_ay_n6,
         prince_inst_sbox_inst12_c_inst0_ay_n5,
         prince_inst_sbox_inst12_c_inst1_msk0_xr,
         prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_msk1_xr,
         prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_msk2_xr,
         prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_msk3_xr,
         prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_msk4_xr,
         prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_msk5_xr,
         prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_msk6_xr,
         prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_msk7_xr,
         prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst1_ax_n6,
         prince_inst_sbox_inst12_c_inst1_ax_n5,
         prince_inst_sbox_inst12_c_inst1_ay_n6,
         prince_inst_sbox_inst12_c_inst1_ay_n5,
         prince_inst_sbox_inst12_c_inst2_msk0_xr,
         prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_msk1_xr,
         prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_msk2_xr,
         prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_msk3_xr,
         prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_msk4_xr,
         prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_msk5_xr,
         prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_msk6_xr,
         prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_msk7_xr,
         prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst2_ax_n6,
         prince_inst_sbox_inst12_c_inst2_ax_n5,
         prince_inst_sbox_inst12_c_inst2_ay_n6,
         prince_inst_sbox_inst12_c_inst2_ay_n5,
         prince_inst_sbox_inst12_c_inst3_msk0_xr,
         prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_msk1_xr,
         prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_msk2_xr,
         prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_msk3_xr,
         prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_msk4_xr,
         prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_msk5_xr,
         prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_msk6_xr,
         prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_msk7_xr,
         prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst12_c_inst3_ax_n6,
         prince_inst_sbox_inst12_c_inst3_ax_n5,
         prince_inst_sbox_inst12_c_inst3_ay_n6,
         prince_inst_sbox_inst12_c_inst3_ay_n5, prince_inst_sbox_inst13_n13,
         prince_inst_sbox_inst13_n12, prince_inst_sbox_inst13_n11,
         prince_inst_sbox_inst13_n10, prince_inst_sbox_inst13_n9,
         prince_inst_sbox_inst13_n8, prince_inst_sbox_inst13_n7,
         prince_inst_sbox_inst13_xxxy_inst_n69,
         prince_inst_sbox_inst13_xxxy_inst_n68,
         prince_inst_sbox_inst13_xxxy_inst_n67,
         prince_inst_sbox_inst13_xxxy_inst_n66,
         prince_inst_sbox_inst13_xxxy_inst_n65,
         prince_inst_sbox_inst13_xxxy_inst_n64,
         prince_inst_sbox_inst13_xxxy_inst_n63,
         prince_inst_sbox_inst13_xxxy_inst_n62,
         prince_inst_sbox_inst13_xxxy_inst_n61,
         prince_inst_sbox_inst13_xxxy_inst_n60,
         prince_inst_sbox_inst13_xxxy_inst_n59,
         prince_inst_sbox_inst13_xxxy_inst_n58,
         prince_inst_sbox_inst13_xxxy_inst_n57,
         prince_inst_sbox_inst13_xxxy_inst_n56,
         prince_inst_sbox_inst13_xxxy_inst_n55,
         prince_inst_sbox_inst13_xxxy_inst_n54,
         prince_inst_sbox_inst13_xxxy_inst_n53,
         prince_inst_sbox_inst13_xxxy_inst_n52,
         prince_inst_sbox_inst13_xxxy_inst_n51,
         prince_inst_sbox_inst13_xxyx_inst_n55,
         prince_inst_sbox_inst13_xxyx_inst_n54,
         prince_inst_sbox_inst13_xxyx_inst_n53,
         prince_inst_sbox_inst13_xxyx_inst_n52,
         prince_inst_sbox_inst13_xxyx_inst_n51,
         prince_inst_sbox_inst13_xxyx_inst_n50,
         prince_inst_sbox_inst13_xxyx_inst_n49,
         prince_inst_sbox_inst13_xxyx_inst_n48,
         prince_inst_sbox_inst13_xxyx_inst_n47,
         prince_inst_sbox_inst13_xxyx_inst_n46,
         prince_inst_sbox_inst13_xxyx_inst_n45,
         prince_inst_sbox_inst13_xxyx_inst_n44,
         prince_inst_sbox_inst13_xxyx_inst_n43,
         prince_inst_sbox_inst13_xxyx_inst_n42,
         prince_inst_sbox_inst13_xxyx_inst_n41,
         prince_inst_sbox_inst13_xxyx_inst_n40,
         prince_inst_sbox_inst13_xxyx_inst_n39,
         prince_inst_sbox_inst13_xxyx_inst_n38,
         prince_inst_sbox_inst13_xyxx_inst_n74,
         prince_inst_sbox_inst13_xyxx_inst_n73,
         prince_inst_sbox_inst13_xyxx_inst_n72,
         prince_inst_sbox_inst13_xyxx_inst_n71,
         prince_inst_sbox_inst13_xyxx_inst_n70,
         prince_inst_sbox_inst13_xyxx_inst_n69,
         prince_inst_sbox_inst13_xyxx_inst_n68,
         prince_inst_sbox_inst13_xyxx_inst_n67,
         prince_inst_sbox_inst13_xyxx_inst_n66,
         prince_inst_sbox_inst13_xyxx_inst_n65,
         prince_inst_sbox_inst13_xyxx_inst_n64,
         prince_inst_sbox_inst13_xyxx_inst_n63,
         prince_inst_sbox_inst13_xyxx_inst_n62,
         prince_inst_sbox_inst13_xyxx_inst_n61,
         prince_inst_sbox_inst13_xyxx_inst_n60,
         prince_inst_sbox_inst13_xyxx_inst_n59,
         prince_inst_sbox_inst13_xyxx_inst_n58,
         prince_inst_sbox_inst13_xyxx_inst_n57,
         prince_inst_sbox_inst13_xyxx_inst_n56,
         prince_inst_sbox_inst13_xyxx_inst_n55,
         prince_inst_sbox_inst13_xyxx_inst_n54,
         prince_inst_sbox_inst13_xyxx_inst_n53,
         prince_inst_sbox_inst13_xyyy_inst_n61,
         prince_inst_sbox_inst13_xyyy_inst_n60,
         prince_inst_sbox_inst13_xyyy_inst_n59,
         prince_inst_sbox_inst13_xyyy_inst_n58,
         prince_inst_sbox_inst13_xyyy_inst_n57,
         prince_inst_sbox_inst13_xyyy_inst_n56,
         prince_inst_sbox_inst13_xyyy_inst_n55,
         prince_inst_sbox_inst13_xyyy_inst_n54,
         prince_inst_sbox_inst13_xyyy_inst_n53,
         prince_inst_sbox_inst13_xyyy_inst_n52,
         prince_inst_sbox_inst13_xyyy_inst_n51,
         prince_inst_sbox_inst13_xyyy_inst_n50,
         prince_inst_sbox_inst13_xyyy_inst_n49,
         prince_inst_sbox_inst13_xyyy_inst_n48,
         prince_inst_sbox_inst13_xyyy_inst_n47,
         prince_inst_sbox_inst13_xyyy_inst_n46,
         prince_inst_sbox_inst13_xyyy_inst_n45,
         prince_inst_sbox_inst13_xyyy_inst_n44,
         prince_inst_sbox_inst13_xyyy_inst_n43,
         prince_inst_sbox_inst13_xyyy_inst_n42,
         prince_inst_sbox_inst13_yxxx_inst_n64,
         prince_inst_sbox_inst13_yxxx_inst_n63,
         prince_inst_sbox_inst13_yxxx_inst_n62,
         prince_inst_sbox_inst13_yxxx_inst_n61,
         prince_inst_sbox_inst13_yxxx_inst_n60,
         prince_inst_sbox_inst13_yxxx_inst_n59,
         prince_inst_sbox_inst13_yxxx_inst_n58,
         prince_inst_sbox_inst13_yxxx_inst_n57,
         prince_inst_sbox_inst13_yxxx_inst_n56,
         prince_inst_sbox_inst13_yxxx_inst_n55,
         prince_inst_sbox_inst13_yxxx_inst_n54,
         prince_inst_sbox_inst13_yxxx_inst_n53,
         prince_inst_sbox_inst13_yxxx_inst_n52,
         prince_inst_sbox_inst13_yxxx_inst_n51,
         prince_inst_sbox_inst13_yxxx_inst_n50,
         prince_inst_sbox_inst13_yxxx_inst_n49,
         prince_inst_sbox_inst13_yxxx_inst_n48,
         prince_inst_sbox_inst13_yxxx_inst_n47,
         prince_inst_sbox_inst13_yxxx_inst_n46,
         prince_inst_sbox_inst13_yxxx_inst_n45,
         prince_inst_sbox_inst13_yxyy_inst_n68,
         prince_inst_sbox_inst13_yxyy_inst_n67,
         prince_inst_sbox_inst13_yxyy_inst_n66,
         prince_inst_sbox_inst13_yxyy_inst_n65,
         prince_inst_sbox_inst13_yxyy_inst_n64,
         prince_inst_sbox_inst13_yxyy_inst_n63,
         prince_inst_sbox_inst13_yxyy_inst_n62,
         prince_inst_sbox_inst13_yxyy_inst_n61,
         prince_inst_sbox_inst13_yxyy_inst_n60,
         prince_inst_sbox_inst13_yxyy_inst_n59,
         prince_inst_sbox_inst13_yxyy_inst_n58,
         prince_inst_sbox_inst13_yxyy_inst_n57,
         prince_inst_sbox_inst13_yxyy_inst_n56,
         prince_inst_sbox_inst13_yxyy_inst_n55,
         prince_inst_sbox_inst13_yxyy_inst_n54,
         prince_inst_sbox_inst13_yxyy_inst_n53,
         prince_inst_sbox_inst13_yxyy_inst_n52,
         prince_inst_sbox_inst13_yxyy_inst_n51,
         prince_inst_sbox_inst13_yxyy_inst_n50,
         prince_inst_sbox_inst13_yxyy_inst_n49,
         prince_inst_sbox_inst13_yyxy_inst_n75,
         prince_inst_sbox_inst13_yyxy_inst_n74,
         prince_inst_sbox_inst13_yyxy_inst_n73,
         prince_inst_sbox_inst13_yyxy_inst_n72,
         prince_inst_sbox_inst13_yyxy_inst_n71,
         prince_inst_sbox_inst13_yyxy_inst_n70,
         prince_inst_sbox_inst13_yyxy_inst_n69,
         prince_inst_sbox_inst13_yyxy_inst_n68,
         prince_inst_sbox_inst13_yyxy_inst_n67,
         prince_inst_sbox_inst13_yyxy_inst_n66,
         prince_inst_sbox_inst13_yyxy_inst_n65,
         prince_inst_sbox_inst13_yyxy_inst_n64,
         prince_inst_sbox_inst13_yyxy_inst_n63,
         prince_inst_sbox_inst13_yyxy_inst_n62,
         prince_inst_sbox_inst13_yyxy_inst_n61,
         prince_inst_sbox_inst13_yyxy_inst_n60,
         prince_inst_sbox_inst13_yyxy_inst_n59,
         prince_inst_sbox_inst13_yyxy_inst_n58,
         prince_inst_sbox_inst13_yyxy_inst_n57,
         prince_inst_sbox_inst13_yyxy_inst_n56,
         prince_inst_sbox_inst13_yyxy_inst_n55,
         prince_inst_sbox_inst13_yyxy_inst_n54,
         prince_inst_sbox_inst13_yyxy_inst_n53,
         prince_inst_sbox_inst13_yyyx_inst_n58,
         prince_inst_sbox_inst13_yyyx_inst_n57,
         prince_inst_sbox_inst13_yyyx_inst_n56,
         prince_inst_sbox_inst13_yyyx_inst_n55,
         prince_inst_sbox_inst13_yyyx_inst_n54,
         prince_inst_sbox_inst13_yyyx_inst_n53,
         prince_inst_sbox_inst13_yyyx_inst_n52,
         prince_inst_sbox_inst13_yyyx_inst_n51,
         prince_inst_sbox_inst13_yyyx_inst_n50,
         prince_inst_sbox_inst13_yyyx_inst_n49,
         prince_inst_sbox_inst13_yyyx_inst_n48,
         prince_inst_sbox_inst13_yyyx_inst_n47,
         prince_inst_sbox_inst13_yyyx_inst_n46,
         prince_inst_sbox_inst13_yyyx_inst_n45,
         prince_inst_sbox_inst13_yyyx_inst_n44,
         prince_inst_sbox_inst13_yyyx_inst_n43,
         prince_inst_sbox_inst13_yyyx_inst_n42,
         prince_inst_sbox_inst13_c_inst0_msk0_xr,
         prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_msk1_xr,
         prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_msk2_xr,
         prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_msk3_xr,
         prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_msk4_xr,
         prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_msk5_xr,
         prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_msk6_xr,
         prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_msk7_xr,
         prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst0_ax_n6,
         prince_inst_sbox_inst13_c_inst0_ax_n5,
         prince_inst_sbox_inst13_c_inst0_ay_n6,
         prince_inst_sbox_inst13_c_inst0_ay_n5,
         prince_inst_sbox_inst13_c_inst1_msk0_xr,
         prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_msk1_xr,
         prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_msk2_xr,
         prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_msk3_xr,
         prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_msk4_xr,
         prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_msk5_xr,
         prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_msk6_xr,
         prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_msk7_xr,
         prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst1_ax_n6,
         prince_inst_sbox_inst13_c_inst1_ax_n5,
         prince_inst_sbox_inst13_c_inst1_ay_n6,
         prince_inst_sbox_inst13_c_inst1_ay_n5,
         prince_inst_sbox_inst13_c_inst2_msk0_xr,
         prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_msk1_xr,
         prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_msk2_xr,
         prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_msk3_xr,
         prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_msk4_xr,
         prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_msk5_xr,
         prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_msk6_xr,
         prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_msk7_xr,
         prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst2_ax_n6,
         prince_inst_sbox_inst13_c_inst2_ax_n5,
         prince_inst_sbox_inst13_c_inst2_ay_n6,
         prince_inst_sbox_inst13_c_inst2_ay_n5,
         prince_inst_sbox_inst13_c_inst3_msk0_xr,
         prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_msk1_xr,
         prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_msk2_xr,
         prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_msk3_xr,
         prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_msk4_xr,
         prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_msk5_xr,
         prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_msk6_xr,
         prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_msk7_xr,
         prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst13_c_inst3_ax_n6,
         prince_inst_sbox_inst13_c_inst3_ax_n5,
         prince_inst_sbox_inst13_c_inst3_ay_n6,
         prince_inst_sbox_inst13_c_inst3_ay_n5, prince_inst_sbox_inst14_n13,
         prince_inst_sbox_inst14_n12, prince_inst_sbox_inst14_n11,
         prince_inst_sbox_inst14_n10, prince_inst_sbox_inst14_n9,
         prince_inst_sbox_inst14_n8, prince_inst_sbox_inst14_n7,
         prince_inst_sbox_inst14_xxxy_inst_n69,
         prince_inst_sbox_inst14_xxxy_inst_n68,
         prince_inst_sbox_inst14_xxxy_inst_n67,
         prince_inst_sbox_inst14_xxxy_inst_n66,
         prince_inst_sbox_inst14_xxxy_inst_n65,
         prince_inst_sbox_inst14_xxxy_inst_n64,
         prince_inst_sbox_inst14_xxxy_inst_n63,
         prince_inst_sbox_inst14_xxxy_inst_n62,
         prince_inst_sbox_inst14_xxxy_inst_n61,
         prince_inst_sbox_inst14_xxxy_inst_n60,
         prince_inst_sbox_inst14_xxxy_inst_n59,
         prince_inst_sbox_inst14_xxxy_inst_n58,
         prince_inst_sbox_inst14_xxxy_inst_n57,
         prince_inst_sbox_inst14_xxxy_inst_n56,
         prince_inst_sbox_inst14_xxxy_inst_n55,
         prince_inst_sbox_inst14_xxxy_inst_n54,
         prince_inst_sbox_inst14_xxxy_inst_n53,
         prince_inst_sbox_inst14_xxxy_inst_n52,
         prince_inst_sbox_inst14_xxxy_inst_n51,
         prince_inst_sbox_inst14_xxyx_inst_n55,
         prince_inst_sbox_inst14_xxyx_inst_n54,
         prince_inst_sbox_inst14_xxyx_inst_n53,
         prince_inst_sbox_inst14_xxyx_inst_n52,
         prince_inst_sbox_inst14_xxyx_inst_n51,
         prince_inst_sbox_inst14_xxyx_inst_n50,
         prince_inst_sbox_inst14_xxyx_inst_n49,
         prince_inst_sbox_inst14_xxyx_inst_n48,
         prince_inst_sbox_inst14_xxyx_inst_n47,
         prince_inst_sbox_inst14_xxyx_inst_n46,
         prince_inst_sbox_inst14_xxyx_inst_n45,
         prince_inst_sbox_inst14_xxyx_inst_n44,
         prince_inst_sbox_inst14_xxyx_inst_n43,
         prince_inst_sbox_inst14_xxyx_inst_n42,
         prince_inst_sbox_inst14_xxyx_inst_n41,
         prince_inst_sbox_inst14_xxyx_inst_n40,
         prince_inst_sbox_inst14_xxyx_inst_n39,
         prince_inst_sbox_inst14_xxyx_inst_n38,
         prince_inst_sbox_inst14_xyxx_inst_n74,
         prince_inst_sbox_inst14_xyxx_inst_n73,
         prince_inst_sbox_inst14_xyxx_inst_n72,
         prince_inst_sbox_inst14_xyxx_inst_n71,
         prince_inst_sbox_inst14_xyxx_inst_n70,
         prince_inst_sbox_inst14_xyxx_inst_n69,
         prince_inst_sbox_inst14_xyxx_inst_n68,
         prince_inst_sbox_inst14_xyxx_inst_n67,
         prince_inst_sbox_inst14_xyxx_inst_n66,
         prince_inst_sbox_inst14_xyxx_inst_n65,
         prince_inst_sbox_inst14_xyxx_inst_n64,
         prince_inst_sbox_inst14_xyxx_inst_n63,
         prince_inst_sbox_inst14_xyxx_inst_n62,
         prince_inst_sbox_inst14_xyxx_inst_n61,
         prince_inst_sbox_inst14_xyxx_inst_n60,
         prince_inst_sbox_inst14_xyxx_inst_n59,
         prince_inst_sbox_inst14_xyxx_inst_n58,
         prince_inst_sbox_inst14_xyxx_inst_n57,
         prince_inst_sbox_inst14_xyxx_inst_n56,
         prince_inst_sbox_inst14_xyxx_inst_n55,
         prince_inst_sbox_inst14_xyxx_inst_n54,
         prince_inst_sbox_inst14_xyxx_inst_n53,
         prince_inst_sbox_inst14_xyyy_inst_n61,
         prince_inst_sbox_inst14_xyyy_inst_n60,
         prince_inst_sbox_inst14_xyyy_inst_n59,
         prince_inst_sbox_inst14_xyyy_inst_n58,
         prince_inst_sbox_inst14_xyyy_inst_n57,
         prince_inst_sbox_inst14_xyyy_inst_n56,
         prince_inst_sbox_inst14_xyyy_inst_n55,
         prince_inst_sbox_inst14_xyyy_inst_n54,
         prince_inst_sbox_inst14_xyyy_inst_n53,
         prince_inst_sbox_inst14_xyyy_inst_n52,
         prince_inst_sbox_inst14_xyyy_inst_n51,
         prince_inst_sbox_inst14_xyyy_inst_n50,
         prince_inst_sbox_inst14_xyyy_inst_n49,
         prince_inst_sbox_inst14_xyyy_inst_n48,
         prince_inst_sbox_inst14_xyyy_inst_n47,
         prince_inst_sbox_inst14_xyyy_inst_n46,
         prince_inst_sbox_inst14_xyyy_inst_n45,
         prince_inst_sbox_inst14_xyyy_inst_n44,
         prince_inst_sbox_inst14_xyyy_inst_n43,
         prince_inst_sbox_inst14_xyyy_inst_n42,
         prince_inst_sbox_inst14_yxxx_inst_n64,
         prince_inst_sbox_inst14_yxxx_inst_n63,
         prince_inst_sbox_inst14_yxxx_inst_n62,
         prince_inst_sbox_inst14_yxxx_inst_n61,
         prince_inst_sbox_inst14_yxxx_inst_n60,
         prince_inst_sbox_inst14_yxxx_inst_n59,
         prince_inst_sbox_inst14_yxxx_inst_n58,
         prince_inst_sbox_inst14_yxxx_inst_n57,
         prince_inst_sbox_inst14_yxxx_inst_n56,
         prince_inst_sbox_inst14_yxxx_inst_n55,
         prince_inst_sbox_inst14_yxxx_inst_n54,
         prince_inst_sbox_inst14_yxxx_inst_n53,
         prince_inst_sbox_inst14_yxxx_inst_n52,
         prince_inst_sbox_inst14_yxxx_inst_n51,
         prince_inst_sbox_inst14_yxxx_inst_n50,
         prince_inst_sbox_inst14_yxxx_inst_n49,
         prince_inst_sbox_inst14_yxxx_inst_n48,
         prince_inst_sbox_inst14_yxxx_inst_n47,
         prince_inst_sbox_inst14_yxxx_inst_n46,
         prince_inst_sbox_inst14_yxxx_inst_n45,
         prince_inst_sbox_inst14_yxyy_inst_n68,
         prince_inst_sbox_inst14_yxyy_inst_n67,
         prince_inst_sbox_inst14_yxyy_inst_n66,
         prince_inst_sbox_inst14_yxyy_inst_n65,
         prince_inst_sbox_inst14_yxyy_inst_n64,
         prince_inst_sbox_inst14_yxyy_inst_n63,
         prince_inst_sbox_inst14_yxyy_inst_n62,
         prince_inst_sbox_inst14_yxyy_inst_n61,
         prince_inst_sbox_inst14_yxyy_inst_n60,
         prince_inst_sbox_inst14_yxyy_inst_n59,
         prince_inst_sbox_inst14_yxyy_inst_n58,
         prince_inst_sbox_inst14_yxyy_inst_n57,
         prince_inst_sbox_inst14_yxyy_inst_n56,
         prince_inst_sbox_inst14_yxyy_inst_n55,
         prince_inst_sbox_inst14_yxyy_inst_n54,
         prince_inst_sbox_inst14_yxyy_inst_n53,
         prince_inst_sbox_inst14_yxyy_inst_n52,
         prince_inst_sbox_inst14_yxyy_inst_n51,
         prince_inst_sbox_inst14_yxyy_inst_n50,
         prince_inst_sbox_inst14_yxyy_inst_n49,
         prince_inst_sbox_inst14_yyxy_inst_n75,
         prince_inst_sbox_inst14_yyxy_inst_n74,
         prince_inst_sbox_inst14_yyxy_inst_n73,
         prince_inst_sbox_inst14_yyxy_inst_n72,
         prince_inst_sbox_inst14_yyxy_inst_n71,
         prince_inst_sbox_inst14_yyxy_inst_n70,
         prince_inst_sbox_inst14_yyxy_inst_n69,
         prince_inst_sbox_inst14_yyxy_inst_n68,
         prince_inst_sbox_inst14_yyxy_inst_n67,
         prince_inst_sbox_inst14_yyxy_inst_n66,
         prince_inst_sbox_inst14_yyxy_inst_n65,
         prince_inst_sbox_inst14_yyxy_inst_n64,
         prince_inst_sbox_inst14_yyxy_inst_n63,
         prince_inst_sbox_inst14_yyxy_inst_n62,
         prince_inst_sbox_inst14_yyxy_inst_n61,
         prince_inst_sbox_inst14_yyxy_inst_n60,
         prince_inst_sbox_inst14_yyxy_inst_n59,
         prince_inst_sbox_inst14_yyxy_inst_n58,
         prince_inst_sbox_inst14_yyxy_inst_n57,
         prince_inst_sbox_inst14_yyxy_inst_n56,
         prince_inst_sbox_inst14_yyxy_inst_n55,
         prince_inst_sbox_inst14_yyxy_inst_n54,
         prince_inst_sbox_inst14_yyxy_inst_n53,
         prince_inst_sbox_inst14_yyyx_inst_n58,
         prince_inst_sbox_inst14_yyyx_inst_n57,
         prince_inst_sbox_inst14_yyyx_inst_n56,
         prince_inst_sbox_inst14_yyyx_inst_n55,
         prince_inst_sbox_inst14_yyyx_inst_n54,
         prince_inst_sbox_inst14_yyyx_inst_n53,
         prince_inst_sbox_inst14_yyyx_inst_n52,
         prince_inst_sbox_inst14_yyyx_inst_n51,
         prince_inst_sbox_inst14_yyyx_inst_n50,
         prince_inst_sbox_inst14_yyyx_inst_n49,
         prince_inst_sbox_inst14_yyyx_inst_n48,
         prince_inst_sbox_inst14_yyyx_inst_n47,
         prince_inst_sbox_inst14_yyyx_inst_n46,
         prince_inst_sbox_inst14_yyyx_inst_n45,
         prince_inst_sbox_inst14_yyyx_inst_n44,
         prince_inst_sbox_inst14_yyyx_inst_n43,
         prince_inst_sbox_inst14_yyyx_inst_n42,
         prince_inst_sbox_inst14_c_inst0_msk0_xr,
         prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_msk1_xr,
         prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_msk2_xr,
         prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_msk3_xr,
         prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_msk4_xr,
         prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_msk5_xr,
         prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_msk6_xr,
         prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_msk7_xr,
         prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst0_ax_n6,
         prince_inst_sbox_inst14_c_inst0_ax_n5,
         prince_inst_sbox_inst14_c_inst0_ay_n6,
         prince_inst_sbox_inst14_c_inst0_ay_n5,
         prince_inst_sbox_inst14_c_inst1_msk0_xr,
         prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_msk1_xr,
         prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_msk2_xr,
         prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_msk3_xr,
         prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_msk4_xr,
         prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_msk5_xr,
         prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_msk6_xr,
         prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_msk7_xr,
         prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst1_ax_n6,
         prince_inst_sbox_inst14_c_inst1_ax_n5,
         prince_inst_sbox_inst14_c_inst1_ay_n6,
         prince_inst_sbox_inst14_c_inst1_ay_n5,
         prince_inst_sbox_inst14_c_inst2_msk0_xr,
         prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_msk1_xr,
         prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_msk2_xr,
         prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_msk3_xr,
         prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_msk4_xr,
         prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_msk5_xr,
         prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_msk6_xr,
         prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_msk7_xr,
         prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst2_ax_n6,
         prince_inst_sbox_inst14_c_inst2_ax_n5,
         prince_inst_sbox_inst14_c_inst2_ay_n6,
         prince_inst_sbox_inst14_c_inst2_ay_n5,
         prince_inst_sbox_inst14_c_inst3_msk0_xr,
         prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_msk1_xr,
         prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_msk2_xr,
         prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_msk3_xr,
         prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_msk4_xr,
         prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_msk5_xr,
         prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_msk6_xr,
         prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_msk7_xr,
         prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst14_c_inst3_ax_n6,
         prince_inst_sbox_inst14_c_inst3_ax_n5,
         prince_inst_sbox_inst14_c_inst3_ay_n6,
         prince_inst_sbox_inst14_c_inst3_ay_n5, prince_inst_sbox_inst15_n10,
         prince_inst_sbox_inst15_n9, prince_inst_sbox_inst15_n8,
         prince_inst_sbox_inst15_n7, prince_inst_sbox_inst15_n6,
         prince_inst_sbox_inst15_xxxy_inst_n69,
         prince_inst_sbox_inst15_xxxy_inst_n68,
         prince_inst_sbox_inst15_xxxy_inst_n67,
         prince_inst_sbox_inst15_xxxy_inst_n66,
         prince_inst_sbox_inst15_xxxy_inst_n65,
         prince_inst_sbox_inst15_xxxy_inst_n64,
         prince_inst_sbox_inst15_xxxy_inst_n63,
         prince_inst_sbox_inst15_xxxy_inst_n62,
         prince_inst_sbox_inst15_xxxy_inst_n61,
         prince_inst_sbox_inst15_xxxy_inst_n60,
         prince_inst_sbox_inst15_xxxy_inst_n59,
         prince_inst_sbox_inst15_xxxy_inst_n58,
         prince_inst_sbox_inst15_xxxy_inst_n57,
         prince_inst_sbox_inst15_xxxy_inst_n56,
         prince_inst_sbox_inst15_xxxy_inst_n55,
         prince_inst_sbox_inst15_xxxy_inst_n54,
         prince_inst_sbox_inst15_xxxy_inst_n53,
         prince_inst_sbox_inst15_xxxy_inst_n52,
         prince_inst_sbox_inst15_xxxy_inst_n51,
         prince_inst_sbox_inst15_xxyx_inst_n55,
         prince_inst_sbox_inst15_xxyx_inst_n54,
         prince_inst_sbox_inst15_xxyx_inst_n53,
         prince_inst_sbox_inst15_xxyx_inst_n52,
         prince_inst_sbox_inst15_xxyx_inst_n51,
         prince_inst_sbox_inst15_xxyx_inst_n50,
         prince_inst_sbox_inst15_xxyx_inst_n49,
         prince_inst_sbox_inst15_xxyx_inst_n48,
         prince_inst_sbox_inst15_xxyx_inst_n47,
         prince_inst_sbox_inst15_xxyx_inst_n46,
         prince_inst_sbox_inst15_xxyx_inst_n45,
         prince_inst_sbox_inst15_xxyx_inst_n44,
         prince_inst_sbox_inst15_xxyx_inst_n43,
         prince_inst_sbox_inst15_xxyx_inst_n42,
         prince_inst_sbox_inst15_xxyx_inst_n41,
         prince_inst_sbox_inst15_xxyx_inst_n40,
         prince_inst_sbox_inst15_xxyx_inst_n39,
         prince_inst_sbox_inst15_xxyx_inst_n38,
         prince_inst_sbox_inst15_xyxx_inst_n74,
         prince_inst_sbox_inst15_xyxx_inst_n73,
         prince_inst_sbox_inst15_xyxx_inst_n72,
         prince_inst_sbox_inst15_xyxx_inst_n71,
         prince_inst_sbox_inst15_xyxx_inst_n70,
         prince_inst_sbox_inst15_xyxx_inst_n69,
         prince_inst_sbox_inst15_xyxx_inst_n68,
         prince_inst_sbox_inst15_xyxx_inst_n67,
         prince_inst_sbox_inst15_xyxx_inst_n66,
         prince_inst_sbox_inst15_xyxx_inst_n65,
         prince_inst_sbox_inst15_xyxx_inst_n64,
         prince_inst_sbox_inst15_xyxx_inst_n63,
         prince_inst_sbox_inst15_xyxx_inst_n62,
         prince_inst_sbox_inst15_xyxx_inst_n61,
         prince_inst_sbox_inst15_xyxx_inst_n60,
         prince_inst_sbox_inst15_xyxx_inst_n59,
         prince_inst_sbox_inst15_xyxx_inst_n58,
         prince_inst_sbox_inst15_xyxx_inst_n57,
         prince_inst_sbox_inst15_xyxx_inst_n56,
         prince_inst_sbox_inst15_xyxx_inst_n55,
         prince_inst_sbox_inst15_xyxx_inst_n54,
         prince_inst_sbox_inst15_xyxx_inst_n53,
         prince_inst_sbox_inst15_xyyy_inst_n61,
         prince_inst_sbox_inst15_xyyy_inst_n60,
         prince_inst_sbox_inst15_xyyy_inst_n59,
         prince_inst_sbox_inst15_xyyy_inst_n58,
         prince_inst_sbox_inst15_xyyy_inst_n57,
         prince_inst_sbox_inst15_xyyy_inst_n56,
         prince_inst_sbox_inst15_xyyy_inst_n55,
         prince_inst_sbox_inst15_xyyy_inst_n54,
         prince_inst_sbox_inst15_xyyy_inst_n53,
         prince_inst_sbox_inst15_xyyy_inst_n52,
         prince_inst_sbox_inst15_xyyy_inst_n51,
         prince_inst_sbox_inst15_xyyy_inst_n50,
         prince_inst_sbox_inst15_xyyy_inst_n49,
         prince_inst_sbox_inst15_xyyy_inst_n48,
         prince_inst_sbox_inst15_xyyy_inst_n47,
         prince_inst_sbox_inst15_xyyy_inst_n46,
         prince_inst_sbox_inst15_xyyy_inst_n45,
         prince_inst_sbox_inst15_xyyy_inst_n44,
         prince_inst_sbox_inst15_xyyy_inst_n43,
         prince_inst_sbox_inst15_xyyy_inst_n42,
         prince_inst_sbox_inst15_yxxx_inst_n64,
         prince_inst_sbox_inst15_yxxx_inst_n63,
         prince_inst_sbox_inst15_yxxx_inst_n62,
         prince_inst_sbox_inst15_yxxx_inst_n61,
         prince_inst_sbox_inst15_yxxx_inst_n60,
         prince_inst_sbox_inst15_yxxx_inst_n59,
         prince_inst_sbox_inst15_yxxx_inst_n58,
         prince_inst_sbox_inst15_yxxx_inst_n57,
         prince_inst_sbox_inst15_yxxx_inst_n56,
         prince_inst_sbox_inst15_yxxx_inst_n55,
         prince_inst_sbox_inst15_yxxx_inst_n54,
         prince_inst_sbox_inst15_yxxx_inst_n53,
         prince_inst_sbox_inst15_yxxx_inst_n52,
         prince_inst_sbox_inst15_yxxx_inst_n51,
         prince_inst_sbox_inst15_yxxx_inst_n50,
         prince_inst_sbox_inst15_yxxx_inst_n49,
         prince_inst_sbox_inst15_yxxx_inst_n48,
         prince_inst_sbox_inst15_yxxx_inst_n47,
         prince_inst_sbox_inst15_yxxx_inst_n46,
         prince_inst_sbox_inst15_yxxx_inst_n45,
         prince_inst_sbox_inst15_yxyy_inst_n68,
         prince_inst_sbox_inst15_yxyy_inst_n67,
         prince_inst_sbox_inst15_yxyy_inst_n66,
         prince_inst_sbox_inst15_yxyy_inst_n65,
         prince_inst_sbox_inst15_yxyy_inst_n64,
         prince_inst_sbox_inst15_yxyy_inst_n63,
         prince_inst_sbox_inst15_yxyy_inst_n62,
         prince_inst_sbox_inst15_yxyy_inst_n61,
         prince_inst_sbox_inst15_yxyy_inst_n60,
         prince_inst_sbox_inst15_yxyy_inst_n59,
         prince_inst_sbox_inst15_yxyy_inst_n58,
         prince_inst_sbox_inst15_yxyy_inst_n57,
         prince_inst_sbox_inst15_yxyy_inst_n56,
         prince_inst_sbox_inst15_yxyy_inst_n55,
         prince_inst_sbox_inst15_yxyy_inst_n54,
         prince_inst_sbox_inst15_yxyy_inst_n53,
         prince_inst_sbox_inst15_yxyy_inst_n52,
         prince_inst_sbox_inst15_yxyy_inst_n51,
         prince_inst_sbox_inst15_yxyy_inst_n50,
         prince_inst_sbox_inst15_yxyy_inst_n49,
         prince_inst_sbox_inst15_yyxy_inst_n75,
         prince_inst_sbox_inst15_yyxy_inst_n74,
         prince_inst_sbox_inst15_yyxy_inst_n73,
         prince_inst_sbox_inst15_yyxy_inst_n72,
         prince_inst_sbox_inst15_yyxy_inst_n71,
         prince_inst_sbox_inst15_yyxy_inst_n70,
         prince_inst_sbox_inst15_yyxy_inst_n69,
         prince_inst_sbox_inst15_yyxy_inst_n68,
         prince_inst_sbox_inst15_yyxy_inst_n67,
         prince_inst_sbox_inst15_yyxy_inst_n66,
         prince_inst_sbox_inst15_yyxy_inst_n65,
         prince_inst_sbox_inst15_yyxy_inst_n64,
         prince_inst_sbox_inst15_yyxy_inst_n63,
         prince_inst_sbox_inst15_yyxy_inst_n62,
         prince_inst_sbox_inst15_yyxy_inst_n61,
         prince_inst_sbox_inst15_yyxy_inst_n60,
         prince_inst_sbox_inst15_yyxy_inst_n59,
         prince_inst_sbox_inst15_yyxy_inst_n58,
         prince_inst_sbox_inst15_yyxy_inst_n57,
         prince_inst_sbox_inst15_yyxy_inst_n56,
         prince_inst_sbox_inst15_yyxy_inst_n55,
         prince_inst_sbox_inst15_yyxy_inst_n54,
         prince_inst_sbox_inst15_yyxy_inst_n53,
         prince_inst_sbox_inst15_yyyx_inst_n58,
         prince_inst_sbox_inst15_yyyx_inst_n57,
         prince_inst_sbox_inst15_yyyx_inst_n56,
         prince_inst_sbox_inst15_yyyx_inst_n55,
         prince_inst_sbox_inst15_yyyx_inst_n54,
         prince_inst_sbox_inst15_yyyx_inst_n53,
         prince_inst_sbox_inst15_yyyx_inst_n52,
         prince_inst_sbox_inst15_yyyx_inst_n51,
         prince_inst_sbox_inst15_yyyx_inst_n50,
         prince_inst_sbox_inst15_yyyx_inst_n49,
         prince_inst_sbox_inst15_yyyx_inst_n48,
         prince_inst_sbox_inst15_yyyx_inst_n47,
         prince_inst_sbox_inst15_yyyx_inst_n46,
         prince_inst_sbox_inst15_yyyx_inst_n45,
         prince_inst_sbox_inst15_yyyx_inst_n44,
         prince_inst_sbox_inst15_yyyx_inst_n43,
         prince_inst_sbox_inst15_yyyx_inst_n42,
         prince_inst_sbox_inst15_c_inst0_msk0_xr,
         prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_msk1_xr,
         prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_msk2_xr,
         prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_msk3_xr,
         prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_msk4_xr,
         prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_msk5_xr,
         prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_msk6_xr,
         prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_msk7_xr,
         prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst0_ax_n6,
         prince_inst_sbox_inst15_c_inst0_ax_n5,
         prince_inst_sbox_inst15_c_inst0_ay_n6,
         prince_inst_sbox_inst15_c_inst0_ay_n5,
         prince_inst_sbox_inst15_c_inst1_msk0_xr,
         prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_msk1_xr,
         prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_msk2_xr,
         prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_msk3_xr,
         prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_msk4_xr,
         prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_msk5_xr,
         prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_msk6_xr,
         prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_msk7_xr,
         prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst1_ax_n6,
         prince_inst_sbox_inst15_c_inst1_ax_n5,
         prince_inst_sbox_inst15_c_inst1_ay_n6,
         prince_inst_sbox_inst15_c_inst1_ay_n5,
         prince_inst_sbox_inst15_c_inst2_msk0_xr,
         prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_msk1_xr,
         prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_msk2_xr,
         prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_msk3_xr,
         prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_msk4_xr,
         prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_msk5_xr,
         prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_msk6_xr,
         prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_msk7_xr,
         prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst2_ax_n6,
         prince_inst_sbox_inst15_c_inst2_ax_n5,
         prince_inst_sbox_inst15_c_inst2_ay_n6,
         prince_inst_sbox_inst15_c_inst2_ay_n5,
         prince_inst_sbox_inst15_c_inst3_msk0_xr,
         prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_msk1_xr,
         prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_msk2_xr,
         prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_msk3_xr,
         prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_msk4_xr,
         prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_msk5_xr,
         prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_msk6_xr,
         prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_msk7_xr,
         prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n12,
         prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n11,
         prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n10,
         prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n6,
         prince_inst_sbox_inst15_c_inst3_ax_n6,
         prince_inst_sbox_inst15_c_inst3_ax_n5,
         prince_inst_sbox_inst15_c_inst3_ay_n6,
         prince_inst_sbox_inst15_c_inst3_ay_n5,
         prince_inst_mx_inst_m1_inst1_a0_n1,
         prince_inst_mx_inst_m1_inst1_a1_n3,
         prince_inst_mx_inst_m1_inst1_a2_n3,
         prince_inst_mx_inst_m1_inst1_a3_n3,
         prince_inst_mx_inst_m1_inst1_a4_n3,
         prince_inst_mx_inst_m1_inst1_a5_n3,
         prince_inst_mx_inst_m1_inst1_a6_n3,
         prince_inst_mx_inst_m1_inst1_a7_n3,
         prince_inst_mx_inst_m1_inst1_a8_n3,
         prince_inst_mx_inst_m1_inst1_a9_n3,
         prince_inst_mx_inst_m1_inst1_a10_n3,
         prince_inst_mx_inst_m1_inst1_a11_n3,
         prince_inst_mx_inst_m1_inst1_a12_n3,
         prince_inst_mx_inst_m1_inst1_a13_n3,
         prince_inst_mx_inst_m1_inst1_a14_n3,
         prince_inst_mx_inst_m1_inst1_a15_n3,
         prince_inst_mx_inst_m2_inst1_a0_n3,
         prince_inst_mx_inst_m2_inst1_a1_n3,
         prince_inst_mx_inst_m2_inst1_a2_n3,
         prince_inst_mx_inst_m2_inst1_a3_n3,
         prince_inst_mx_inst_m2_inst1_a4_n3,
         prince_inst_mx_inst_m2_inst1_a5_n3,
         prince_inst_mx_inst_m2_inst1_a6_n3,
         prince_inst_mx_inst_m2_inst1_a7_n3,
         prince_inst_mx_inst_m2_inst1_a8_n3,
         prince_inst_mx_inst_m2_inst1_a9_n3,
         prince_inst_mx_inst_m2_inst1_a10_n3,
         prince_inst_mx_inst_m2_inst1_a11_n3,
         prince_inst_mx_inst_m2_inst1_a12_n3,
         prince_inst_mx_inst_m2_inst1_a13_n3,
         prince_inst_mx_inst_m2_inst1_a14_n3,
         prince_inst_mx_inst_m2_inst1_a15_n3,
         prince_inst_mx_inst_m2_inst2_a0_n3,
         prince_inst_mx_inst_m2_inst2_a1_n3,
         prince_inst_mx_inst_m2_inst2_a2_n3,
         prince_inst_mx_inst_m2_inst2_a3_n3,
         prince_inst_mx_inst_m2_inst2_a4_n3,
         prince_inst_mx_inst_m2_inst2_a5_n3,
         prince_inst_mx_inst_m2_inst2_a6_n3,
         prince_inst_mx_inst_m2_inst2_a7_n3,
         prince_inst_mx_inst_m2_inst2_a8_n3,
         prince_inst_mx_inst_m2_inst2_a9_n3,
         prince_inst_mx_inst_m2_inst2_a10_n3,
         prince_inst_mx_inst_m2_inst2_a11_n3,
         prince_inst_mx_inst_m2_inst2_a12_n3,
         prince_inst_mx_inst_m2_inst2_a13_n3,
         prince_inst_mx_inst_m2_inst2_a14_n3,
         prince_inst_mx_inst_m2_inst2_a15_n3,
         prince_inst_mx_inst_m1_inst2_a0_n3,
         prince_inst_mx_inst_m1_inst2_a1_n3,
         prince_inst_mx_inst_m1_inst2_a2_n3,
         prince_inst_mx_inst_m1_inst2_a3_n3,
         prince_inst_mx_inst_m1_inst2_a4_n3,
         prince_inst_mx_inst_m1_inst2_a5_n3,
         prince_inst_mx_inst_m1_inst2_a6_n3,
         prince_inst_mx_inst_m1_inst2_a7_n3,
         prince_inst_mx_inst_m1_inst2_a8_n3,
         prince_inst_mx_inst_m1_inst2_a9_n3,
         prince_inst_mx_inst_m1_inst2_a10_n3,
         prince_inst_mx_inst_m1_inst2_a11_n3,
         prince_inst_mx_inst_m1_inst2_a12_n3,
         prince_inst_mx_inst_m1_inst2_a13_n3,
         prince_inst_mx_inst_m1_inst2_a14_n3,
         prince_inst_mx_inst_m1_inst2_a15_n3,
         prince_inst_my_inst_m1_inst1_a0_n3,
         prince_inst_my_inst_m1_inst1_a1_n3,
         prince_inst_my_inst_m1_inst1_a2_n3,
         prince_inst_my_inst_m1_inst1_a3_n3,
         prince_inst_my_inst_m1_inst1_a4_n3,
         prince_inst_my_inst_m1_inst1_a5_n3,
         prince_inst_my_inst_m1_inst1_a6_n3,
         prince_inst_my_inst_m1_inst1_a7_n3,
         prince_inst_my_inst_m1_inst1_a8_n3,
         prince_inst_my_inst_m1_inst1_a9_n3,
         prince_inst_my_inst_m1_inst1_a10_n3,
         prince_inst_my_inst_m1_inst1_a11_n3,
         prince_inst_my_inst_m1_inst1_a12_n3,
         prince_inst_my_inst_m1_inst1_a13_n3,
         prince_inst_my_inst_m1_inst1_a14_n3,
         prince_inst_my_inst_m1_inst1_a15_n3,
         prince_inst_my_inst_m2_inst1_a0_n3,
         prince_inst_my_inst_m2_inst1_a1_n3,
         prince_inst_my_inst_m2_inst1_a2_n3,
         prince_inst_my_inst_m2_inst1_a3_n3,
         prince_inst_my_inst_m2_inst1_a4_n3,
         prince_inst_my_inst_m2_inst1_a5_n3,
         prince_inst_my_inst_m2_inst1_a6_n3,
         prince_inst_my_inst_m2_inst1_a7_n3,
         prince_inst_my_inst_m2_inst1_a8_n3,
         prince_inst_my_inst_m2_inst1_a9_n3,
         prince_inst_my_inst_m2_inst1_a10_n3,
         prince_inst_my_inst_m2_inst1_a11_n3,
         prince_inst_my_inst_m2_inst1_a12_n3,
         prince_inst_my_inst_m2_inst1_a13_n3,
         prince_inst_my_inst_m2_inst1_a14_n3,
         prince_inst_my_inst_m2_inst1_a15_n3,
         prince_inst_my_inst_m2_inst2_a0_n3,
         prince_inst_my_inst_m2_inst2_a1_n3,
         prince_inst_my_inst_m2_inst2_a2_n3,
         prince_inst_my_inst_m2_inst2_a3_n3,
         prince_inst_my_inst_m2_inst2_a4_n3,
         prince_inst_my_inst_m2_inst2_a5_n3,
         prince_inst_my_inst_m2_inst2_a6_n3,
         prince_inst_my_inst_m2_inst2_a7_n3,
         prince_inst_my_inst_m2_inst2_a8_n3,
         prince_inst_my_inst_m2_inst2_a9_n3,
         prince_inst_my_inst_m2_inst2_a10_n3,
         prince_inst_my_inst_m2_inst2_a11_n3,
         prince_inst_my_inst_m2_inst2_a12_n3,
         prince_inst_my_inst_m2_inst2_a13_n3,
         prince_inst_my_inst_m2_inst2_a14_n3,
         prince_inst_my_inst_m2_inst2_a15_n3,
         prince_inst_my_inst_m1_inst2_a0_n3,
         prince_inst_my_inst_m1_inst2_a1_n3,
         prince_inst_my_inst_m1_inst2_a2_n3,
         prince_inst_my_inst_m1_inst2_a3_n3,
         prince_inst_my_inst_m1_inst2_a4_n3,
         prince_inst_my_inst_m1_inst2_a5_n3,
         prince_inst_my_inst_m1_inst2_a6_n3,
         prince_inst_my_inst_m1_inst2_a7_n3,
         prince_inst_my_inst_m1_inst2_a8_n3,
         prince_inst_my_inst_m1_inst2_a9_n3,
         prince_inst_my_inst_m1_inst2_a10_n3,
         prince_inst_my_inst_m1_inst2_a11_n3,
         prince_inst_my_inst_m1_inst2_a12_n3,
         prince_inst_my_inst_m1_inst2_a13_n3,
         prince_inst_my_inst_m1_inst2_a14_n3,
         prince_inst_my_inst_m1_inst2_a15_n3, mux_c0_n265, mux_c0_n264,
         mux_c0_n263, mux_c1_n264, mux_c1_n263, mux_c1_n262;
  wire   [191:1] kext;
  wire   [63:0] p0_reg;
  wire   [63:0] init_x;
  wire   [63:0] init_y;
  wire   [63:0] rout_x;
  wire   [63:0] rout_y;
  wire   [63:0] rc;
  wire   [63:0] final_x;
  wire   [63:0] final_y;
  wire   [63:0] final_x_k;
  wire   [63:0] prince_inst_min_y;
  wire   [63:0] prince_inst_min_x;
  wire   [63:0] prince_inst_sin_y;
  wire   [63:0] prince_inst_sin_x;
  wire   [63:0] prince_inst_sout_x;
  wire   [63:0] prince_inst_xout_x;
  wire   [63:0] prince_inst_srin_y;
  wire   [63:0] prince_inst_srin_x;
  wire   [63:0] prince_inst_rc2_inv;
  wire   [7:0] prince_inst_sbox_inst0_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst0_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst0_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst0_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst0_t3_sh;
  wire   [7:0] prince_inst_sbox_inst0_t2_sh;
  wire   [7:0] prince_inst_sbox_inst0_t1_sh;
  wire   [7:0] prince_inst_sbox_inst0_t0_sh;
  wire   [7:0] prince_inst_sbox_inst0_s3_sh;
  wire   [7:0] prince_inst_sbox_inst0_s2_sh;
  wire   [7:0] prince_inst_sbox_inst0_s1_sh;
  wire   [7:0] prince_inst_sbox_inst0_s0_sh;
  wire   [7:0] prince_inst_sbox_inst0_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst0_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst0_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst0_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst1_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst1_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst1_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst1_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst1_t3_sh;
  wire   [7:0] prince_inst_sbox_inst1_t2_sh;
  wire   [7:0] prince_inst_sbox_inst1_t1_sh;
  wire   [7:0] prince_inst_sbox_inst1_t0_sh;
  wire   [7:0] prince_inst_sbox_inst1_s3_sh;
  wire   [7:0] prince_inst_sbox_inst1_s2_sh;
  wire   [7:0] prince_inst_sbox_inst1_s1_sh;
  wire   [7:0] prince_inst_sbox_inst1_s0_sh;
  wire   [7:0] prince_inst_sbox_inst1_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst1_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst1_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst1_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst2_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst2_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst2_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst2_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst2_t3_sh;
  wire   [7:0] prince_inst_sbox_inst2_t2_sh;
  wire   [7:0] prince_inst_sbox_inst2_t1_sh;
  wire   [7:0] prince_inst_sbox_inst2_t0_sh;
  wire   [7:0] prince_inst_sbox_inst2_s3_sh;
  wire   [7:0] prince_inst_sbox_inst2_s2_sh;
  wire   [7:0] prince_inst_sbox_inst2_s1_sh;
  wire   [7:0] prince_inst_sbox_inst2_s0_sh;
  wire   [7:0] prince_inst_sbox_inst2_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst2_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst2_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst2_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst3_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst3_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst3_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst3_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst3_t3_sh;
  wire   [7:0] prince_inst_sbox_inst3_t2_sh;
  wire   [7:0] prince_inst_sbox_inst3_t1_sh;
  wire   [7:0] prince_inst_sbox_inst3_t0_sh;
  wire   [7:0] prince_inst_sbox_inst3_s3_sh;
  wire   [7:0] prince_inst_sbox_inst3_s2_sh;
  wire   [7:0] prince_inst_sbox_inst3_s1_sh;
  wire   [7:0] prince_inst_sbox_inst3_s0_sh;
  wire   [7:0] prince_inst_sbox_inst3_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst3_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst3_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst3_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst4_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst4_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst4_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst4_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst4_t3_sh;
  wire   [7:0] prince_inst_sbox_inst4_t2_sh;
  wire   [7:0] prince_inst_sbox_inst4_t1_sh;
  wire   [7:0] prince_inst_sbox_inst4_t0_sh;
  wire   [7:0] prince_inst_sbox_inst4_s3_sh;
  wire   [7:0] prince_inst_sbox_inst4_s2_sh;
  wire   [7:0] prince_inst_sbox_inst4_s1_sh;
  wire   [7:0] prince_inst_sbox_inst4_s0_sh;
  wire   [7:0] prince_inst_sbox_inst4_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst4_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst4_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst4_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst5_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst5_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst5_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst5_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst5_t3_sh;
  wire   [7:0] prince_inst_sbox_inst5_t2_sh;
  wire   [7:0] prince_inst_sbox_inst5_t1_sh;
  wire   [7:0] prince_inst_sbox_inst5_t0_sh;
  wire   [7:0] prince_inst_sbox_inst5_s3_sh;
  wire   [7:0] prince_inst_sbox_inst5_s2_sh;
  wire   [7:0] prince_inst_sbox_inst5_s1_sh;
  wire   [7:0] prince_inst_sbox_inst5_s0_sh;
  wire   [7:0] prince_inst_sbox_inst5_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst5_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst5_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst5_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst6_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst6_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst6_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst6_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst6_t3_sh;
  wire   [7:0] prince_inst_sbox_inst6_t2_sh;
  wire   [7:0] prince_inst_sbox_inst6_t1_sh;
  wire   [7:0] prince_inst_sbox_inst6_t0_sh;
  wire   [7:0] prince_inst_sbox_inst6_s3_sh;
  wire   [7:0] prince_inst_sbox_inst6_s2_sh;
  wire   [7:0] prince_inst_sbox_inst6_s1_sh;
  wire   [7:0] prince_inst_sbox_inst6_s0_sh;
  wire   [7:0] prince_inst_sbox_inst6_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst6_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst6_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst6_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst7_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst7_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst7_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst7_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst7_t3_sh;
  wire   [7:0] prince_inst_sbox_inst7_t2_sh;
  wire   [7:0] prince_inst_sbox_inst7_t1_sh;
  wire   [7:0] prince_inst_sbox_inst7_t0_sh;
  wire   [7:0] prince_inst_sbox_inst7_s3_sh;
  wire   [7:0] prince_inst_sbox_inst7_s2_sh;
  wire   [7:0] prince_inst_sbox_inst7_s1_sh;
  wire   [7:0] prince_inst_sbox_inst7_s0_sh;
  wire   [7:0] prince_inst_sbox_inst7_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst7_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst7_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst7_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst8_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst8_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst8_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst8_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst8_t3_sh;
  wire   [7:0] prince_inst_sbox_inst8_t2_sh;
  wire   [7:0] prince_inst_sbox_inst8_t1_sh;
  wire   [7:0] prince_inst_sbox_inst8_t0_sh;
  wire   [7:0] prince_inst_sbox_inst8_s3_sh;
  wire   [7:0] prince_inst_sbox_inst8_s2_sh;
  wire   [7:0] prince_inst_sbox_inst8_s1_sh;
  wire   [7:0] prince_inst_sbox_inst8_s0_sh;
  wire   [7:0] prince_inst_sbox_inst8_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst8_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst8_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst8_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst9_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst9_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst9_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst9_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst9_t3_sh;
  wire   [7:0] prince_inst_sbox_inst9_t2_sh;
  wire   [7:0] prince_inst_sbox_inst9_t1_sh;
  wire   [7:0] prince_inst_sbox_inst9_t0_sh;
  wire   [7:0] prince_inst_sbox_inst9_s3_sh;
  wire   [7:0] prince_inst_sbox_inst9_s2_sh;
  wire   [7:0] prince_inst_sbox_inst9_s1_sh;
  wire   [7:0] prince_inst_sbox_inst9_s0_sh;
  wire   [7:0] prince_inst_sbox_inst9_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst9_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst9_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst9_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst10_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst10_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst10_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst10_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst10_t3_sh;
  wire   [7:0] prince_inst_sbox_inst10_t2_sh;
  wire   [7:0] prince_inst_sbox_inst10_t1_sh;
  wire   [7:0] prince_inst_sbox_inst10_t0_sh;
  wire   [7:0] prince_inst_sbox_inst10_s3_sh;
  wire   [7:0] prince_inst_sbox_inst10_s2_sh;
  wire   [7:0] prince_inst_sbox_inst10_s1_sh;
  wire   [7:0] prince_inst_sbox_inst10_s0_sh;
  wire   [7:0] prince_inst_sbox_inst10_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst10_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst10_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst10_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst11_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst11_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst11_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst11_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst11_t3_sh;
  wire   [7:0] prince_inst_sbox_inst11_t2_sh;
  wire   [7:0] prince_inst_sbox_inst11_t1_sh;
  wire   [7:0] prince_inst_sbox_inst11_t0_sh;
  wire   [7:0] prince_inst_sbox_inst11_s3_sh;
  wire   [7:0] prince_inst_sbox_inst11_s2_sh;
  wire   [7:0] prince_inst_sbox_inst11_s1_sh;
  wire   [7:0] prince_inst_sbox_inst11_s0_sh;
  wire   [7:0] prince_inst_sbox_inst11_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst11_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst11_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst11_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst12_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst12_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst12_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst12_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst12_t3_sh;
  wire   [7:0] prince_inst_sbox_inst12_t2_sh;
  wire   [7:0] prince_inst_sbox_inst12_t1_sh;
  wire   [7:0] prince_inst_sbox_inst12_t0_sh;
  wire   [7:0] prince_inst_sbox_inst12_s3_sh;
  wire   [7:0] prince_inst_sbox_inst12_s2_sh;
  wire   [7:0] prince_inst_sbox_inst12_s1_sh;
  wire   [7:0] prince_inst_sbox_inst12_s0_sh;
  wire   [7:0] prince_inst_sbox_inst12_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst12_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst12_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst12_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst13_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst13_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst13_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst13_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst13_t3_sh;
  wire   [7:0] prince_inst_sbox_inst13_t2_sh;
  wire   [7:0] prince_inst_sbox_inst13_t1_sh;
  wire   [7:0] prince_inst_sbox_inst13_t0_sh;
  wire   [7:0] prince_inst_sbox_inst13_s3_sh;
  wire   [7:0] prince_inst_sbox_inst13_s2_sh;
  wire   [7:0] prince_inst_sbox_inst13_s1_sh;
  wire   [7:0] prince_inst_sbox_inst13_s0_sh;
  wire   [7:0] prince_inst_sbox_inst13_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst13_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst13_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst13_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst14_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst14_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst14_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst14_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst14_t3_sh;
  wire   [7:0] prince_inst_sbox_inst14_t2_sh;
  wire   [7:0] prince_inst_sbox_inst14_t1_sh;
  wire   [7:0] prince_inst_sbox_inst14_t0_sh;
  wire   [7:0] prince_inst_sbox_inst14_s3_sh;
  wire   [7:0] prince_inst_sbox_inst14_s2_sh;
  wire   [7:0] prince_inst_sbox_inst14_s1_sh;
  wire   [7:0] prince_inst_sbox_inst14_s0_sh;
  wire   [7:0] prince_inst_sbox_inst14_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst14_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst14_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst14_c_inst3_y;
  wire   [7:0] prince_inst_sbox_inst15_sh3_tmp;
  wire   [7:0] prince_inst_sbox_inst15_sh2_tmp;
  wire   [7:0] prince_inst_sbox_inst15_sh1_tmp;
  wire   [7:0] prince_inst_sbox_inst15_sh0_tmp;
  wire   [7:0] prince_inst_sbox_inst15_t3_sh;
  wire   [7:0] prince_inst_sbox_inst15_t2_sh;
  wire   [7:0] prince_inst_sbox_inst15_t1_sh;
  wire   [7:0] prince_inst_sbox_inst15_t0_sh;
  wire   [7:0] prince_inst_sbox_inst15_s3_sh;
  wire   [7:0] prince_inst_sbox_inst15_s2_sh;
  wire   [7:0] prince_inst_sbox_inst15_s1_sh;
  wire   [7:0] prince_inst_sbox_inst15_s0_sh;
  wire   [7:0] prince_inst_sbox_inst15_c_inst0_y;
  wire   [7:0] prince_inst_sbox_inst15_c_inst1_y;
  wire   [7:0] prince_inst_sbox_inst15_c_inst2_y;
  wire   [7:0] prince_inst_sbox_inst15_c_inst3_y;

  MUX2_X1 U773 ( .A(kext[73]), .B(kext[72]), .S(enc), .Z(n521) );
  XOR2_X1 U774 ( .A(p0_reg[9]), .B(n521), .Z(init_x[57]) );
  MUX2_X1 U775 ( .A(kext[72]), .B(kext[71]), .S(enc), .Z(n522) );
  XOR2_X1 U776 ( .A(p0_reg[8]), .B(n522), .Z(init_x[56]) );
  MUX2_X1 U777 ( .A(kext[71]), .B(kext[70]), .S(enc), .Z(n523) );
  XOR2_X1 U778 ( .A(p0_reg[7]), .B(n523), .Z(init_x[39]) );
  MUX2_X1 U779 ( .A(kext[70]), .B(kext[69]), .S(enc), .Z(n524) );
  XOR2_X1 U780 ( .A(p0_reg[6]), .B(n524), .Z(init_x[38]) );
  MUX2_X1 U781 ( .A(kext[127]), .B(kext[126]), .S(enc), .Z(n525) );
  XOR2_X1 U782 ( .A(p0_reg[63]), .B(n525), .Z(init_x[63]) );
  MUX2_X1 U783 ( .A(kext[126]), .B(kext[125]), .S(enc), .Z(n526) );
  XOR2_X1 U784 ( .A(p0_reg[62]), .B(n526), .Z(init_x[62]) );
  MUX2_X1 U785 ( .A(kext[125]), .B(kext[124]), .S(enc), .Z(n527) );
  XOR2_X1 U786 ( .A(p0_reg[61]), .B(n527), .Z(init_x[61]) );
  MUX2_X1 U787 ( .A(kext[124]), .B(kext[123]), .S(enc), .Z(n528) );
  XOR2_X1 U788 ( .A(p0_reg[60]), .B(n528), .Z(init_x[60]) );
  MUX2_X1 U789 ( .A(kext[69]), .B(kext[68]), .S(enc), .Z(n529) );
  XOR2_X1 U790 ( .A(p0_reg[5]), .B(n529), .Z(init_x[37]) );
  MUX2_X1 U791 ( .A(kext[123]), .B(kext[122]), .S(enc), .Z(n530) );
  XOR2_X1 U792 ( .A(p0_reg[59]), .B(n530), .Z(init_x[43]) );
  MUX2_X1 U793 ( .A(kext[122]), .B(kext[121]), .S(enc), .Z(n531) );
  XOR2_X1 U794 ( .A(p0_reg[58]), .B(n531), .Z(init_x[42]) );
  MUX2_X1 U795 ( .A(kext[121]), .B(kext[120]), .S(enc), .Z(n532) );
  XOR2_X1 U796 ( .A(p0_reg[57]), .B(n532), .Z(init_x[41]) );
  MUX2_X1 U797 ( .A(kext[120]), .B(kext[119]), .S(enc), .Z(n533) );
  XOR2_X1 U798 ( .A(p0_reg[56]), .B(n533), .Z(init_x[40]) );
  MUX2_X1 U799 ( .A(kext[119]), .B(kext[118]), .S(enc), .Z(n534) );
  XOR2_X1 U800 ( .A(p0_reg[55]), .B(n534), .Z(init_x[23]) );
  MUX2_X1 U801 ( .A(kext[118]), .B(kext[117]), .S(enc), .Z(n535) );
  XOR2_X1 U802 ( .A(p0_reg[54]), .B(n535), .Z(init_x[22]) );
  MUX2_X1 U803 ( .A(kext[117]), .B(kext[116]), .S(enc), .Z(n536) );
  XOR2_X1 U804 ( .A(p0_reg[53]), .B(n536), .Z(init_x[21]) );
  MUX2_X1 U805 ( .A(kext[116]), .B(kext[115]), .S(enc), .Z(n537) );
  XOR2_X1 U806 ( .A(p0_reg[52]), .B(n537), .Z(init_x[20]) );
  MUX2_X1 U807 ( .A(kext[115]), .B(kext[114]), .S(enc), .Z(n538) );
  XOR2_X1 U808 ( .A(p0_reg[51]), .B(n538), .Z(init_x[3]) );
  MUX2_X1 U809 ( .A(kext[114]), .B(kext[113]), .S(enc), .Z(n539) );
  XOR2_X1 U810 ( .A(p0_reg[50]), .B(n539), .Z(init_x[2]) );
  MUX2_X1 U811 ( .A(kext[68]), .B(kext[67]), .S(enc), .Z(n540) );
  XOR2_X1 U812 ( .A(p0_reg[4]), .B(n540), .Z(init_x[36]) );
  MUX2_X1 U813 ( .A(kext[113]), .B(kext[112]), .S(enc), .Z(n541) );
  XOR2_X1 U814 ( .A(p0_reg[49]), .B(n541), .Z(init_x[1]) );
  MUX2_X1 U815 ( .A(kext[112]), .B(kext[111]), .S(enc), .Z(n542) );
  XOR2_X1 U816 ( .A(p0_reg[48]), .B(n542), .Z(init_x[0]) );
  MUX2_X1 U817 ( .A(kext[111]), .B(kext[110]), .S(enc), .Z(n543) );
  XOR2_X1 U818 ( .A(p0_reg[47]), .B(n543), .Z(init_x[47]) );
  MUX2_X1 U819 ( .A(kext[110]), .B(kext[109]), .S(enc), .Z(n544) );
  XOR2_X1 U820 ( .A(p0_reg[46]), .B(n544), .Z(init_x[46]) );
  MUX2_X1 U821 ( .A(kext[109]), .B(kext[108]), .S(enc), .Z(n545) );
  XOR2_X1 U822 ( .A(p0_reg[45]), .B(n545), .Z(init_x[45]) );
  MUX2_X1 U823 ( .A(kext[108]), .B(kext[107]), .S(enc), .Z(n546) );
  XOR2_X1 U824 ( .A(p0_reg[44]), .B(n546), .Z(init_x[44]) );
  MUX2_X1 U825 ( .A(kext[107]), .B(kext[106]), .S(enc), .Z(n547) );
  XOR2_X1 U826 ( .A(p0_reg[43]), .B(n547), .Z(init_x[27]) );
  MUX2_X1 U827 ( .A(kext[106]), .B(kext[105]), .S(enc), .Z(n548) );
  XOR2_X1 U828 ( .A(p0_reg[42]), .B(n548), .Z(init_x[26]) );
  MUX2_X1 U829 ( .A(kext[105]), .B(kext[104]), .S(enc), .Z(n549) );
  XOR2_X1 U830 ( .A(p0_reg[41]), .B(n549), .Z(init_x[25]) );
  MUX2_X1 U831 ( .A(kext[104]), .B(kext[103]), .S(enc), .Z(n550) );
  XOR2_X1 U832 ( .A(p0_reg[40]), .B(n550), .Z(init_x[24]) );
  MUX2_X1 U833 ( .A(kext[67]), .B(kext[66]), .S(enc), .Z(n551) );
  XOR2_X1 U834 ( .A(p0_reg[3]), .B(n551), .Z(init_x[19]) );
  MUX2_X1 U835 ( .A(kext[103]), .B(kext[102]), .S(enc), .Z(n552) );
  XOR2_X1 U836 ( .A(p0_reg[39]), .B(n552), .Z(init_x[7]) );
  MUX2_X1 U837 ( .A(kext[102]), .B(kext[101]), .S(enc), .Z(n553) );
  XOR2_X1 U838 ( .A(p0_reg[38]), .B(n553), .Z(init_x[6]) );
  MUX2_X1 U839 ( .A(kext[101]), .B(kext[100]), .S(enc), .Z(n554) );
  XOR2_X1 U840 ( .A(p0_reg[37]), .B(n554), .Z(init_x[5]) );
  MUX2_X1 U841 ( .A(kext[100]), .B(kext[99]), .S(enc), .Z(n555) );
  XOR2_X1 U842 ( .A(p0_reg[36]), .B(n555), .Z(init_x[4]) );
  MUX2_X1 U843 ( .A(kext[99]), .B(kext[98]), .S(enc), .Z(n556) );
  XOR2_X1 U844 ( .A(p0_reg[35]), .B(n556), .Z(init_x[51]) );
  MUX2_X1 U845 ( .A(kext[98]), .B(kext[97]), .S(enc), .Z(n557) );
  XOR2_X1 U846 ( .A(p0_reg[34]), .B(n557), .Z(init_x[50]) );
  MUX2_X1 U847 ( .A(kext[97]), .B(kext[96]), .S(enc), .Z(n558) );
  XOR2_X1 U848 ( .A(p0_reg[33]), .B(n558), .Z(init_x[49]) );
  MUX2_X1 U849 ( .A(kext[96]), .B(kext[95]), .S(enc), .Z(n559) );
  XOR2_X1 U850 ( .A(p0_reg[32]), .B(n559), .Z(init_x[48]) );
  MUX2_X1 U851 ( .A(kext[95]), .B(kext[94]), .S(enc), .Z(n560) );
  XOR2_X1 U852 ( .A(p0_reg[31]), .B(n560), .Z(init_x[31]) );
  MUX2_X1 U853 ( .A(kext[94]), .B(kext[93]), .S(enc), .Z(n561) );
  XOR2_X1 U854 ( .A(p0_reg[30]), .B(n561), .Z(init_x[30]) );
  MUX2_X1 U855 ( .A(kext[66]), .B(kext[65]), .S(enc), .Z(n562) );
  XOR2_X1 U856 ( .A(p0_reg[2]), .B(n562), .Z(init_x[18]) );
  MUX2_X1 U857 ( .A(kext[93]), .B(kext[92]), .S(enc), .Z(n563) );
  XOR2_X1 U858 ( .A(p0_reg[29]), .B(n563), .Z(init_x[29]) );
  MUX2_X1 U859 ( .A(kext[92]), .B(kext[91]), .S(enc), .Z(n564) );
  XOR2_X1 U860 ( .A(p0_reg[28]), .B(n564), .Z(init_x[28]) );
  MUX2_X1 U861 ( .A(kext[91]), .B(kext[90]), .S(enc), .Z(n565) );
  XOR2_X1 U862 ( .A(p0_reg[27]), .B(n565), .Z(init_x[11]) );
  MUX2_X1 U863 ( .A(kext[90]), .B(kext[89]), .S(enc), .Z(n566) );
  XOR2_X1 U864 ( .A(p0_reg[26]), .B(n566), .Z(init_x[10]) );
  MUX2_X1 U865 ( .A(kext[89]), .B(kext[88]), .S(enc), .Z(n567) );
  XOR2_X1 U866 ( .A(p0_reg[25]), .B(n567), .Z(init_x[9]) );
  MUX2_X1 U867 ( .A(kext[88]), .B(kext[87]), .S(enc), .Z(n568) );
  XOR2_X1 U868 ( .A(p0_reg[24]), .B(n568), .Z(init_x[8]) );
  MUX2_X1 U869 ( .A(kext[87]), .B(kext[86]), .S(enc), .Z(n569) );
  XOR2_X1 U870 ( .A(p0_reg[23]), .B(n569), .Z(init_x[55]) );
  MUX2_X1 U871 ( .A(kext[86]), .B(kext[85]), .S(enc), .Z(n570) );
  XOR2_X1 U872 ( .A(p0_reg[22]), .B(n570), .Z(init_x[54]) );
  MUX2_X1 U873 ( .A(kext[85]), .B(kext[84]), .S(enc), .Z(n571) );
  XOR2_X1 U874 ( .A(p0_reg[21]), .B(n571), .Z(init_x[53]) );
  MUX2_X1 U875 ( .A(kext[84]), .B(kext[83]), .S(enc), .Z(n572) );
  XOR2_X1 U876 ( .A(p0_reg[20]), .B(n572), .Z(init_x[52]) );
  MUX2_X1 U877 ( .A(kext[65]), .B(kext[1]), .S(enc), .Z(n573) );
  XOR2_X1 U878 ( .A(p0_reg[1]), .B(n573), .Z(init_x[17]) );
  MUX2_X1 U879 ( .A(kext[83]), .B(kext[82]), .S(enc), .Z(n574) );
  XOR2_X1 U880 ( .A(p0_reg[19]), .B(n574), .Z(init_x[35]) );
  MUX2_X1 U881 ( .A(kext[82]), .B(kext[81]), .S(enc), .Z(n575) );
  XOR2_X1 U882 ( .A(p0_reg[18]), .B(n575), .Z(init_x[34]) );
  MUX2_X1 U883 ( .A(kext[81]), .B(kext[80]), .S(enc), .Z(n576) );
  XOR2_X1 U884 ( .A(p0_reg[17]), .B(n576), .Z(init_x[33]) );
  MUX2_X1 U885 ( .A(kext[80]), .B(kext[79]), .S(enc), .Z(n577) );
  XOR2_X1 U886 ( .A(p0_reg[16]), .B(n577), .Z(init_x[32]) );
  MUX2_X1 U887 ( .A(kext[79]), .B(kext[78]), .S(enc), .Z(n578) );
  XOR2_X1 U888 ( .A(p0_reg[15]), .B(n578), .Z(init_x[15]) );
  MUX2_X1 U889 ( .A(kext[78]), .B(kext[77]), .S(enc), .Z(n579) );
  XOR2_X1 U890 ( .A(p0_reg[14]), .B(n579), .Z(init_x[14]) );
  MUX2_X1 U891 ( .A(kext[77]), .B(kext[76]), .S(enc), .Z(n580) );
  XOR2_X1 U892 ( .A(p0_reg[13]), .B(n580), .Z(init_x[13]) );
  MUX2_X1 U893 ( .A(kext[76]), .B(kext[75]), .S(enc), .Z(n581) );
  XOR2_X1 U894 ( .A(p0_reg[12]), .B(n581), .Z(init_x[12]) );
  MUX2_X1 U895 ( .A(kext[75]), .B(kext[74]), .S(enc), .Z(n582) );
  XOR2_X1 U896 ( .A(p0_reg[11]), .B(n582), .Z(init_x[59]) );
  MUX2_X1 U897 ( .A(kext[74]), .B(kext[73]), .S(enc), .Z(n583) );
  XOR2_X1 U898 ( .A(p0_reg[10]), .B(n583), .Z(init_x[58]) );
  MUX2_X1 U899 ( .A(kext[64]), .B(kext[127]), .S(enc), .Z(n584) );
  XOR2_X1 U900 ( .A(p0_reg[0]), .B(n584), .Z(init_x[16]) );
  MUX2_X1 U901 ( .A(kext[72]), .B(kext[73]), .S(enc), .Z(n585) );
  XOR2_X1 U902 ( .A(final_x[9]), .B(n585), .Z(final_x_k[9]) );
  MUX2_X1 U903 ( .A(kext[71]), .B(kext[72]), .S(enc), .Z(n586) );
  XOR2_X1 U904 ( .A(final_x[8]), .B(n586), .Z(final_x_k[8]) );
  MUX2_X1 U905 ( .A(kext[70]), .B(kext[71]), .S(enc), .Z(n587) );
  XOR2_X1 U906 ( .A(final_x[7]), .B(n587), .Z(final_x_k[7]) );
  MUX2_X1 U907 ( .A(kext[69]), .B(kext[70]), .S(enc), .Z(n588) );
  XOR2_X1 U908 ( .A(final_x[6]), .B(n588), .Z(final_x_k[6]) );
  MUX2_X1 U909 ( .A(kext[126]), .B(kext[127]), .S(enc), .Z(n589) );
  XOR2_X1 U910 ( .A(final_x[63]), .B(n589), .Z(final_x_k[63]) );
  MUX2_X1 U911 ( .A(kext[125]), .B(kext[126]), .S(enc), .Z(n590) );
  XOR2_X1 U912 ( .A(final_x[62]), .B(n590), .Z(final_x_k[62]) );
  MUX2_X1 U913 ( .A(kext[124]), .B(kext[125]), .S(enc), .Z(n591) );
  XOR2_X1 U914 ( .A(final_x[61]), .B(n591), .Z(final_x_k[61]) );
  MUX2_X1 U915 ( .A(kext[123]), .B(kext[124]), .S(enc), .Z(n592) );
  XOR2_X1 U916 ( .A(final_x[60]), .B(n592), .Z(final_x_k[60]) );
  MUX2_X1 U917 ( .A(kext[68]), .B(kext[69]), .S(enc), .Z(n593) );
  XOR2_X1 U918 ( .A(final_x[5]), .B(n593), .Z(final_x_k[5]) );
  MUX2_X1 U919 ( .A(kext[122]), .B(kext[123]), .S(enc), .Z(n594) );
  XOR2_X1 U920 ( .A(final_x[59]), .B(n594), .Z(final_x_k[59]) );
  MUX2_X1 U921 ( .A(kext[121]), .B(kext[122]), .S(enc), .Z(n595) );
  XOR2_X1 U922 ( .A(final_x[58]), .B(n595), .Z(final_x_k[58]) );
  MUX2_X1 U923 ( .A(kext[120]), .B(kext[121]), .S(enc), .Z(n596) );
  XOR2_X1 U924 ( .A(final_x[57]), .B(n596), .Z(final_x_k[57]) );
  MUX2_X1 U925 ( .A(kext[119]), .B(kext[120]), .S(enc), .Z(n597) );
  XOR2_X1 U926 ( .A(final_x[56]), .B(n597), .Z(final_x_k[56]) );
  MUX2_X1 U927 ( .A(kext[118]), .B(kext[119]), .S(enc), .Z(n598) );
  XOR2_X1 U928 ( .A(final_x[55]), .B(n598), .Z(final_x_k[55]) );
  MUX2_X1 U929 ( .A(kext[117]), .B(kext[118]), .S(enc), .Z(n599) );
  XOR2_X1 U930 ( .A(final_x[54]), .B(n599), .Z(final_x_k[54]) );
  MUX2_X1 U931 ( .A(kext[116]), .B(kext[117]), .S(enc), .Z(n600) );
  XOR2_X1 U932 ( .A(final_x[53]), .B(n600), .Z(final_x_k[53]) );
  MUX2_X1 U933 ( .A(kext[115]), .B(kext[116]), .S(enc), .Z(n601) );
  XOR2_X1 U934 ( .A(final_x[52]), .B(n601), .Z(final_x_k[52]) );
  MUX2_X1 U935 ( .A(kext[114]), .B(kext[115]), .S(enc), .Z(n602) );
  XOR2_X1 U936 ( .A(final_x[51]), .B(n602), .Z(final_x_k[51]) );
  MUX2_X1 U937 ( .A(kext[113]), .B(kext[114]), .S(enc), .Z(n603) );
  XOR2_X1 U938 ( .A(final_x[50]), .B(n603), .Z(final_x_k[50]) );
  MUX2_X1 U939 ( .A(kext[67]), .B(kext[68]), .S(enc), .Z(n604) );
  XOR2_X1 U940 ( .A(final_x[4]), .B(n604), .Z(final_x_k[4]) );
  MUX2_X1 U941 ( .A(kext[112]), .B(kext[113]), .S(enc), .Z(n605) );
  XOR2_X1 U942 ( .A(final_x[49]), .B(n605), .Z(final_x_k[49]) );
  MUX2_X1 U943 ( .A(kext[111]), .B(kext[112]), .S(enc), .Z(n606) );
  XOR2_X1 U944 ( .A(final_x[48]), .B(n606), .Z(final_x_k[48]) );
  MUX2_X1 U945 ( .A(kext[110]), .B(kext[111]), .S(enc), .Z(n607) );
  XOR2_X1 U946 ( .A(final_x[47]), .B(n607), .Z(final_x_k[47]) );
  MUX2_X1 U947 ( .A(kext[109]), .B(kext[110]), .S(enc), .Z(n608) );
  XOR2_X1 U948 ( .A(final_x[46]), .B(n608), .Z(final_x_k[46]) );
  MUX2_X1 U949 ( .A(kext[108]), .B(kext[109]), .S(enc), .Z(n609) );
  XOR2_X1 U950 ( .A(final_x[45]), .B(n609), .Z(final_x_k[45]) );
  MUX2_X1 U951 ( .A(kext[107]), .B(kext[108]), .S(enc), .Z(n610) );
  XOR2_X1 U952 ( .A(final_x[44]), .B(n610), .Z(final_x_k[44]) );
  MUX2_X1 U953 ( .A(kext[106]), .B(kext[107]), .S(enc), .Z(n611) );
  XOR2_X1 U954 ( .A(final_x[43]), .B(n611), .Z(final_x_k[43]) );
  MUX2_X1 U955 ( .A(kext[105]), .B(kext[106]), .S(enc), .Z(n612) );
  XOR2_X1 U956 ( .A(final_x[42]), .B(n612), .Z(final_x_k[42]) );
  MUX2_X1 U957 ( .A(kext[104]), .B(kext[105]), .S(enc), .Z(n613) );
  XOR2_X1 U958 ( .A(final_x[41]), .B(n613), .Z(final_x_k[41]) );
  MUX2_X1 U959 ( .A(kext[103]), .B(kext[104]), .S(enc), .Z(n614) );
  XOR2_X1 U960 ( .A(final_x[40]), .B(n614), .Z(final_x_k[40]) );
  MUX2_X1 U961 ( .A(kext[66]), .B(kext[67]), .S(enc), .Z(n615) );
  XOR2_X1 U962 ( .A(final_x[3]), .B(n615), .Z(final_x_k[3]) );
  MUX2_X1 U963 ( .A(kext[102]), .B(kext[103]), .S(enc), .Z(n616) );
  XOR2_X1 U964 ( .A(final_x[39]), .B(n616), .Z(final_x_k[39]) );
  MUX2_X1 U965 ( .A(kext[101]), .B(kext[102]), .S(enc), .Z(n617) );
  XOR2_X1 U966 ( .A(final_x[38]), .B(n617), .Z(final_x_k[38]) );
  MUX2_X1 U967 ( .A(kext[100]), .B(kext[101]), .S(enc), .Z(n618) );
  XOR2_X1 U968 ( .A(final_x[37]), .B(n618), .Z(final_x_k[37]) );
  MUX2_X1 U969 ( .A(kext[99]), .B(kext[100]), .S(enc), .Z(n619) );
  XOR2_X1 U970 ( .A(final_x[36]), .B(n619), .Z(final_x_k[36]) );
  MUX2_X1 U971 ( .A(kext[98]), .B(kext[99]), .S(enc), .Z(n620) );
  XOR2_X1 U972 ( .A(final_x[35]), .B(n620), .Z(final_x_k[35]) );
  MUX2_X1 U973 ( .A(kext[97]), .B(kext[98]), .S(enc), .Z(n621) );
  XOR2_X1 U974 ( .A(final_x[34]), .B(n621), .Z(final_x_k[34]) );
  MUX2_X1 U975 ( .A(kext[96]), .B(kext[97]), .S(enc), .Z(n622) );
  XOR2_X1 U976 ( .A(final_x[33]), .B(n622), .Z(final_x_k[33]) );
  MUX2_X1 U977 ( .A(kext[95]), .B(kext[96]), .S(enc), .Z(n623) );
  XOR2_X1 U978 ( .A(final_x[32]), .B(n623), .Z(final_x_k[32]) );
  MUX2_X1 U979 ( .A(kext[94]), .B(kext[95]), .S(enc), .Z(n624) );
  XOR2_X1 U980 ( .A(final_x[31]), .B(n624), .Z(final_x_k[31]) );
  MUX2_X1 U981 ( .A(kext[93]), .B(kext[94]), .S(enc), .Z(n625) );
  XOR2_X1 U982 ( .A(final_x[30]), .B(n625), .Z(final_x_k[30]) );
  MUX2_X1 U983 ( .A(kext[65]), .B(kext[66]), .S(enc), .Z(n626) );
  XOR2_X1 U984 ( .A(final_x[2]), .B(n626), .Z(final_x_k[2]) );
  MUX2_X1 U985 ( .A(kext[92]), .B(kext[93]), .S(enc), .Z(n627) );
  XOR2_X1 U986 ( .A(final_x[29]), .B(n627), .Z(final_x_k[29]) );
  MUX2_X1 U987 ( .A(kext[91]), .B(kext[92]), .S(enc), .Z(n628) );
  XOR2_X1 U988 ( .A(final_x[28]), .B(n628), .Z(final_x_k[28]) );
  MUX2_X1 U989 ( .A(kext[90]), .B(kext[91]), .S(enc), .Z(n629) );
  XOR2_X1 U990 ( .A(final_x[27]), .B(n629), .Z(final_x_k[27]) );
  MUX2_X1 U991 ( .A(kext[89]), .B(kext[90]), .S(enc), .Z(n630) );
  XOR2_X1 U992 ( .A(final_x[26]), .B(n630), .Z(final_x_k[26]) );
  MUX2_X1 U993 ( .A(kext[88]), .B(kext[89]), .S(enc), .Z(n631) );
  XOR2_X1 U994 ( .A(final_x[25]), .B(n631), .Z(final_x_k[25]) );
  MUX2_X1 U995 ( .A(kext[87]), .B(kext[88]), .S(enc), .Z(n632) );
  XOR2_X1 U996 ( .A(final_x[24]), .B(n632), .Z(final_x_k[24]) );
  MUX2_X1 U997 ( .A(kext[86]), .B(kext[87]), .S(enc), .Z(n633) );
  XOR2_X1 U998 ( .A(final_x[23]), .B(n633), .Z(final_x_k[23]) );
  MUX2_X1 U999 ( .A(kext[85]), .B(kext[86]), .S(enc), .Z(n634) );
  XOR2_X1 U1000 ( .A(final_x[22]), .B(n634), .Z(final_x_k[22]) );
  MUX2_X1 U1001 ( .A(kext[84]), .B(kext[85]), .S(enc), .Z(n635) );
  XOR2_X1 U1002 ( .A(final_x[21]), .B(n635), .Z(final_x_k[21]) );
  MUX2_X1 U1003 ( .A(kext[83]), .B(kext[84]), .S(enc), .Z(n636) );
  XOR2_X1 U1004 ( .A(final_x[20]), .B(n636), .Z(final_x_k[20]) );
  MUX2_X1 U1005 ( .A(kext[1]), .B(kext[65]), .S(enc), .Z(n637) );
  XOR2_X1 U1006 ( .A(final_x[1]), .B(n637), .Z(final_x_k[1]) );
  MUX2_X1 U1007 ( .A(kext[82]), .B(kext[83]), .S(enc), .Z(n638) );
  XOR2_X1 U1008 ( .A(final_x[19]), .B(n638), .Z(final_x_k[19]) );
  MUX2_X1 U1009 ( .A(kext[81]), .B(kext[82]), .S(enc), .Z(n639) );
  XOR2_X1 U1010 ( .A(final_x[18]), .B(n639), .Z(final_x_k[18]) );
  MUX2_X1 U1011 ( .A(kext[80]), .B(kext[81]), .S(enc), .Z(n640) );
  XOR2_X1 U1012 ( .A(final_x[17]), .B(n640), .Z(final_x_k[17]) );
  MUX2_X1 U1013 ( .A(kext[79]), .B(kext[80]), .S(enc), .Z(n641) );
  XOR2_X1 U1014 ( .A(final_x[16]), .B(n641), .Z(final_x_k[16]) );
  MUX2_X1 U1015 ( .A(kext[78]), .B(kext[79]), .S(enc), .Z(n642) );
  XOR2_X1 U1016 ( .A(final_x[15]), .B(n642), .Z(final_x_k[15]) );
  MUX2_X1 U1017 ( .A(kext[77]), .B(kext[78]), .S(enc), .Z(n643) );
  XOR2_X1 U1018 ( .A(final_x[14]), .B(n643), .Z(final_x_k[14]) );
  MUX2_X1 U1019 ( .A(kext[76]), .B(kext[77]), .S(enc), .Z(n644) );
  XOR2_X1 U1020 ( .A(final_x[13]), .B(n644), .Z(final_x_k[13]) );
  MUX2_X1 U1021 ( .A(kext[75]), .B(kext[76]), .S(enc), .Z(n645) );
  XOR2_X1 U1022 ( .A(final_x[12]), .B(n645), .Z(final_x_k[12]) );
  MUX2_X1 U1023 ( .A(kext[74]), .B(kext[75]), .S(enc), .Z(n646) );
  XOR2_X1 U1024 ( .A(final_x[11]), .B(n646), .Z(final_x_k[11]) );
  MUX2_X1 U1025 ( .A(kext[73]), .B(kext[74]), .S(enc), .Z(n647) );
  XOR2_X1 U1026 ( .A(final_x[10]), .B(n647), .Z(final_x_k[10]) );
  MUX2_X1 U1027 ( .A(kext[127]), .B(kext[64]), .S(enc), .Z(n648) );
  XOR2_X1 U1028 ( .A(final_x[0]), .B(n648), .Z(final_x_k[0]) );
  XOR2_X1 k_inst_U1 ( .A(kext[1]), .B(kext[126]), .Z(kext[64]) );
  NAND2_X1 reg_k0_U205 ( .A1(reg_k0_n340), .A2(reg_k0_n339), .ZN(reg_k0_n195)
         );
  NAND2_X1 reg_k0_U204 ( .A1(k[63]), .A2(reg_k0_n338), .ZN(reg_k0_n339) );
  NAND2_X1 reg_k0_U203 ( .A1(kext[191]), .A2(reg_k0_n337), .ZN(reg_k0_n340) );
  NAND2_X1 reg_k0_U202 ( .A1(reg_k0_n336), .A2(reg_k0_n335), .ZN(reg_k0_n194)
         );
  NAND2_X1 reg_k0_U201 ( .A1(k[62]), .A2(reg_k0_n338), .ZN(reg_k0_n335) );
  NAND2_X1 reg_k0_U200 ( .A1(kext[190]), .A2(reg_k0_n337), .ZN(reg_k0_n336) );
  NAND2_X1 reg_k0_U199 ( .A1(reg_k0_n334), .A2(reg_k0_n333), .ZN(reg_k0_n193)
         );
  NAND2_X1 reg_k0_U198 ( .A1(k[61]), .A2(reg_k0_n338), .ZN(reg_k0_n333) );
  NAND2_X1 reg_k0_U197 ( .A1(kext[189]), .A2(reg_k0_n337), .ZN(reg_k0_n334) );
  NAND2_X1 reg_k0_U196 ( .A1(reg_k0_n332), .A2(reg_k0_n331), .ZN(reg_k0_n192)
         );
  NAND2_X1 reg_k0_U195 ( .A1(k[60]), .A2(reg_k0_n338), .ZN(reg_k0_n331) );
  NAND2_X1 reg_k0_U194 ( .A1(kext[188]), .A2(reg_k0_n337), .ZN(reg_k0_n332) );
  NAND2_X1 reg_k0_U193 ( .A1(reg_k0_n330), .A2(reg_k0_n329), .ZN(reg_k0_n167)
         );
  NAND2_X1 reg_k0_U192 ( .A1(k[35]), .A2(reg_k0_n338), .ZN(reg_k0_n329) );
  NAND2_X1 reg_k0_U191 ( .A1(kext[163]), .A2(reg_k0_n337), .ZN(reg_k0_n330) );
  NAND2_X1 reg_k0_U190 ( .A1(reg_k0_n328), .A2(reg_k0_n327), .ZN(reg_k0_n166)
         );
  NAND2_X1 reg_k0_U189 ( .A1(k[34]), .A2(reg_k0_n338), .ZN(reg_k0_n327) );
  NAND2_X1 reg_k0_U188 ( .A1(kext[162]), .A2(reg_k0_n337), .ZN(reg_k0_n328) );
  NAND2_X1 reg_k0_U187 ( .A1(reg_k0_n326), .A2(reg_k0_n325), .ZN(reg_k0_n165)
         );
  NAND2_X1 reg_k0_U186 ( .A1(k[33]), .A2(reg_k0_n338), .ZN(reg_k0_n325) );
  NAND2_X1 reg_k0_U185 ( .A1(kext[161]), .A2(reg_k0_n337), .ZN(reg_k0_n326) );
  NAND2_X1 reg_k0_U184 ( .A1(reg_k0_n324), .A2(reg_k0_n323), .ZN(reg_k0_n164)
         );
  NAND2_X1 reg_k0_U183 ( .A1(k[32]), .A2(reg_k0_n338), .ZN(reg_k0_n323) );
  NAND2_X1 reg_k0_U182 ( .A1(kext[160]), .A2(reg_k0_n337), .ZN(reg_k0_n324) );
  NAND2_X1 reg_k0_U181 ( .A1(reg_k0_n322), .A2(reg_k0_n321), .ZN(reg_k0_n163)
         );
  NAND2_X1 reg_k0_U180 ( .A1(k[31]), .A2(reg_k0_n338), .ZN(reg_k0_n321) );
  NAND2_X1 reg_k0_U179 ( .A1(kext[159]), .A2(reg_k0_n337), .ZN(reg_k0_n322) );
  NAND2_X1 reg_k0_U178 ( .A1(reg_k0_n320), .A2(reg_k0_n319), .ZN(reg_k0_n162)
         );
  NAND2_X1 reg_k0_U177 ( .A1(k[30]), .A2(reg_k0_n338), .ZN(reg_k0_n319) );
  NAND2_X1 reg_k0_U176 ( .A1(kext[158]), .A2(reg_k0_n337), .ZN(reg_k0_n320) );
  NAND2_X1 reg_k0_U175 ( .A1(reg_k0_n318), .A2(reg_k0_n317), .ZN(reg_k0_n161)
         );
  NAND2_X1 reg_k0_U174 ( .A1(k[29]), .A2(reg_k0_n338), .ZN(reg_k0_n317) );
  NAND2_X1 reg_k0_U173 ( .A1(kext[157]), .A2(reg_k0_n337), .ZN(reg_k0_n318) );
  NAND2_X1 reg_k0_U172 ( .A1(reg_k0_n316), .A2(reg_k0_n315), .ZN(reg_k0_n160)
         );
  NAND2_X1 reg_k0_U171 ( .A1(k[28]), .A2(reg_k0_n338), .ZN(reg_k0_n315) );
  NAND2_X1 reg_k0_U170 ( .A1(kext[156]), .A2(reg_k0_n337), .ZN(reg_k0_n316) );
  NAND2_X1 reg_k0_U169 ( .A1(reg_k0_n314), .A2(reg_k0_n313), .ZN(reg_k0_n159)
         );
  NAND2_X1 reg_k0_U168 ( .A1(k[27]), .A2(reg_k0_n312), .ZN(reg_k0_n313) );
  NAND2_X1 reg_k0_U167 ( .A1(kext[155]), .A2(reg_k0_n311), .ZN(reg_k0_n314) );
  NAND2_X1 reg_k0_U166 ( .A1(reg_k0_n310), .A2(reg_k0_n309), .ZN(reg_k0_n158)
         );
  NAND2_X1 reg_k0_U165 ( .A1(k[26]), .A2(reg_k0_n312), .ZN(reg_k0_n309) );
  NAND2_X1 reg_k0_U164 ( .A1(kext[154]), .A2(reg_k0_n311), .ZN(reg_k0_n310) );
  NAND2_X1 reg_k0_U163 ( .A1(reg_k0_n308), .A2(reg_k0_n307), .ZN(reg_k0_n157)
         );
  NAND2_X1 reg_k0_U162 ( .A1(k[25]), .A2(reg_k0_n312), .ZN(reg_k0_n307) );
  NAND2_X1 reg_k0_U161 ( .A1(kext[153]), .A2(reg_k0_n311), .ZN(reg_k0_n308) );
  NAND2_X1 reg_k0_U160 ( .A1(reg_k0_n306), .A2(reg_k0_n305), .ZN(reg_k0_n156)
         );
  NAND2_X1 reg_k0_U159 ( .A1(k[24]), .A2(reg_k0_n312), .ZN(reg_k0_n305) );
  NAND2_X1 reg_k0_U158 ( .A1(kext[152]), .A2(reg_k0_n311), .ZN(reg_k0_n306) );
  NAND2_X1 reg_k0_U157 ( .A1(reg_k0_n304), .A2(reg_k0_n303), .ZN(reg_k0_n155)
         );
  NAND2_X1 reg_k0_U156 ( .A1(k[23]), .A2(reg_k0_n312), .ZN(reg_k0_n303) );
  NAND2_X1 reg_k0_U155 ( .A1(kext[151]), .A2(reg_k0_n311), .ZN(reg_k0_n304) );
  NAND2_X1 reg_k0_U154 ( .A1(reg_k0_n302), .A2(reg_k0_n301), .ZN(reg_k0_n154)
         );
  NAND2_X1 reg_k0_U153 ( .A1(k[22]), .A2(reg_k0_n312), .ZN(reg_k0_n301) );
  NAND2_X1 reg_k0_U152 ( .A1(kext[150]), .A2(reg_k0_n311), .ZN(reg_k0_n302) );
  NAND2_X1 reg_k0_U151 ( .A1(reg_k0_n300), .A2(reg_k0_n299), .ZN(reg_k0_n153)
         );
  NAND2_X1 reg_k0_U150 ( .A1(k[21]), .A2(reg_k0_n312), .ZN(reg_k0_n299) );
  NAND2_X1 reg_k0_U149 ( .A1(kext[149]), .A2(reg_k0_n311), .ZN(reg_k0_n300) );
  NAND2_X1 reg_k0_U148 ( .A1(reg_k0_n298), .A2(reg_k0_n297), .ZN(reg_k0_n152)
         );
  NAND2_X1 reg_k0_U147 ( .A1(k[20]), .A2(reg_k0_n312), .ZN(reg_k0_n297) );
  NAND2_X1 reg_k0_U146 ( .A1(kext[148]), .A2(reg_k0_n311), .ZN(reg_k0_n298) );
  NAND2_X1 reg_k0_U145 ( .A1(reg_k0_n296), .A2(reg_k0_n295), .ZN(reg_k0_n151)
         );
  NAND2_X1 reg_k0_U144 ( .A1(k[19]), .A2(reg_k0_n312), .ZN(reg_k0_n295) );
  NAND2_X1 reg_k0_U143 ( .A1(kext[147]), .A2(reg_k0_n311), .ZN(reg_k0_n296) );
  NAND2_X1 reg_k0_U142 ( .A1(reg_k0_n294), .A2(reg_k0_n293), .ZN(reg_k0_n150)
         );
  NAND2_X1 reg_k0_U141 ( .A1(k[18]), .A2(reg_k0_n312), .ZN(reg_k0_n293) );
  NAND2_X1 reg_k0_U140 ( .A1(kext[146]), .A2(reg_k0_n311), .ZN(reg_k0_n294) );
  NAND2_X1 reg_k0_U139 ( .A1(reg_k0_n292), .A2(reg_k0_n291), .ZN(reg_k0_n149)
         );
  NAND2_X1 reg_k0_U138 ( .A1(k[17]), .A2(reg_k0_n312), .ZN(reg_k0_n291) );
  NAND2_X1 reg_k0_U137 ( .A1(kext[145]), .A2(reg_k0_n311), .ZN(reg_k0_n292) );
  NAND2_X1 reg_k0_U136 ( .A1(reg_k0_n290), .A2(reg_k0_n289), .ZN(reg_k0_n148)
         );
  NAND2_X1 reg_k0_U135 ( .A1(k[16]), .A2(reg_k0_n312), .ZN(reg_k0_n289) );
  NAND2_X1 reg_k0_U134 ( .A1(kext[144]), .A2(reg_k0_n311), .ZN(reg_k0_n290) );
  NAND2_X1 reg_k0_U133 ( .A1(reg_k0_n288), .A2(reg_k0_n287), .ZN(reg_k0_n147)
         );
  NAND2_X1 reg_k0_U132 ( .A1(k[15]), .A2(reg_k0_n312), .ZN(reg_k0_n287) );
  NAND2_X1 reg_k0_U131 ( .A1(prince_inst_rc2_inv[15]), .A2(reg_k0_n311), .ZN(
        reg_k0_n288) );
  NAND2_X1 reg_k0_U130 ( .A1(reg_k0_n286), .A2(reg_k0_n285), .ZN(reg_k0_n146)
         );
  NAND2_X1 reg_k0_U129 ( .A1(k[14]), .A2(reg_k0_n338), .ZN(reg_k0_n285) );
  NAND2_X1 reg_k0_U128 ( .A1(kext[142]), .A2(reg_k0_n337), .ZN(reg_k0_n286) );
  NAND2_X1 reg_k0_U127 ( .A1(reg_k0_n284), .A2(reg_k0_n283), .ZN(reg_k0_n145)
         );
  NAND2_X1 reg_k0_U126 ( .A1(k[13]), .A2(reg_k0_n312), .ZN(reg_k0_n283) );
  NAND2_X1 reg_k0_U125 ( .A1(kext[141]), .A2(reg_k0_n311), .ZN(reg_k0_n284) );
  NAND2_X1 reg_k0_U124 ( .A1(reg_k0_n282), .A2(reg_k0_n281), .ZN(reg_k0_n144)
         );
  NAND2_X1 reg_k0_U123 ( .A1(k[12]), .A2(reg_k0_n338), .ZN(reg_k0_n281) );
  NAND2_X1 reg_k0_U122 ( .A1(kext[140]), .A2(reg_k0_n337), .ZN(reg_k0_n282) );
  NAND2_X1 reg_k0_U121 ( .A1(reg_k0_n280), .A2(reg_k0_n279), .ZN(reg_k0_n143)
         );
  NAND2_X1 reg_k0_U120 ( .A1(k[11]), .A2(reg_k0_n312), .ZN(reg_k0_n279) );
  NAND2_X1 reg_k0_U119 ( .A1(kext[139]), .A2(reg_k0_n311), .ZN(reg_k0_n280) );
  NAND2_X1 reg_k0_U118 ( .A1(reg_k0_n278), .A2(reg_k0_n277), .ZN(reg_k0_n142)
         );
  NAND2_X1 reg_k0_U117 ( .A1(k[10]), .A2(reg_k0_n338), .ZN(reg_k0_n277) );
  NAND2_X1 reg_k0_U116 ( .A1(kext[138]), .A2(reg_k0_n337), .ZN(reg_k0_n278) );
  NAND2_X1 reg_k0_U115 ( .A1(reg_k0_n276), .A2(reg_k0_n275), .ZN(reg_k0_n141)
         );
  NAND2_X1 reg_k0_U114 ( .A1(k[9]), .A2(reg_k0_n312), .ZN(reg_k0_n275) );
  NAND2_X1 reg_k0_U113 ( .A1(kext[137]), .A2(reg_k0_n311), .ZN(reg_k0_n276) );
  NAND2_X1 reg_k0_U112 ( .A1(reg_k0_n274), .A2(reg_k0_n273), .ZN(reg_k0_n140)
         );
  NAND2_X1 reg_k0_U111 ( .A1(k[8]), .A2(reg_k0_n338), .ZN(reg_k0_n273) );
  NAND2_X1 reg_k0_U110 ( .A1(kext[136]), .A2(reg_k0_n337), .ZN(reg_k0_n274) );
  NAND2_X1 reg_k0_U109 ( .A1(reg_k0_n272), .A2(reg_k0_n271), .ZN(reg_k0_n139)
         );
  NAND2_X1 reg_k0_U108 ( .A1(k[7]), .A2(reg_k0_n312), .ZN(reg_k0_n271) );
  NAND2_X1 reg_k0_U107 ( .A1(kext[135]), .A2(reg_k0_n311), .ZN(reg_k0_n272) );
  NAND2_X1 reg_k0_U106 ( .A1(reg_k0_n270), .A2(reg_k0_n269), .ZN(reg_k0_n138)
         );
  NAND2_X1 reg_k0_U105 ( .A1(k[6]), .A2(reg_k0_n338), .ZN(reg_k0_n269) );
  NAND2_X1 reg_k0_U104 ( .A1(kext[134]), .A2(reg_k0_n337), .ZN(reg_k0_n270) );
  NAND2_X1 reg_k0_U103 ( .A1(reg_k0_n268), .A2(reg_k0_n267), .ZN(reg_k0_n137)
         );
  NAND2_X1 reg_k0_U102 ( .A1(k[5]), .A2(reg_k0_n312), .ZN(reg_k0_n267) );
  INV_X1 reg_k0_U101 ( .A(reg_k0_n266), .ZN(reg_k0_n312) );
  NAND2_X1 reg_k0_U100 ( .A1(kext[133]), .A2(reg_k0_n311), .ZN(reg_k0_n268) );
  INV_X1 reg_k0_U99 ( .A(reg_k0_n265), .ZN(reg_k0_n311) );
  NAND2_X1 reg_k0_U98 ( .A1(reg_k0_n264), .A2(reg_k0_n263), .ZN(reg_k0_n136)
         );
  NAND2_X1 reg_k0_U97 ( .A1(k[4]), .A2(reg_k0_n338), .ZN(reg_k0_n263) );
  INV_X1 reg_k0_U96 ( .A(reg_k0_n266), .ZN(reg_k0_n338) );
  NAND2_X1 reg_k0_U95 ( .A1(kext[132]), .A2(reg_k0_n337), .ZN(reg_k0_n264) );
  INV_X1 reg_k0_U94 ( .A(reg_k0_n265), .ZN(reg_k0_n337) );
  NAND2_X1 reg_k0_U93 ( .A1(reg_k0_n262), .A2(reg_k0_n261), .ZN(reg_k0_n135)
         );
  NAND2_X1 reg_k0_U92 ( .A1(k[3]), .A2(reg_k0_n260), .ZN(reg_k0_n261) );
  NAND2_X1 reg_k0_U91 ( .A1(kext[131]), .A2(reg_k0_n259), .ZN(reg_k0_n262) );
  NAND2_X1 reg_k0_U90 ( .A1(reg_k0_n258), .A2(reg_k0_n257), .ZN(reg_k0_n134)
         );
  NAND2_X1 reg_k0_U89 ( .A1(k[2]), .A2(reg_k0_n260), .ZN(reg_k0_n257) );
  NAND2_X1 reg_k0_U88 ( .A1(kext[130]), .A2(reg_k0_n259), .ZN(reg_k0_n258) );
  NAND2_X1 reg_k0_U87 ( .A1(reg_k0_n256), .A2(reg_k0_n255), .ZN(reg_k0_n133)
         );
  NAND2_X1 reg_k0_U86 ( .A1(k[1]), .A2(reg_k0_n260), .ZN(reg_k0_n255) );
  NAND2_X1 reg_k0_U85 ( .A1(kext[129]), .A2(reg_k0_n259), .ZN(reg_k0_n256) );
  NAND2_X1 reg_k0_U84 ( .A1(reg_k0_n254), .A2(reg_k0_n253), .ZN(reg_k0_n132)
         );
  NAND2_X1 reg_k0_U83 ( .A1(k[0]), .A2(reg_k0_n260), .ZN(reg_k0_n253) );
  NAND2_X1 reg_k0_U82 ( .A1(kext[128]), .A2(reg_k0_n259), .ZN(reg_k0_n254) );
  NAND2_X1 reg_k0_U81 ( .A1(reg_k0_n252), .A2(reg_k0_n251), .ZN(reg_k0_n191)
         );
  NAND2_X1 reg_k0_U80 ( .A1(k[59]), .A2(reg_k0_n260), .ZN(reg_k0_n251) );
  NAND2_X1 reg_k0_U79 ( .A1(kext[187]), .A2(reg_k0_n259), .ZN(reg_k0_n252) );
  NAND2_X1 reg_k0_U78 ( .A1(reg_k0_n250), .A2(reg_k0_n249), .ZN(reg_k0_n190)
         );
  NAND2_X1 reg_k0_U77 ( .A1(k[58]), .A2(reg_k0_n260), .ZN(reg_k0_n249) );
  NAND2_X1 reg_k0_U76 ( .A1(kext[186]), .A2(reg_k0_n259), .ZN(reg_k0_n250) );
  NAND2_X1 reg_k0_U75 ( .A1(reg_k0_n248), .A2(reg_k0_n247), .ZN(reg_k0_n189)
         );
  NAND2_X1 reg_k0_U74 ( .A1(k[57]), .A2(reg_k0_n260), .ZN(reg_k0_n247) );
  NAND2_X1 reg_k0_U73 ( .A1(kext[185]), .A2(reg_k0_n259), .ZN(reg_k0_n248) );
  NAND2_X1 reg_k0_U72 ( .A1(reg_k0_n246), .A2(reg_k0_n245), .ZN(reg_k0_n188)
         );
  NAND2_X1 reg_k0_U71 ( .A1(k[56]), .A2(reg_k0_n260), .ZN(reg_k0_n245) );
  NAND2_X1 reg_k0_U70 ( .A1(kext[184]), .A2(reg_k0_n259), .ZN(reg_k0_n246) );
  NAND2_X1 reg_k0_U69 ( .A1(reg_k0_n244), .A2(reg_k0_n243), .ZN(reg_k0_n187)
         );
  NAND2_X1 reg_k0_U68 ( .A1(k[55]), .A2(reg_k0_n260), .ZN(reg_k0_n243) );
  NAND2_X1 reg_k0_U67 ( .A1(kext[183]), .A2(reg_k0_n259), .ZN(reg_k0_n244) );
  NAND2_X1 reg_k0_U66 ( .A1(reg_k0_n242), .A2(reg_k0_n241), .ZN(reg_k0_n186)
         );
  NAND2_X1 reg_k0_U65 ( .A1(k[54]), .A2(reg_k0_n240), .ZN(reg_k0_n241) );
  NAND2_X1 reg_k0_U64 ( .A1(kext[182]), .A2(reg_k0_n259), .ZN(reg_k0_n242) );
  NAND2_X1 reg_k0_U63 ( .A1(reg_k0_n239), .A2(reg_k0_n238), .ZN(reg_k0_n185)
         );
  NAND2_X1 reg_k0_U62 ( .A1(k[53]), .A2(reg_k0_n240), .ZN(reg_k0_n238) );
  NAND2_X1 reg_k0_U61 ( .A1(kext[181]), .A2(reg_k0_n259), .ZN(reg_k0_n239) );
  NAND2_X1 reg_k0_U60 ( .A1(reg_k0_n237), .A2(reg_k0_n236), .ZN(reg_k0_n184)
         );
  NAND2_X1 reg_k0_U59 ( .A1(k[52]), .A2(reg_k0_n240), .ZN(reg_k0_n236) );
  NAND2_X1 reg_k0_U58 ( .A1(kext[180]), .A2(reg_k0_n259), .ZN(reg_k0_n237) );
  NAND2_X1 reg_k0_U57 ( .A1(reg_k0_n235), .A2(reg_k0_n234), .ZN(reg_k0_n183)
         );
  NAND2_X1 reg_k0_U56 ( .A1(k[51]), .A2(reg_k0_n240), .ZN(reg_k0_n234) );
  NAND2_X1 reg_k0_U55 ( .A1(kext[179]), .A2(reg_k0_n259), .ZN(reg_k0_n235) );
  NAND2_X1 reg_k0_U54 ( .A1(reg_k0_n233), .A2(reg_k0_n232), .ZN(reg_k0_n182)
         );
  NAND2_X1 reg_k0_U53 ( .A1(k[50]), .A2(reg_k0_n240), .ZN(reg_k0_n232) );
  NAND2_X1 reg_k0_U52 ( .A1(kext[178]), .A2(reg_k0_n259), .ZN(reg_k0_n233) );
  NAND2_X1 reg_k0_U51 ( .A1(reg_k0_n231), .A2(reg_k0_n230), .ZN(reg_k0_n181)
         );
  NAND2_X1 reg_k0_U50 ( .A1(k[49]), .A2(reg_k0_n240), .ZN(reg_k0_n230) );
  NAND2_X1 reg_k0_U49 ( .A1(kext[177]), .A2(reg_k0_n229), .ZN(reg_k0_n231) );
  NAND2_X1 reg_k0_U48 ( .A1(reg_k0_n228), .A2(reg_k0_n227), .ZN(reg_k0_n180)
         );
  NAND2_X1 reg_k0_U47 ( .A1(k[48]), .A2(reg_k0_n240), .ZN(reg_k0_n227) );
  NAND2_X1 reg_k0_U46 ( .A1(kext[176]), .A2(reg_k0_n229), .ZN(reg_k0_n228) );
  NAND2_X1 reg_k0_U45 ( .A1(reg_k0_n226), .A2(reg_k0_n225), .ZN(reg_k0_n179)
         );
  NAND2_X1 reg_k0_U44 ( .A1(k[47]), .A2(reg_k0_n240), .ZN(reg_k0_n225) );
  NAND2_X1 reg_k0_U43 ( .A1(kext[175]), .A2(reg_k0_n229), .ZN(reg_k0_n226) );
  NAND2_X1 reg_k0_U42 ( .A1(reg_k0_n224), .A2(reg_k0_n223), .ZN(reg_k0_n178)
         );
  NAND2_X1 reg_k0_U41 ( .A1(k[46]), .A2(reg_k0_n240), .ZN(reg_k0_n223) );
  NAND2_X1 reg_k0_U40 ( .A1(kext[174]), .A2(reg_k0_n229), .ZN(reg_k0_n224) );
  NAND2_X1 reg_k0_U39 ( .A1(reg_k0_n222), .A2(reg_k0_n221), .ZN(reg_k0_n177)
         );
  NAND2_X1 reg_k0_U38 ( .A1(k[45]), .A2(reg_k0_n240), .ZN(reg_k0_n221) );
  NAND2_X1 reg_k0_U37 ( .A1(kext[173]), .A2(reg_k0_n229), .ZN(reg_k0_n222) );
  NAND2_X1 reg_k0_U36 ( .A1(reg_k0_n220), .A2(reg_k0_n219), .ZN(reg_k0_n176)
         );
  NAND2_X1 reg_k0_U35 ( .A1(k[44]), .A2(reg_k0_n240), .ZN(reg_k0_n219) );
  NAND2_X1 reg_k0_U34 ( .A1(kext[172]), .A2(reg_k0_n229), .ZN(reg_k0_n220) );
  NAND2_X1 reg_k0_U33 ( .A1(reg_k0_n218), .A2(reg_k0_n217), .ZN(reg_k0_n175)
         );
  NAND2_X1 reg_k0_U32 ( .A1(k[43]), .A2(reg_k0_n240), .ZN(reg_k0_n217) );
  NAND2_X1 reg_k0_U31 ( .A1(kext[171]), .A2(reg_k0_n229), .ZN(reg_k0_n218) );
  NAND2_X1 reg_k0_U30 ( .A1(reg_k0_n216), .A2(reg_k0_n215), .ZN(reg_k0_n174)
         );
  NAND2_X1 reg_k0_U29 ( .A1(k[42]), .A2(reg_k0_n240), .ZN(reg_k0_n215) );
  NAND2_X1 reg_k0_U28 ( .A1(kext[170]), .A2(reg_k0_n229), .ZN(reg_k0_n216) );
  NAND2_X1 reg_k0_U27 ( .A1(reg_k0_n214), .A2(reg_k0_n213), .ZN(reg_k0_n173)
         );
  NAND2_X1 reg_k0_U26 ( .A1(k[41]), .A2(reg_k0_n240), .ZN(reg_k0_n213) );
  NAND2_X1 reg_k0_U25 ( .A1(kext[169]), .A2(reg_k0_n229), .ZN(reg_k0_n214) );
  NAND2_X1 reg_k0_U24 ( .A1(reg_k0_n212), .A2(reg_k0_n211), .ZN(reg_k0_n172)
         );
  NAND2_X1 reg_k0_U23 ( .A1(k[40]), .A2(reg_k0_n240), .ZN(reg_k0_n211) );
  NAND2_X1 reg_k0_U22 ( .A1(kext[168]), .A2(reg_k0_n259), .ZN(reg_k0_n212) );
  NAND2_X1 reg_k0_U21 ( .A1(reg_k0_n210), .A2(reg_k0_n209), .ZN(reg_k0_n171)
         );
  NAND2_X1 reg_k0_U20 ( .A1(k[39]), .A2(reg_k0_n240), .ZN(reg_k0_n209) );
  NAND2_X1 reg_k0_U19 ( .A1(kext[167]), .A2(reg_k0_n259), .ZN(reg_k0_n210) );
  NAND2_X1 reg_k0_U18 ( .A1(reg_k0_n208), .A2(reg_k0_n207), .ZN(reg_k0_n170)
         );
  NAND2_X1 reg_k0_U17 ( .A1(k[38]), .A2(reg_k0_n240), .ZN(reg_k0_n207) );
  NAND2_X1 reg_k0_U16 ( .A1(kext[166]), .A2(reg_k0_n259), .ZN(reg_k0_n208) );
  NAND2_X1 reg_k0_U15 ( .A1(reg_k0_n206), .A2(reg_k0_n205), .ZN(reg_k0_n169)
         );
  NAND2_X1 reg_k0_U14 ( .A1(k[37]), .A2(reg_k0_n240), .ZN(reg_k0_n205) );
  NAND2_X1 reg_k0_U13 ( .A1(kext[165]), .A2(reg_k0_n259), .ZN(reg_k0_n206) );
  NAND2_X1 reg_k0_U12 ( .A1(reg_k0_n204), .A2(reg_k0_n203), .ZN(reg_k0_n168)
         );
  NAND2_X1 reg_k0_U11 ( .A1(reg_k0_n259), .A2(kext[164]), .ZN(reg_k0_n203) );
  INV_X1 reg_k0_U10 ( .A(reg_k0_n265), .ZN(reg_k0_n259) );
  INV_X1 reg_k0_U9 ( .A(reg_k0_n229), .ZN(reg_k0_n265) );
  NAND2_X1 reg_k0_U8 ( .A1(reg_k0_n240), .A2(k[36]), .ZN(reg_k0_n204) );
  INV_X1 reg_k0_U7 ( .A(reg_k0_n266), .ZN(reg_k0_n240) );
  INV_X1 reg_k0_U6 ( .A(reg_k0_n260), .ZN(reg_k0_n266) );
  INV_X1 reg_k0_U5 ( .A(en_sig), .ZN(reg_k0_n202) );
  NOR2_X1 reg_k0_U4 ( .A1(rst), .A2(reg_k0_n202), .ZN(reg_k0_n260) );
  NOR2_X1 reg_k0_U3 ( .A1(rst), .A2(en_sig), .ZN(reg_k0_n229) );
  DFF_X1 reg_k0_s_current_state_reg_0_ ( .D(reg_k0_n132), .CK(clk), .Q(
        kext[128]) );
  DFF_X1 reg_k0_s_current_state_reg_1_ ( .D(reg_k0_n133), .CK(clk), .Q(
        kext[129]) );
  DFF_X1 reg_k0_s_current_state_reg_2_ ( .D(reg_k0_n134), .CK(clk), .Q(
        kext[130]) );
  DFF_X1 reg_k0_s_current_state_reg_3_ ( .D(reg_k0_n135), .CK(clk), .Q(
        kext[131]) );
  DFF_X1 reg_k0_s_current_state_reg_4_ ( .D(reg_k0_n136), .CK(clk), .Q(
        kext[132]) );
  DFF_X1 reg_k0_s_current_state_reg_5_ ( .D(reg_k0_n137), .CK(clk), .Q(
        kext[133]) );
  DFF_X1 reg_k0_s_current_state_reg_6_ ( .D(reg_k0_n138), .CK(clk), .Q(
        kext[134]) );
  DFF_X1 reg_k0_s_current_state_reg_7_ ( .D(reg_k0_n139), .CK(clk), .Q(
        kext[135]) );
  DFF_X1 reg_k0_s_current_state_reg_8_ ( .D(reg_k0_n140), .CK(clk), .Q(
        kext[136]) );
  DFF_X1 reg_k0_s_current_state_reg_9_ ( .D(reg_k0_n141), .CK(clk), .Q(
        kext[137]) );
  DFF_X1 reg_k0_s_current_state_reg_10_ ( .D(reg_k0_n142), .CK(clk), .Q(
        kext[138]) );
  DFF_X1 reg_k0_s_current_state_reg_11_ ( .D(reg_k0_n143), .CK(clk), .Q(
        kext[139]) );
  DFF_X1 reg_k0_s_current_state_reg_12_ ( .D(reg_k0_n144), .CK(clk), .Q(
        kext[140]) );
  DFF_X1 reg_k0_s_current_state_reg_13_ ( .D(reg_k0_n145), .CK(clk), .Q(
        kext[141]) );
  DFF_X1 reg_k0_s_current_state_reg_14_ ( .D(reg_k0_n146), .CK(clk), .Q(
        kext[142]) );
  DFF_X1 reg_k0_s_current_state_reg_15_ ( .D(reg_k0_n147), .CK(clk), .Q(
        prince_inst_rc2_inv[15]) );
  DFF_X1 reg_k0_s_current_state_reg_16_ ( .D(reg_k0_n148), .CK(clk), .Q(
        kext[144]) );
  DFF_X1 reg_k0_s_current_state_reg_17_ ( .D(reg_k0_n149), .CK(clk), .Q(
        kext[145]) );
  DFF_X1 reg_k0_s_current_state_reg_18_ ( .D(reg_k0_n150), .CK(clk), .Q(
        kext[146]) );
  DFF_X1 reg_k0_s_current_state_reg_19_ ( .D(reg_k0_n151), .CK(clk), .Q(
        kext[147]) );
  DFF_X1 reg_k0_s_current_state_reg_20_ ( .D(reg_k0_n152), .CK(clk), .Q(
        kext[148]) );
  DFF_X1 reg_k0_s_current_state_reg_21_ ( .D(reg_k0_n153), .CK(clk), .Q(
        kext[149]) );
  DFF_X1 reg_k0_s_current_state_reg_22_ ( .D(reg_k0_n154), .CK(clk), .Q(
        kext[150]) );
  DFF_X1 reg_k0_s_current_state_reg_23_ ( .D(reg_k0_n155), .CK(clk), .Q(
        kext[151]) );
  DFF_X1 reg_k0_s_current_state_reg_24_ ( .D(reg_k0_n156), .CK(clk), .Q(
        kext[152]) );
  DFF_X1 reg_k0_s_current_state_reg_25_ ( .D(reg_k0_n157), .CK(clk), .Q(
        kext[153]) );
  DFF_X1 reg_k0_s_current_state_reg_26_ ( .D(reg_k0_n158), .CK(clk), .Q(
        kext[154]) );
  DFF_X1 reg_k0_s_current_state_reg_27_ ( .D(reg_k0_n159), .CK(clk), .Q(
        kext[155]) );
  DFF_X1 reg_k0_s_current_state_reg_28_ ( .D(reg_k0_n160), .CK(clk), .Q(
        kext[156]) );
  DFF_X1 reg_k0_s_current_state_reg_29_ ( .D(reg_k0_n161), .CK(clk), .Q(
        kext[157]) );
  DFF_X1 reg_k0_s_current_state_reg_30_ ( .D(reg_k0_n162), .CK(clk), .Q(
        kext[158]) );
  DFF_X1 reg_k0_s_current_state_reg_31_ ( .D(reg_k0_n163), .CK(clk), .Q(
        kext[159]) );
  DFF_X1 reg_k0_s_current_state_reg_32_ ( .D(reg_k0_n164), .CK(clk), .Q(
        kext[160]) );
  DFF_X1 reg_k0_s_current_state_reg_33_ ( .D(reg_k0_n165), .CK(clk), .Q(
        kext[161]) );
  DFF_X1 reg_k0_s_current_state_reg_34_ ( .D(reg_k0_n166), .CK(clk), .Q(
        kext[162]) );
  DFF_X1 reg_k0_s_current_state_reg_35_ ( .D(reg_k0_n167), .CK(clk), .Q(
        kext[163]) );
  DFF_X1 reg_k0_s_current_state_reg_36_ ( .D(reg_k0_n168), .CK(clk), .Q(
        kext[164]) );
  DFF_X1 reg_k0_s_current_state_reg_37_ ( .D(reg_k0_n169), .CK(clk), .Q(
        kext[165]) );
  DFF_X1 reg_k0_s_current_state_reg_38_ ( .D(reg_k0_n170), .CK(clk), .Q(
        kext[166]) );
  DFF_X1 reg_k0_s_current_state_reg_39_ ( .D(reg_k0_n171), .CK(clk), .Q(
        kext[167]) );
  DFF_X1 reg_k0_s_current_state_reg_40_ ( .D(reg_k0_n172), .CK(clk), .Q(
        kext[168]) );
  DFF_X1 reg_k0_s_current_state_reg_41_ ( .D(reg_k0_n173), .CK(clk), .Q(
        kext[169]) );
  DFF_X1 reg_k0_s_current_state_reg_42_ ( .D(reg_k0_n174), .CK(clk), .Q(
        kext[170]) );
  DFF_X1 reg_k0_s_current_state_reg_43_ ( .D(reg_k0_n175), .CK(clk), .Q(
        kext[171]) );
  DFF_X1 reg_k0_s_current_state_reg_44_ ( .D(reg_k0_n176), .CK(clk), .Q(
        kext[172]) );
  DFF_X1 reg_k0_s_current_state_reg_45_ ( .D(reg_k0_n177), .CK(clk), .Q(
        kext[173]) );
  DFF_X1 reg_k0_s_current_state_reg_46_ ( .D(reg_k0_n178), .CK(clk), .Q(
        kext[174]) );
  DFF_X1 reg_k0_s_current_state_reg_47_ ( .D(reg_k0_n179), .CK(clk), .Q(
        kext[175]) );
  DFF_X1 reg_k0_s_current_state_reg_48_ ( .D(reg_k0_n180), .CK(clk), .Q(
        kext[176]) );
  DFF_X1 reg_k0_s_current_state_reg_49_ ( .D(reg_k0_n181), .CK(clk), .Q(
        kext[177]) );
  DFF_X1 reg_k0_s_current_state_reg_50_ ( .D(reg_k0_n182), .CK(clk), .Q(
        kext[178]) );
  DFF_X1 reg_k0_s_current_state_reg_51_ ( .D(reg_k0_n183), .CK(clk), .Q(
        kext[179]) );
  DFF_X1 reg_k0_s_current_state_reg_52_ ( .D(reg_k0_n184), .CK(clk), .Q(
        kext[180]) );
  DFF_X1 reg_k0_s_current_state_reg_53_ ( .D(reg_k0_n185), .CK(clk), .Q(
        kext[181]) );
  DFF_X1 reg_k0_s_current_state_reg_54_ ( .D(reg_k0_n186), .CK(clk), .Q(
        kext[182]) );
  DFF_X1 reg_k0_s_current_state_reg_55_ ( .D(reg_k0_n187), .CK(clk), .Q(
        kext[183]) );
  DFF_X1 reg_k0_s_current_state_reg_56_ ( .D(reg_k0_n188), .CK(clk), .Q(
        kext[184]) );
  DFF_X1 reg_k0_s_current_state_reg_57_ ( .D(reg_k0_n189), .CK(clk), .Q(
        kext[185]) );
  DFF_X1 reg_k0_s_current_state_reg_58_ ( .D(reg_k0_n190), .CK(clk), .Q(
        kext[186]) );
  DFF_X1 reg_k0_s_current_state_reg_59_ ( .D(reg_k0_n191), .CK(clk), .Q(
        kext[187]) );
  DFF_X1 reg_k0_s_current_state_reg_60_ ( .D(reg_k0_n192), .CK(clk), .Q(
        kext[188]) );
  DFF_X1 reg_k0_s_current_state_reg_61_ ( .D(reg_k0_n193), .CK(clk), .Q(
        kext[189]) );
  DFF_X1 reg_k0_s_current_state_reg_62_ ( .D(reg_k0_n194), .CK(clk), .Q(
        kext[190]) );
  DFF_X1 reg_k0_s_current_state_reg_63_ ( .D(reg_k0_n195), .CK(clk), .Q(
        kext[191]) );
  NAND2_X1 reg_k1_U205 ( .A1(reg_k1_n532), .A2(reg_k1_n531), .ZN(reg_k1_n203)
         );
  NAND2_X1 reg_k1_U204 ( .A1(k[126]), .A2(reg_k1_n530), .ZN(reg_k1_n531) );
  NAND2_X1 reg_k1_U203 ( .A1(kext[125]), .A2(reg_k1_n529), .ZN(reg_k1_n532) );
  NAND2_X1 reg_k1_U202 ( .A1(reg_k1_n528), .A2(reg_k1_n527), .ZN(reg_k1_n204)
         );
  NAND2_X1 reg_k1_U201 ( .A1(k[125]), .A2(reg_k1_n530), .ZN(reg_k1_n527) );
  NAND2_X1 reg_k1_U200 ( .A1(kext[124]), .A2(reg_k1_n529), .ZN(reg_k1_n528) );
  NAND2_X1 reg_k1_U199 ( .A1(reg_k1_n526), .A2(reg_k1_n525), .ZN(reg_k1_n205)
         );
  NAND2_X1 reg_k1_U198 ( .A1(k[124]), .A2(reg_k1_n530), .ZN(reg_k1_n525) );
  NAND2_X1 reg_k1_U197 ( .A1(kext[123]), .A2(reg_k1_n529), .ZN(reg_k1_n526) );
  NAND2_X1 reg_k1_U196 ( .A1(reg_k1_n524), .A2(reg_k1_n523), .ZN(reg_k1_n230)
         );
  NAND2_X1 reg_k1_U195 ( .A1(k[99]), .A2(reg_k1_n530), .ZN(reg_k1_n523) );
  NAND2_X1 reg_k1_U194 ( .A1(kext[98]), .A2(reg_k1_n529), .ZN(reg_k1_n524) );
  NAND2_X1 reg_k1_U193 ( .A1(reg_k1_n522), .A2(reg_k1_n521), .ZN(reg_k1_n231)
         );
  NAND2_X1 reg_k1_U192 ( .A1(k[98]), .A2(reg_k1_n530), .ZN(reg_k1_n521) );
  NAND2_X1 reg_k1_U191 ( .A1(kext[97]), .A2(reg_k1_n529), .ZN(reg_k1_n522) );
  NAND2_X1 reg_k1_U190 ( .A1(reg_k1_n520), .A2(reg_k1_n519), .ZN(reg_k1_n232)
         );
  NAND2_X1 reg_k1_U189 ( .A1(k[97]), .A2(reg_k1_n530), .ZN(reg_k1_n519) );
  NAND2_X1 reg_k1_U188 ( .A1(kext[96]), .A2(reg_k1_n529), .ZN(reg_k1_n520) );
  NAND2_X1 reg_k1_U187 ( .A1(reg_k1_n518), .A2(reg_k1_n517), .ZN(reg_k1_n233)
         );
  NAND2_X1 reg_k1_U186 ( .A1(k[96]), .A2(reg_k1_n530), .ZN(reg_k1_n517) );
  NAND2_X1 reg_k1_U185 ( .A1(kext[95]), .A2(reg_k1_n529), .ZN(reg_k1_n518) );
  NAND2_X1 reg_k1_U184 ( .A1(reg_k1_n516), .A2(reg_k1_n515), .ZN(reg_k1_n234)
         );
  NAND2_X1 reg_k1_U183 ( .A1(k[95]), .A2(reg_k1_n530), .ZN(reg_k1_n515) );
  NAND2_X1 reg_k1_U182 ( .A1(kext[94]), .A2(reg_k1_n529), .ZN(reg_k1_n516) );
  NAND2_X1 reg_k1_U181 ( .A1(reg_k1_n514), .A2(reg_k1_n513), .ZN(reg_k1_n235)
         );
  NAND2_X1 reg_k1_U180 ( .A1(k[94]), .A2(reg_k1_n530), .ZN(reg_k1_n513) );
  NAND2_X1 reg_k1_U179 ( .A1(kext[93]), .A2(reg_k1_n529), .ZN(reg_k1_n514) );
  NAND2_X1 reg_k1_U178 ( .A1(reg_k1_n512), .A2(reg_k1_n511), .ZN(reg_k1_n236)
         );
  NAND2_X1 reg_k1_U177 ( .A1(k[93]), .A2(reg_k1_n530), .ZN(reg_k1_n511) );
  NAND2_X1 reg_k1_U176 ( .A1(kext[92]), .A2(reg_k1_n529), .ZN(reg_k1_n512) );
  NAND2_X1 reg_k1_U175 ( .A1(reg_k1_n510), .A2(reg_k1_n509), .ZN(reg_k1_n237)
         );
  NAND2_X1 reg_k1_U174 ( .A1(k[92]), .A2(reg_k1_n530), .ZN(reg_k1_n509) );
  NAND2_X1 reg_k1_U173 ( .A1(kext[91]), .A2(reg_k1_n529), .ZN(reg_k1_n510) );
  NAND2_X1 reg_k1_U172 ( .A1(reg_k1_n508), .A2(reg_k1_n507), .ZN(reg_k1_n238)
         );
  NAND2_X1 reg_k1_U171 ( .A1(k[91]), .A2(reg_k1_n530), .ZN(reg_k1_n507) );
  NAND2_X1 reg_k1_U170 ( .A1(kext[90]), .A2(reg_k1_n529), .ZN(reg_k1_n508) );
  NAND2_X1 reg_k1_U169 ( .A1(reg_k1_n506), .A2(reg_k1_n505), .ZN(reg_k1_n239)
         );
  NAND2_X1 reg_k1_U168 ( .A1(k[90]), .A2(reg_k1_n504), .ZN(reg_k1_n505) );
  NAND2_X1 reg_k1_U167 ( .A1(kext[89]), .A2(reg_k1_n503), .ZN(reg_k1_n506) );
  NAND2_X1 reg_k1_U166 ( .A1(reg_k1_n502), .A2(reg_k1_n501), .ZN(reg_k1_n240)
         );
  NAND2_X1 reg_k1_U165 ( .A1(k[89]), .A2(reg_k1_n504), .ZN(reg_k1_n501) );
  NAND2_X1 reg_k1_U164 ( .A1(kext[88]), .A2(reg_k1_n503), .ZN(reg_k1_n502) );
  NAND2_X1 reg_k1_U163 ( .A1(reg_k1_n500), .A2(reg_k1_n499), .ZN(reg_k1_n241)
         );
  NAND2_X1 reg_k1_U162 ( .A1(k[88]), .A2(reg_k1_n504), .ZN(reg_k1_n499) );
  NAND2_X1 reg_k1_U161 ( .A1(kext[87]), .A2(reg_k1_n503), .ZN(reg_k1_n500) );
  NAND2_X1 reg_k1_U160 ( .A1(reg_k1_n498), .A2(reg_k1_n497), .ZN(reg_k1_n242)
         );
  NAND2_X1 reg_k1_U159 ( .A1(k[87]), .A2(reg_k1_n504), .ZN(reg_k1_n497) );
  NAND2_X1 reg_k1_U158 ( .A1(kext[86]), .A2(reg_k1_n503), .ZN(reg_k1_n498) );
  NAND2_X1 reg_k1_U157 ( .A1(reg_k1_n496), .A2(reg_k1_n495), .ZN(reg_k1_n243)
         );
  NAND2_X1 reg_k1_U156 ( .A1(k[86]), .A2(reg_k1_n504), .ZN(reg_k1_n495) );
  NAND2_X1 reg_k1_U155 ( .A1(kext[85]), .A2(reg_k1_n503), .ZN(reg_k1_n496) );
  NAND2_X1 reg_k1_U154 ( .A1(reg_k1_n494), .A2(reg_k1_n493), .ZN(reg_k1_n244)
         );
  NAND2_X1 reg_k1_U153 ( .A1(k[85]), .A2(reg_k1_n504), .ZN(reg_k1_n493) );
  NAND2_X1 reg_k1_U152 ( .A1(kext[84]), .A2(reg_k1_n503), .ZN(reg_k1_n494) );
  NAND2_X1 reg_k1_U151 ( .A1(reg_k1_n492), .A2(reg_k1_n491), .ZN(reg_k1_n245)
         );
  NAND2_X1 reg_k1_U150 ( .A1(k[84]), .A2(reg_k1_n504), .ZN(reg_k1_n491) );
  NAND2_X1 reg_k1_U149 ( .A1(kext[83]), .A2(reg_k1_n503), .ZN(reg_k1_n492) );
  NAND2_X1 reg_k1_U148 ( .A1(reg_k1_n490), .A2(reg_k1_n489), .ZN(reg_k1_n246)
         );
  NAND2_X1 reg_k1_U147 ( .A1(k[83]), .A2(reg_k1_n504), .ZN(reg_k1_n489) );
  NAND2_X1 reg_k1_U146 ( .A1(kext[82]), .A2(reg_k1_n503), .ZN(reg_k1_n490) );
  NAND2_X1 reg_k1_U145 ( .A1(reg_k1_n488), .A2(reg_k1_n487), .ZN(reg_k1_n247)
         );
  NAND2_X1 reg_k1_U144 ( .A1(k[82]), .A2(reg_k1_n504), .ZN(reg_k1_n487) );
  NAND2_X1 reg_k1_U143 ( .A1(kext[81]), .A2(reg_k1_n503), .ZN(reg_k1_n488) );
  NAND2_X1 reg_k1_U142 ( .A1(reg_k1_n486), .A2(reg_k1_n485), .ZN(reg_k1_n248)
         );
  NAND2_X1 reg_k1_U141 ( .A1(k[81]), .A2(reg_k1_n504), .ZN(reg_k1_n485) );
  NAND2_X1 reg_k1_U140 ( .A1(kext[80]), .A2(reg_k1_n503), .ZN(reg_k1_n486) );
  NAND2_X1 reg_k1_U139 ( .A1(reg_k1_n484), .A2(reg_k1_n483), .ZN(reg_k1_n249)
         );
  NAND2_X1 reg_k1_U138 ( .A1(k[80]), .A2(reg_k1_n504), .ZN(reg_k1_n483) );
  NAND2_X1 reg_k1_U137 ( .A1(kext[79]), .A2(reg_k1_n503), .ZN(reg_k1_n484) );
  NAND2_X1 reg_k1_U136 ( .A1(reg_k1_n482), .A2(reg_k1_n481), .ZN(reg_k1_n250)
         );
  NAND2_X1 reg_k1_U135 ( .A1(k[79]), .A2(reg_k1_n504), .ZN(reg_k1_n481) );
  NAND2_X1 reg_k1_U134 ( .A1(kext[78]), .A2(reg_k1_n503), .ZN(reg_k1_n482) );
  NAND2_X1 reg_k1_U133 ( .A1(reg_k1_n480), .A2(reg_k1_n479), .ZN(reg_k1_n251)
         );
  NAND2_X1 reg_k1_U132 ( .A1(k[78]), .A2(reg_k1_n504), .ZN(reg_k1_n479) );
  NAND2_X1 reg_k1_U131 ( .A1(kext[77]), .A2(reg_k1_n503), .ZN(reg_k1_n480) );
  NAND2_X1 reg_k1_U130 ( .A1(reg_k1_n478), .A2(reg_k1_n477), .ZN(reg_k1_n252)
         );
  NAND2_X1 reg_k1_U129 ( .A1(k[77]), .A2(reg_k1_n530), .ZN(reg_k1_n477) );
  NAND2_X1 reg_k1_U128 ( .A1(kext[76]), .A2(reg_k1_n529), .ZN(reg_k1_n478) );
  NAND2_X1 reg_k1_U127 ( .A1(reg_k1_n476), .A2(reg_k1_n475), .ZN(reg_k1_n253)
         );
  NAND2_X1 reg_k1_U126 ( .A1(k[76]), .A2(reg_k1_n504), .ZN(reg_k1_n475) );
  NAND2_X1 reg_k1_U125 ( .A1(kext[75]), .A2(reg_k1_n503), .ZN(reg_k1_n476) );
  NAND2_X1 reg_k1_U124 ( .A1(reg_k1_n474), .A2(reg_k1_n473), .ZN(reg_k1_n254)
         );
  NAND2_X1 reg_k1_U123 ( .A1(k[75]), .A2(reg_k1_n530), .ZN(reg_k1_n473) );
  NAND2_X1 reg_k1_U122 ( .A1(kext[74]), .A2(reg_k1_n529), .ZN(reg_k1_n474) );
  NAND2_X1 reg_k1_U121 ( .A1(reg_k1_n472), .A2(reg_k1_n471), .ZN(reg_k1_n255)
         );
  NAND2_X1 reg_k1_U120 ( .A1(k[74]), .A2(reg_k1_n504), .ZN(reg_k1_n471) );
  NAND2_X1 reg_k1_U119 ( .A1(kext[73]), .A2(reg_k1_n503), .ZN(reg_k1_n472) );
  NAND2_X1 reg_k1_U118 ( .A1(reg_k1_n470), .A2(reg_k1_n469), .ZN(reg_k1_n256)
         );
  NAND2_X1 reg_k1_U117 ( .A1(k[73]), .A2(reg_k1_n530), .ZN(reg_k1_n469) );
  NAND2_X1 reg_k1_U116 ( .A1(kext[72]), .A2(reg_k1_n529), .ZN(reg_k1_n470) );
  NAND2_X1 reg_k1_U115 ( .A1(reg_k1_n468), .A2(reg_k1_n467), .ZN(reg_k1_n257)
         );
  NAND2_X1 reg_k1_U114 ( .A1(k[72]), .A2(reg_k1_n504), .ZN(reg_k1_n467) );
  NAND2_X1 reg_k1_U113 ( .A1(kext[71]), .A2(reg_k1_n503), .ZN(reg_k1_n468) );
  NAND2_X1 reg_k1_U112 ( .A1(reg_k1_n466), .A2(reg_k1_n465), .ZN(reg_k1_n258)
         );
  NAND2_X1 reg_k1_U111 ( .A1(k[71]), .A2(reg_k1_n530), .ZN(reg_k1_n465) );
  NAND2_X1 reg_k1_U110 ( .A1(kext[70]), .A2(reg_k1_n529), .ZN(reg_k1_n466) );
  NAND2_X1 reg_k1_U109 ( .A1(reg_k1_n464), .A2(reg_k1_n463), .ZN(reg_k1_n259)
         );
  NAND2_X1 reg_k1_U108 ( .A1(k[70]), .A2(reg_k1_n504), .ZN(reg_k1_n463) );
  NAND2_X1 reg_k1_U107 ( .A1(kext[69]), .A2(reg_k1_n503), .ZN(reg_k1_n464) );
  NAND2_X1 reg_k1_U106 ( .A1(reg_k1_n462), .A2(reg_k1_n461), .ZN(reg_k1_n260)
         );
  NAND2_X1 reg_k1_U105 ( .A1(k[69]), .A2(reg_k1_n530), .ZN(reg_k1_n461) );
  NAND2_X1 reg_k1_U104 ( .A1(kext[68]), .A2(reg_k1_n529), .ZN(reg_k1_n462) );
  NAND2_X1 reg_k1_U103 ( .A1(reg_k1_n460), .A2(reg_k1_n459), .ZN(reg_k1_n261)
         );
  NAND2_X1 reg_k1_U102 ( .A1(k[68]), .A2(reg_k1_n504), .ZN(reg_k1_n459) );
  INV_X1 reg_k1_U101 ( .A(reg_k1_n458), .ZN(reg_k1_n504) );
  NAND2_X1 reg_k1_U100 ( .A1(kext[67]), .A2(reg_k1_n503), .ZN(reg_k1_n460) );
  INV_X1 reg_k1_U99 ( .A(reg_k1_n457), .ZN(reg_k1_n503) );
  NAND2_X1 reg_k1_U98 ( .A1(reg_k1_n456), .A2(reg_k1_n455), .ZN(reg_k1_n262)
         );
  NAND2_X1 reg_k1_U97 ( .A1(k[67]), .A2(reg_k1_n530), .ZN(reg_k1_n455) );
  INV_X1 reg_k1_U96 ( .A(reg_k1_n458), .ZN(reg_k1_n530) );
  NAND2_X1 reg_k1_U95 ( .A1(kext[66]), .A2(reg_k1_n529), .ZN(reg_k1_n456) );
  INV_X1 reg_k1_U94 ( .A(reg_k1_n457), .ZN(reg_k1_n529) );
  NAND2_X1 reg_k1_U93 ( .A1(reg_k1_n454), .A2(reg_k1_n453), .ZN(reg_k1_n263)
         );
  NAND2_X1 reg_k1_U92 ( .A1(k[66]), .A2(reg_k1_n452), .ZN(reg_k1_n453) );
  NAND2_X1 reg_k1_U91 ( .A1(kext[65]), .A2(reg_k1_n451), .ZN(reg_k1_n454) );
  NAND2_X1 reg_k1_U90 ( .A1(reg_k1_n450), .A2(reg_k1_n449), .ZN(reg_k1_n264)
         );
  NAND2_X1 reg_k1_U89 ( .A1(k[65]), .A2(reg_k1_n452), .ZN(reg_k1_n449) );
  NAND2_X1 reg_k1_U88 ( .A1(kext[1]), .A2(reg_k1_n451), .ZN(reg_k1_n450) );
  NAND2_X1 reg_k1_U87 ( .A1(reg_k1_n448), .A2(reg_k1_n447), .ZN(reg_k1_n265)
         );
  NAND2_X1 reg_k1_U86 ( .A1(k[64]), .A2(reg_k1_n452), .ZN(reg_k1_n447) );
  NAND2_X1 reg_k1_U85 ( .A1(kext[127]), .A2(reg_k1_n451), .ZN(reg_k1_n448) );
  NAND2_X1 reg_k1_U84 ( .A1(reg_k1_n446), .A2(reg_k1_n445), .ZN(reg_k1_n206)
         );
  NAND2_X1 reg_k1_U83 ( .A1(k[123]), .A2(reg_k1_n452), .ZN(reg_k1_n445) );
  NAND2_X1 reg_k1_U82 ( .A1(kext[122]), .A2(reg_k1_n451), .ZN(reg_k1_n446) );
  NAND2_X1 reg_k1_U81 ( .A1(reg_k1_n444), .A2(reg_k1_n443), .ZN(reg_k1_n207)
         );
  NAND2_X1 reg_k1_U80 ( .A1(k[122]), .A2(reg_k1_n452), .ZN(reg_k1_n443) );
  NAND2_X1 reg_k1_U79 ( .A1(kext[121]), .A2(reg_k1_n451), .ZN(reg_k1_n444) );
  NAND2_X1 reg_k1_U78 ( .A1(reg_k1_n442), .A2(reg_k1_n441), .ZN(reg_k1_n208)
         );
  NAND2_X1 reg_k1_U77 ( .A1(k[121]), .A2(reg_k1_n452), .ZN(reg_k1_n441) );
  NAND2_X1 reg_k1_U76 ( .A1(kext[120]), .A2(reg_k1_n451), .ZN(reg_k1_n442) );
  NAND2_X1 reg_k1_U75 ( .A1(reg_k1_n440), .A2(reg_k1_n439), .ZN(reg_k1_n209)
         );
  NAND2_X1 reg_k1_U74 ( .A1(k[120]), .A2(reg_k1_n452), .ZN(reg_k1_n439) );
  NAND2_X1 reg_k1_U73 ( .A1(kext[119]), .A2(reg_k1_n451), .ZN(reg_k1_n440) );
  NAND2_X1 reg_k1_U72 ( .A1(reg_k1_n438), .A2(reg_k1_n437), .ZN(reg_k1_n210)
         );
  NAND2_X1 reg_k1_U71 ( .A1(k[119]), .A2(reg_k1_n452), .ZN(reg_k1_n437) );
  NAND2_X1 reg_k1_U70 ( .A1(kext[118]), .A2(reg_k1_n451), .ZN(reg_k1_n438) );
  NAND2_X1 reg_k1_U69 ( .A1(reg_k1_n436), .A2(reg_k1_n435), .ZN(reg_k1_n211)
         );
  NAND2_X1 reg_k1_U68 ( .A1(k[118]), .A2(reg_k1_n452), .ZN(reg_k1_n435) );
  NAND2_X1 reg_k1_U67 ( .A1(kext[117]), .A2(reg_k1_n451), .ZN(reg_k1_n436) );
  NAND2_X1 reg_k1_U66 ( .A1(reg_k1_n434), .A2(reg_k1_n433), .ZN(reg_k1_n212)
         );
  NAND2_X1 reg_k1_U65 ( .A1(k[117]), .A2(reg_k1_n432), .ZN(reg_k1_n433) );
  NAND2_X1 reg_k1_U64 ( .A1(kext[116]), .A2(reg_k1_n451), .ZN(reg_k1_n434) );
  NAND2_X1 reg_k1_U63 ( .A1(reg_k1_n431), .A2(reg_k1_n430), .ZN(reg_k1_n213)
         );
  NAND2_X1 reg_k1_U62 ( .A1(k[116]), .A2(reg_k1_n432), .ZN(reg_k1_n430) );
  NAND2_X1 reg_k1_U61 ( .A1(kext[115]), .A2(reg_k1_n451), .ZN(reg_k1_n431) );
  NAND2_X1 reg_k1_U60 ( .A1(reg_k1_n429), .A2(reg_k1_n428), .ZN(reg_k1_n214)
         );
  NAND2_X1 reg_k1_U59 ( .A1(k[115]), .A2(reg_k1_n432), .ZN(reg_k1_n428) );
  NAND2_X1 reg_k1_U58 ( .A1(kext[114]), .A2(reg_k1_n451), .ZN(reg_k1_n429) );
  NAND2_X1 reg_k1_U57 ( .A1(reg_k1_n427), .A2(reg_k1_n426), .ZN(reg_k1_n215)
         );
  NAND2_X1 reg_k1_U56 ( .A1(k[114]), .A2(reg_k1_n432), .ZN(reg_k1_n426) );
  NAND2_X1 reg_k1_U55 ( .A1(kext[113]), .A2(reg_k1_n451), .ZN(reg_k1_n427) );
  NAND2_X1 reg_k1_U54 ( .A1(reg_k1_n425), .A2(reg_k1_n424), .ZN(reg_k1_n216)
         );
  NAND2_X1 reg_k1_U53 ( .A1(k[113]), .A2(reg_k1_n432), .ZN(reg_k1_n424) );
  NAND2_X1 reg_k1_U52 ( .A1(kext[112]), .A2(reg_k1_n451), .ZN(reg_k1_n425) );
  NAND2_X1 reg_k1_U51 ( .A1(reg_k1_n423), .A2(reg_k1_n422), .ZN(reg_k1_n217)
         );
  NAND2_X1 reg_k1_U50 ( .A1(k[112]), .A2(reg_k1_n432), .ZN(reg_k1_n422) );
  NAND2_X1 reg_k1_U49 ( .A1(kext[111]), .A2(reg_k1_n421), .ZN(reg_k1_n423) );
  NAND2_X1 reg_k1_U48 ( .A1(reg_k1_n420), .A2(reg_k1_n419), .ZN(reg_k1_n218)
         );
  NAND2_X1 reg_k1_U47 ( .A1(k[111]), .A2(reg_k1_n432), .ZN(reg_k1_n419) );
  NAND2_X1 reg_k1_U46 ( .A1(kext[110]), .A2(reg_k1_n421), .ZN(reg_k1_n420) );
  NAND2_X1 reg_k1_U45 ( .A1(reg_k1_n418), .A2(reg_k1_n417), .ZN(reg_k1_n219)
         );
  NAND2_X1 reg_k1_U44 ( .A1(k[110]), .A2(reg_k1_n432), .ZN(reg_k1_n417) );
  NAND2_X1 reg_k1_U43 ( .A1(kext[109]), .A2(reg_k1_n421), .ZN(reg_k1_n418) );
  NAND2_X1 reg_k1_U42 ( .A1(reg_k1_n416), .A2(reg_k1_n415), .ZN(reg_k1_n220)
         );
  NAND2_X1 reg_k1_U41 ( .A1(k[109]), .A2(reg_k1_n432), .ZN(reg_k1_n415) );
  NAND2_X1 reg_k1_U40 ( .A1(kext[108]), .A2(reg_k1_n421), .ZN(reg_k1_n416) );
  NAND2_X1 reg_k1_U39 ( .A1(reg_k1_n414), .A2(reg_k1_n413), .ZN(reg_k1_n221)
         );
  NAND2_X1 reg_k1_U38 ( .A1(k[108]), .A2(reg_k1_n432), .ZN(reg_k1_n413) );
  NAND2_X1 reg_k1_U37 ( .A1(kext[107]), .A2(reg_k1_n421), .ZN(reg_k1_n414) );
  NAND2_X1 reg_k1_U36 ( .A1(reg_k1_n412), .A2(reg_k1_n411), .ZN(reg_k1_n222)
         );
  NAND2_X1 reg_k1_U35 ( .A1(k[107]), .A2(reg_k1_n432), .ZN(reg_k1_n411) );
  NAND2_X1 reg_k1_U34 ( .A1(kext[106]), .A2(reg_k1_n421), .ZN(reg_k1_n412) );
  NAND2_X1 reg_k1_U33 ( .A1(reg_k1_n410), .A2(reg_k1_n409), .ZN(reg_k1_n223)
         );
  NAND2_X1 reg_k1_U32 ( .A1(k[106]), .A2(reg_k1_n432), .ZN(reg_k1_n409) );
  NAND2_X1 reg_k1_U31 ( .A1(kext[105]), .A2(reg_k1_n421), .ZN(reg_k1_n410) );
  NAND2_X1 reg_k1_U30 ( .A1(reg_k1_n408), .A2(reg_k1_n407), .ZN(reg_k1_n224)
         );
  NAND2_X1 reg_k1_U29 ( .A1(k[105]), .A2(reg_k1_n432), .ZN(reg_k1_n407) );
  NAND2_X1 reg_k1_U28 ( .A1(kext[104]), .A2(reg_k1_n421), .ZN(reg_k1_n408) );
  NAND2_X1 reg_k1_U27 ( .A1(reg_k1_n406), .A2(reg_k1_n405), .ZN(reg_k1_n225)
         );
  NAND2_X1 reg_k1_U26 ( .A1(k[104]), .A2(reg_k1_n432), .ZN(reg_k1_n405) );
  NAND2_X1 reg_k1_U25 ( .A1(kext[103]), .A2(reg_k1_n421), .ZN(reg_k1_n406) );
  NAND2_X1 reg_k1_U24 ( .A1(reg_k1_n404), .A2(reg_k1_n403), .ZN(reg_k1_n226)
         );
  NAND2_X1 reg_k1_U23 ( .A1(k[103]), .A2(reg_k1_n432), .ZN(reg_k1_n403) );
  NAND2_X1 reg_k1_U22 ( .A1(kext[102]), .A2(reg_k1_n451), .ZN(reg_k1_n404) );
  NAND2_X1 reg_k1_U21 ( .A1(reg_k1_n402), .A2(reg_k1_n401), .ZN(reg_k1_n227)
         );
  NAND2_X1 reg_k1_U20 ( .A1(k[102]), .A2(reg_k1_n432), .ZN(reg_k1_n401) );
  NAND2_X1 reg_k1_U19 ( .A1(kext[101]), .A2(reg_k1_n451), .ZN(reg_k1_n402) );
  NAND2_X1 reg_k1_U18 ( .A1(reg_k1_n400), .A2(reg_k1_n399), .ZN(reg_k1_n228)
         );
  NAND2_X1 reg_k1_U17 ( .A1(k[101]), .A2(reg_k1_n432), .ZN(reg_k1_n399) );
  NAND2_X1 reg_k1_U16 ( .A1(kext[100]), .A2(reg_k1_n451), .ZN(reg_k1_n400) );
  NAND2_X1 reg_k1_U15 ( .A1(reg_k1_n398), .A2(reg_k1_n397), .ZN(reg_k1_n229)
         );
  NAND2_X1 reg_k1_U14 ( .A1(k[100]), .A2(reg_k1_n432), .ZN(reg_k1_n397) );
  NAND2_X1 reg_k1_U13 ( .A1(kext[99]), .A2(reg_k1_n451), .ZN(reg_k1_n398) );
  NAND2_X1 reg_k1_U12 ( .A1(reg_k1_n396), .A2(reg_k1_n395), .ZN(reg_k1_n202)
         );
  NAND2_X1 reg_k1_U11 ( .A1(reg_k1_n451), .A2(kext[126]), .ZN(reg_k1_n395) );
  INV_X1 reg_k1_U10 ( .A(reg_k1_n457), .ZN(reg_k1_n451) );
  INV_X1 reg_k1_U9 ( .A(reg_k1_n421), .ZN(reg_k1_n457) );
  NAND2_X1 reg_k1_U8 ( .A1(reg_k1_n432), .A2(k[127]), .ZN(reg_k1_n396) );
  INV_X1 reg_k1_U7 ( .A(reg_k1_n458), .ZN(reg_k1_n432) );
  INV_X1 reg_k1_U6 ( .A(reg_k1_n452), .ZN(reg_k1_n458) );
  INV_X1 reg_k1_U5 ( .A(en_sig), .ZN(reg_k1_n394) );
  NOR2_X1 reg_k1_U4 ( .A1(rst), .A2(reg_k1_n394), .ZN(reg_k1_n452) );
  NOR2_X1 reg_k1_U3 ( .A1(rst), .A2(en_sig), .ZN(reg_k1_n421) );
  DFF_X1 reg_k1_s_current_state_reg_0_ ( .D(reg_k1_n265), .CK(clk), .Q(
        kext[127]) );
  DFF_X1 reg_k1_s_current_state_reg_1_ ( .D(reg_k1_n264), .CK(clk), .Q(kext[1]) );
  DFF_X1 reg_k1_s_current_state_reg_2_ ( .D(reg_k1_n263), .CK(clk), .Q(
        kext[65]) );
  DFF_X1 reg_k1_s_current_state_reg_3_ ( .D(reg_k1_n262), .CK(clk), .Q(
        kext[66]) );
  DFF_X1 reg_k1_s_current_state_reg_4_ ( .D(reg_k1_n261), .CK(clk), .Q(
        kext[67]) );
  DFF_X1 reg_k1_s_current_state_reg_5_ ( .D(reg_k1_n260), .CK(clk), .Q(
        kext[68]) );
  DFF_X1 reg_k1_s_current_state_reg_6_ ( .D(reg_k1_n259), .CK(clk), .Q(
        kext[69]) );
  DFF_X1 reg_k1_s_current_state_reg_7_ ( .D(reg_k1_n258), .CK(clk), .Q(
        kext[70]) );
  DFF_X1 reg_k1_s_current_state_reg_8_ ( .D(reg_k1_n257), .CK(clk), .Q(
        kext[71]) );
  DFF_X1 reg_k1_s_current_state_reg_9_ ( .D(reg_k1_n256), .CK(clk), .Q(
        kext[72]) );
  DFF_X1 reg_k1_s_current_state_reg_10_ ( .D(reg_k1_n255), .CK(clk), .Q(
        kext[73]) );
  DFF_X1 reg_k1_s_current_state_reg_11_ ( .D(reg_k1_n254), .CK(clk), .Q(
        kext[74]) );
  DFF_X1 reg_k1_s_current_state_reg_12_ ( .D(reg_k1_n253), .CK(clk), .Q(
        kext[75]) );
  DFF_X1 reg_k1_s_current_state_reg_13_ ( .D(reg_k1_n252), .CK(clk), .Q(
        kext[76]) );
  DFF_X1 reg_k1_s_current_state_reg_14_ ( .D(reg_k1_n251), .CK(clk), .Q(
        kext[77]) );
  DFF_X1 reg_k1_s_current_state_reg_15_ ( .D(reg_k1_n250), .CK(clk), .Q(
        kext[78]) );
  DFF_X1 reg_k1_s_current_state_reg_16_ ( .D(reg_k1_n249), .CK(clk), .Q(
        kext[79]) );
  DFF_X1 reg_k1_s_current_state_reg_17_ ( .D(reg_k1_n248), .CK(clk), .Q(
        kext[80]) );
  DFF_X1 reg_k1_s_current_state_reg_18_ ( .D(reg_k1_n247), .CK(clk), .Q(
        kext[81]) );
  DFF_X1 reg_k1_s_current_state_reg_19_ ( .D(reg_k1_n246), .CK(clk), .Q(
        kext[82]) );
  DFF_X1 reg_k1_s_current_state_reg_20_ ( .D(reg_k1_n245), .CK(clk), .Q(
        kext[83]) );
  DFF_X1 reg_k1_s_current_state_reg_21_ ( .D(reg_k1_n244), .CK(clk), .Q(
        kext[84]) );
  DFF_X1 reg_k1_s_current_state_reg_22_ ( .D(reg_k1_n243), .CK(clk), .Q(
        kext[85]) );
  DFF_X1 reg_k1_s_current_state_reg_23_ ( .D(reg_k1_n242), .CK(clk), .Q(
        kext[86]) );
  DFF_X1 reg_k1_s_current_state_reg_24_ ( .D(reg_k1_n241), .CK(clk), .Q(
        kext[87]) );
  DFF_X1 reg_k1_s_current_state_reg_25_ ( .D(reg_k1_n240), .CK(clk), .Q(
        kext[88]) );
  DFF_X1 reg_k1_s_current_state_reg_26_ ( .D(reg_k1_n239), .CK(clk), .Q(
        kext[89]) );
  DFF_X1 reg_k1_s_current_state_reg_27_ ( .D(reg_k1_n238), .CK(clk), .Q(
        kext[90]) );
  DFF_X1 reg_k1_s_current_state_reg_28_ ( .D(reg_k1_n237), .CK(clk), .Q(
        kext[91]) );
  DFF_X1 reg_k1_s_current_state_reg_29_ ( .D(reg_k1_n236), .CK(clk), .Q(
        kext[92]) );
  DFF_X1 reg_k1_s_current_state_reg_30_ ( .D(reg_k1_n235), .CK(clk), .Q(
        kext[93]) );
  DFF_X1 reg_k1_s_current_state_reg_31_ ( .D(reg_k1_n234), .CK(clk), .Q(
        kext[94]) );
  DFF_X1 reg_k1_s_current_state_reg_32_ ( .D(reg_k1_n233), .CK(clk), .Q(
        kext[95]) );
  DFF_X1 reg_k1_s_current_state_reg_33_ ( .D(reg_k1_n232), .CK(clk), .Q(
        kext[96]) );
  DFF_X1 reg_k1_s_current_state_reg_34_ ( .D(reg_k1_n231), .CK(clk), .Q(
        kext[97]) );
  DFF_X1 reg_k1_s_current_state_reg_35_ ( .D(reg_k1_n230), .CK(clk), .Q(
        kext[98]) );
  DFF_X1 reg_k1_s_current_state_reg_36_ ( .D(reg_k1_n229), .CK(clk), .Q(
        kext[99]) );
  DFF_X1 reg_k1_s_current_state_reg_37_ ( .D(reg_k1_n228), .CK(clk), .Q(
        kext[100]) );
  DFF_X1 reg_k1_s_current_state_reg_38_ ( .D(reg_k1_n227), .CK(clk), .Q(
        kext[101]) );
  DFF_X1 reg_k1_s_current_state_reg_39_ ( .D(reg_k1_n226), .CK(clk), .Q(
        kext[102]) );
  DFF_X1 reg_k1_s_current_state_reg_40_ ( .D(reg_k1_n225), .CK(clk), .Q(
        kext[103]) );
  DFF_X1 reg_k1_s_current_state_reg_41_ ( .D(reg_k1_n224), .CK(clk), .Q(
        kext[104]) );
  DFF_X1 reg_k1_s_current_state_reg_42_ ( .D(reg_k1_n223), .CK(clk), .Q(
        kext[105]) );
  DFF_X1 reg_k1_s_current_state_reg_43_ ( .D(reg_k1_n222), .CK(clk), .Q(
        kext[106]) );
  DFF_X1 reg_k1_s_current_state_reg_44_ ( .D(reg_k1_n221), .CK(clk), .Q(
        kext[107]) );
  DFF_X1 reg_k1_s_current_state_reg_45_ ( .D(reg_k1_n220), .CK(clk), .Q(
        kext[108]) );
  DFF_X1 reg_k1_s_current_state_reg_46_ ( .D(reg_k1_n219), .CK(clk), .Q(
        kext[109]) );
  DFF_X1 reg_k1_s_current_state_reg_47_ ( .D(reg_k1_n218), .CK(clk), .Q(
        kext[110]) );
  DFF_X1 reg_k1_s_current_state_reg_48_ ( .D(reg_k1_n217), .CK(clk), .Q(
        kext[111]) );
  DFF_X1 reg_k1_s_current_state_reg_49_ ( .D(reg_k1_n216), .CK(clk), .Q(
        kext[112]) );
  DFF_X1 reg_k1_s_current_state_reg_50_ ( .D(reg_k1_n215), .CK(clk), .Q(
        kext[113]) );
  DFF_X1 reg_k1_s_current_state_reg_51_ ( .D(reg_k1_n214), .CK(clk), .Q(
        kext[114]) );
  DFF_X1 reg_k1_s_current_state_reg_52_ ( .D(reg_k1_n213), .CK(clk), .Q(
        kext[115]) );
  DFF_X1 reg_k1_s_current_state_reg_53_ ( .D(reg_k1_n212), .CK(clk), .Q(
        kext[116]) );
  DFF_X1 reg_k1_s_current_state_reg_54_ ( .D(reg_k1_n211), .CK(clk), .Q(
        kext[117]) );
  DFF_X1 reg_k1_s_current_state_reg_55_ ( .D(reg_k1_n210), .CK(clk), .Q(
        kext[118]) );
  DFF_X1 reg_k1_s_current_state_reg_56_ ( .D(reg_k1_n209), .CK(clk), .Q(
        kext[119]) );
  DFF_X1 reg_k1_s_current_state_reg_57_ ( .D(reg_k1_n208), .CK(clk), .Q(
        kext[120]) );
  DFF_X1 reg_k1_s_current_state_reg_58_ ( .D(reg_k1_n207), .CK(clk), .Q(
        kext[121]) );
  DFF_X1 reg_k1_s_current_state_reg_59_ ( .D(reg_k1_n206), .CK(clk), .Q(
        kext[122]) );
  DFF_X1 reg_k1_s_current_state_reg_60_ ( .D(reg_k1_n205), .CK(clk), .Q(
        kext[123]) );
  DFF_X1 reg_k1_s_current_state_reg_61_ ( .D(reg_k1_n204), .CK(clk), .Q(
        kext[124]) );
  DFF_X1 reg_k1_s_current_state_reg_62_ ( .D(reg_k1_n203), .CK(clk), .Q(
        kext[125]) );
  DFF_X1 reg_k1_s_current_state_reg_63_ ( .D(reg_k1_n202), .CK(clk), .Q(
        kext[126]) );
  NAND2_X1 reg_p0_U204 ( .A1(reg_p0_n531), .A2(reg_p0_n530), .ZN(reg_p0_n202)
         );
  NAND2_X1 reg_p0_U203 ( .A1(p0[63]), .A2(reg_p0_n529), .ZN(reg_p0_n530) );
  NAND2_X1 reg_p0_U202 ( .A1(p0_reg[63]), .A2(reg_p0_n528), .ZN(reg_p0_n531)
         );
  NAND2_X1 reg_p0_U201 ( .A1(reg_p0_n527), .A2(reg_p0_n526), .ZN(reg_p0_n203)
         );
  NAND2_X1 reg_p0_U200 ( .A1(p0[62]), .A2(reg_p0_n529), .ZN(reg_p0_n526) );
  NAND2_X1 reg_p0_U199 ( .A1(p0_reg[62]), .A2(reg_p0_n528), .ZN(reg_p0_n527)
         );
  NAND2_X1 reg_p0_U198 ( .A1(reg_p0_n525), .A2(reg_p0_n524), .ZN(reg_p0_n204)
         );
  NAND2_X1 reg_p0_U197 ( .A1(p0[61]), .A2(reg_p0_n529), .ZN(reg_p0_n524) );
  NAND2_X1 reg_p0_U196 ( .A1(p0_reg[61]), .A2(reg_p0_n528), .ZN(reg_p0_n525)
         );
  NAND2_X1 reg_p0_U195 ( .A1(reg_p0_n523), .A2(reg_p0_n522), .ZN(reg_p0_n205)
         );
  NAND2_X1 reg_p0_U194 ( .A1(p0[60]), .A2(reg_p0_n529), .ZN(reg_p0_n522) );
  NAND2_X1 reg_p0_U193 ( .A1(p0_reg[60]), .A2(reg_p0_n528), .ZN(reg_p0_n523)
         );
  NAND2_X1 reg_p0_U192 ( .A1(reg_p0_n521), .A2(reg_p0_n520), .ZN(reg_p0_n230)
         );
  NAND2_X1 reg_p0_U191 ( .A1(p0[35]), .A2(reg_p0_n529), .ZN(reg_p0_n520) );
  NAND2_X1 reg_p0_U190 ( .A1(p0_reg[35]), .A2(reg_p0_n528), .ZN(reg_p0_n521)
         );
  NAND2_X1 reg_p0_U189 ( .A1(reg_p0_n519), .A2(reg_p0_n518), .ZN(reg_p0_n231)
         );
  NAND2_X1 reg_p0_U188 ( .A1(p0[34]), .A2(reg_p0_n529), .ZN(reg_p0_n518) );
  NAND2_X1 reg_p0_U187 ( .A1(p0_reg[34]), .A2(reg_p0_n528), .ZN(reg_p0_n519)
         );
  NAND2_X1 reg_p0_U186 ( .A1(reg_p0_n517), .A2(reg_p0_n516), .ZN(reg_p0_n232)
         );
  NAND2_X1 reg_p0_U185 ( .A1(p0[33]), .A2(reg_p0_n529), .ZN(reg_p0_n516) );
  NAND2_X1 reg_p0_U184 ( .A1(p0_reg[33]), .A2(reg_p0_n528), .ZN(reg_p0_n517)
         );
  NAND2_X1 reg_p0_U183 ( .A1(reg_p0_n515), .A2(reg_p0_n514), .ZN(reg_p0_n233)
         );
  NAND2_X1 reg_p0_U182 ( .A1(p0[32]), .A2(reg_p0_n529), .ZN(reg_p0_n514) );
  NAND2_X1 reg_p0_U181 ( .A1(p0_reg[32]), .A2(reg_p0_n528), .ZN(reg_p0_n515)
         );
  NAND2_X1 reg_p0_U180 ( .A1(reg_p0_n513), .A2(reg_p0_n512), .ZN(reg_p0_n234)
         );
  NAND2_X1 reg_p0_U179 ( .A1(p0[31]), .A2(reg_p0_n529), .ZN(reg_p0_n512) );
  NAND2_X1 reg_p0_U178 ( .A1(p0_reg[31]), .A2(reg_p0_n528), .ZN(reg_p0_n513)
         );
  NAND2_X1 reg_p0_U177 ( .A1(reg_p0_n511), .A2(reg_p0_n510), .ZN(reg_p0_n235)
         );
  NAND2_X1 reg_p0_U176 ( .A1(p0[30]), .A2(reg_p0_n529), .ZN(reg_p0_n510) );
  NAND2_X1 reg_p0_U175 ( .A1(p0_reg[30]), .A2(reg_p0_n528), .ZN(reg_p0_n511)
         );
  NAND2_X1 reg_p0_U174 ( .A1(reg_p0_n509), .A2(reg_p0_n508), .ZN(reg_p0_n236)
         );
  NAND2_X1 reg_p0_U173 ( .A1(p0[29]), .A2(reg_p0_n529), .ZN(reg_p0_n508) );
  NAND2_X1 reg_p0_U172 ( .A1(p0_reg[29]), .A2(reg_p0_n528), .ZN(reg_p0_n509)
         );
  NAND2_X1 reg_p0_U171 ( .A1(reg_p0_n507), .A2(reg_p0_n506), .ZN(reg_p0_n237)
         );
  NAND2_X1 reg_p0_U170 ( .A1(p0[28]), .A2(reg_p0_n529), .ZN(reg_p0_n506) );
  NAND2_X1 reg_p0_U169 ( .A1(p0_reg[28]), .A2(reg_p0_n528), .ZN(reg_p0_n507)
         );
  NAND2_X1 reg_p0_U168 ( .A1(reg_p0_n505), .A2(reg_p0_n504), .ZN(reg_p0_n238)
         );
  NAND2_X1 reg_p0_U167 ( .A1(p0[27]), .A2(reg_p0_n452), .ZN(reg_p0_n504) );
  NAND2_X1 reg_p0_U166 ( .A1(p0_reg[27]), .A2(reg_p0_n503), .ZN(reg_p0_n505)
         );
  NAND2_X1 reg_p0_U165 ( .A1(reg_p0_n502), .A2(reg_p0_n501), .ZN(reg_p0_n239)
         );
  NAND2_X1 reg_p0_U164 ( .A1(p0[26]), .A2(reg_p0_n452), .ZN(reg_p0_n501) );
  NAND2_X1 reg_p0_U163 ( .A1(p0_reg[26]), .A2(reg_p0_n503), .ZN(reg_p0_n502)
         );
  NAND2_X1 reg_p0_U162 ( .A1(reg_p0_n500), .A2(reg_p0_n499), .ZN(reg_p0_n240)
         );
  NAND2_X1 reg_p0_U161 ( .A1(p0[25]), .A2(reg_p0_n452), .ZN(reg_p0_n499) );
  NAND2_X1 reg_p0_U160 ( .A1(p0_reg[25]), .A2(reg_p0_n503), .ZN(reg_p0_n500)
         );
  NAND2_X1 reg_p0_U159 ( .A1(reg_p0_n498), .A2(reg_p0_n497), .ZN(reg_p0_n241)
         );
  NAND2_X1 reg_p0_U158 ( .A1(p0[24]), .A2(reg_p0_n452), .ZN(reg_p0_n497) );
  NAND2_X1 reg_p0_U157 ( .A1(p0_reg[24]), .A2(reg_p0_n503), .ZN(reg_p0_n498)
         );
  NAND2_X1 reg_p0_U156 ( .A1(reg_p0_n496), .A2(reg_p0_n495), .ZN(reg_p0_n242)
         );
  NAND2_X1 reg_p0_U155 ( .A1(p0[23]), .A2(reg_p0_n452), .ZN(reg_p0_n495) );
  NAND2_X1 reg_p0_U154 ( .A1(p0_reg[23]), .A2(reg_p0_n503), .ZN(reg_p0_n496)
         );
  NAND2_X1 reg_p0_U153 ( .A1(reg_p0_n494), .A2(reg_p0_n493), .ZN(reg_p0_n243)
         );
  NAND2_X1 reg_p0_U152 ( .A1(p0[22]), .A2(reg_p0_n452), .ZN(reg_p0_n493) );
  NAND2_X1 reg_p0_U151 ( .A1(p0_reg[22]), .A2(reg_p0_n503), .ZN(reg_p0_n494)
         );
  NAND2_X1 reg_p0_U150 ( .A1(reg_p0_n492), .A2(reg_p0_n491), .ZN(reg_p0_n244)
         );
  NAND2_X1 reg_p0_U149 ( .A1(p0[21]), .A2(reg_p0_n452), .ZN(reg_p0_n491) );
  NAND2_X1 reg_p0_U148 ( .A1(p0_reg[21]), .A2(reg_p0_n503), .ZN(reg_p0_n492)
         );
  NAND2_X1 reg_p0_U147 ( .A1(reg_p0_n490), .A2(reg_p0_n489), .ZN(reg_p0_n245)
         );
  NAND2_X1 reg_p0_U146 ( .A1(p0[20]), .A2(reg_p0_n452), .ZN(reg_p0_n489) );
  NAND2_X1 reg_p0_U145 ( .A1(p0_reg[20]), .A2(reg_p0_n503), .ZN(reg_p0_n490)
         );
  NAND2_X1 reg_p0_U144 ( .A1(reg_p0_n488), .A2(reg_p0_n487), .ZN(reg_p0_n246)
         );
  NAND2_X1 reg_p0_U143 ( .A1(p0[19]), .A2(reg_p0_n452), .ZN(reg_p0_n487) );
  NAND2_X1 reg_p0_U142 ( .A1(p0_reg[19]), .A2(reg_p0_n503), .ZN(reg_p0_n488)
         );
  NAND2_X1 reg_p0_U141 ( .A1(reg_p0_n486), .A2(reg_p0_n485), .ZN(reg_p0_n247)
         );
  NAND2_X1 reg_p0_U140 ( .A1(p0[18]), .A2(reg_p0_n452), .ZN(reg_p0_n485) );
  NAND2_X1 reg_p0_U139 ( .A1(p0_reg[18]), .A2(reg_p0_n503), .ZN(reg_p0_n486)
         );
  NAND2_X1 reg_p0_U138 ( .A1(reg_p0_n484), .A2(reg_p0_n483), .ZN(reg_p0_n248)
         );
  NAND2_X1 reg_p0_U137 ( .A1(p0[17]), .A2(reg_p0_n452), .ZN(reg_p0_n483) );
  NAND2_X1 reg_p0_U136 ( .A1(p0_reg[17]), .A2(reg_p0_n503), .ZN(reg_p0_n484)
         );
  NAND2_X1 reg_p0_U135 ( .A1(reg_p0_n482), .A2(reg_p0_n481), .ZN(reg_p0_n249)
         );
  NAND2_X1 reg_p0_U134 ( .A1(p0[16]), .A2(reg_p0_n452), .ZN(reg_p0_n481) );
  NAND2_X1 reg_p0_U133 ( .A1(p0_reg[16]), .A2(reg_p0_n503), .ZN(reg_p0_n482)
         );
  NAND2_X1 reg_p0_U132 ( .A1(reg_p0_n480), .A2(reg_p0_n479), .ZN(reg_p0_n250)
         );
  NAND2_X1 reg_p0_U131 ( .A1(p0[15]), .A2(reg_p0_n452), .ZN(reg_p0_n479) );
  NAND2_X1 reg_p0_U130 ( .A1(p0_reg[15]), .A2(reg_p0_n503), .ZN(reg_p0_n480)
         );
  NAND2_X1 reg_p0_U129 ( .A1(reg_p0_n478), .A2(reg_p0_n477), .ZN(reg_p0_n251)
         );
  NAND2_X1 reg_p0_U128 ( .A1(p0[14]), .A2(reg_p0_n529), .ZN(reg_p0_n477) );
  NAND2_X1 reg_p0_U127 ( .A1(p0_reg[14]), .A2(reg_p0_n528), .ZN(reg_p0_n478)
         );
  NAND2_X1 reg_p0_U126 ( .A1(reg_p0_n476), .A2(reg_p0_n475), .ZN(reg_p0_n252)
         );
  NAND2_X1 reg_p0_U125 ( .A1(p0[13]), .A2(reg_p0_n452), .ZN(reg_p0_n475) );
  NAND2_X1 reg_p0_U124 ( .A1(p0_reg[13]), .A2(reg_p0_n503), .ZN(reg_p0_n476)
         );
  NAND2_X1 reg_p0_U123 ( .A1(reg_p0_n474), .A2(reg_p0_n473), .ZN(reg_p0_n253)
         );
  NAND2_X1 reg_p0_U122 ( .A1(p0[12]), .A2(reg_p0_n529), .ZN(reg_p0_n473) );
  NAND2_X1 reg_p0_U121 ( .A1(p0_reg[12]), .A2(reg_p0_n528), .ZN(reg_p0_n474)
         );
  NAND2_X1 reg_p0_U120 ( .A1(reg_p0_n472), .A2(reg_p0_n471), .ZN(reg_p0_n254)
         );
  NAND2_X1 reg_p0_U119 ( .A1(p0[11]), .A2(reg_p0_n452), .ZN(reg_p0_n471) );
  NAND2_X1 reg_p0_U118 ( .A1(p0_reg[11]), .A2(reg_p0_n503), .ZN(reg_p0_n472)
         );
  NAND2_X1 reg_p0_U117 ( .A1(reg_p0_n470), .A2(reg_p0_n469), .ZN(reg_p0_n255)
         );
  NAND2_X1 reg_p0_U116 ( .A1(p0[10]), .A2(reg_p0_n529), .ZN(reg_p0_n469) );
  NAND2_X1 reg_p0_U115 ( .A1(p0_reg[10]), .A2(reg_p0_n528), .ZN(reg_p0_n470)
         );
  NAND2_X1 reg_p0_U114 ( .A1(reg_p0_n468), .A2(reg_p0_n467), .ZN(reg_p0_n256)
         );
  NAND2_X1 reg_p0_U113 ( .A1(p0[9]), .A2(reg_p0_n452), .ZN(reg_p0_n467) );
  NAND2_X1 reg_p0_U112 ( .A1(p0_reg[9]), .A2(reg_p0_n503), .ZN(reg_p0_n468) );
  NAND2_X1 reg_p0_U111 ( .A1(reg_p0_n466), .A2(reg_p0_n465), .ZN(reg_p0_n257)
         );
  NAND2_X1 reg_p0_U110 ( .A1(p0[8]), .A2(reg_p0_n529), .ZN(reg_p0_n465) );
  NAND2_X1 reg_p0_U109 ( .A1(p0_reg[8]), .A2(reg_p0_n528), .ZN(reg_p0_n466) );
  NAND2_X1 reg_p0_U108 ( .A1(reg_p0_n464), .A2(reg_p0_n463), .ZN(reg_p0_n258)
         );
  NAND2_X1 reg_p0_U107 ( .A1(p0[7]), .A2(reg_p0_n529), .ZN(reg_p0_n463) );
  NAND2_X1 reg_p0_U106 ( .A1(p0_reg[7]), .A2(reg_p0_n503), .ZN(reg_p0_n464) );
  NAND2_X1 reg_p0_U105 ( .A1(reg_p0_n462), .A2(reg_p0_n461), .ZN(reg_p0_n259)
         );
  NAND2_X1 reg_p0_U104 ( .A1(p0[6]), .A2(reg_p0_n529), .ZN(reg_p0_n461) );
  NAND2_X1 reg_p0_U103 ( .A1(p0_reg[6]), .A2(reg_p0_n528), .ZN(reg_p0_n462) );
  NAND2_X1 reg_p0_U102 ( .A1(reg_p0_n460), .A2(reg_p0_n459), .ZN(reg_p0_n260)
         );
  NAND2_X1 reg_p0_U101 ( .A1(p0[5]), .A2(reg_p0_n452), .ZN(reg_p0_n459) );
  NAND2_X1 reg_p0_U100 ( .A1(p0_reg[5]), .A2(reg_p0_n503), .ZN(reg_p0_n460) );
  INV_X1 reg_p0_U99 ( .A(reg_p0_n457), .ZN(reg_p0_n503) );
  NAND2_X1 reg_p0_U98 ( .A1(reg_p0_n456), .A2(reg_p0_n455), .ZN(reg_p0_n261)
         );
  NAND2_X1 reg_p0_U97 ( .A1(p0[4]), .A2(reg_p0_n529), .ZN(reg_p0_n455) );
  INV_X1 reg_p0_U96 ( .A(reg_p0_n458), .ZN(reg_p0_n529) );
  NAND2_X1 reg_p0_U95 ( .A1(p0_reg[4]), .A2(reg_p0_n528), .ZN(reg_p0_n456) );
  INV_X1 reg_p0_U94 ( .A(reg_p0_n457), .ZN(reg_p0_n528) );
  NAND2_X1 reg_p0_U93 ( .A1(reg_p0_n454), .A2(reg_p0_n453), .ZN(reg_p0_n262)
         );
  NAND2_X1 reg_p0_U92 ( .A1(p0[3]), .A2(reg_p0_n452), .ZN(reg_p0_n453) );
  NAND2_X1 reg_p0_U91 ( .A1(p0_reg[3]), .A2(reg_p0_n451), .ZN(reg_p0_n454) );
  NAND2_X1 reg_p0_U90 ( .A1(reg_p0_n450), .A2(reg_p0_n449), .ZN(reg_p0_n263)
         );
  NAND2_X1 reg_p0_U89 ( .A1(p0[2]), .A2(reg_p0_n452), .ZN(reg_p0_n449) );
  NAND2_X1 reg_p0_U88 ( .A1(p0_reg[2]), .A2(reg_p0_n451), .ZN(reg_p0_n450) );
  NAND2_X1 reg_p0_U87 ( .A1(reg_p0_n448), .A2(reg_p0_n447), .ZN(reg_p0_n264)
         );
  NAND2_X1 reg_p0_U86 ( .A1(p0[1]), .A2(reg_p0_n452), .ZN(reg_p0_n447) );
  NAND2_X1 reg_p0_U85 ( .A1(p0_reg[1]), .A2(reg_p0_n451), .ZN(reg_p0_n448) );
  NAND2_X1 reg_p0_U84 ( .A1(reg_p0_n446), .A2(reg_p0_n445), .ZN(reg_p0_n265)
         );
  NAND2_X1 reg_p0_U83 ( .A1(p0[0]), .A2(reg_p0_n452), .ZN(reg_p0_n445) );
  NAND2_X1 reg_p0_U82 ( .A1(p0_reg[0]), .A2(reg_p0_n451), .ZN(reg_p0_n446) );
  NAND2_X1 reg_p0_U81 ( .A1(reg_p0_n444), .A2(reg_p0_n443), .ZN(reg_p0_n206)
         );
  NAND2_X1 reg_p0_U80 ( .A1(p0[59]), .A2(reg_p0_n452), .ZN(reg_p0_n443) );
  NAND2_X1 reg_p0_U79 ( .A1(p0_reg[59]), .A2(reg_p0_n451), .ZN(reg_p0_n444) );
  NAND2_X1 reg_p0_U78 ( .A1(reg_p0_n442), .A2(reg_p0_n441), .ZN(reg_p0_n207)
         );
  NAND2_X1 reg_p0_U77 ( .A1(p0[58]), .A2(reg_p0_n452), .ZN(reg_p0_n441) );
  NAND2_X1 reg_p0_U76 ( .A1(p0_reg[58]), .A2(reg_p0_n451), .ZN(reg_p0_n442) );
  NAND2_X1 reg_p0_U75 ( .A1(reg_p0_n440), .A2(reg_p0_n439), .ZN(reg_p0_n208)
         );
  NAND2_X1 reg_p0_U74 ( .A1(p0[57]), .A2(reg_p0_n452), .ZN(reg_p0_n439) );
  NAND2_X1 reg_p0_U73 ( .A1(p0_reg[57]), .A2(reg_p0_n451), .ZN(reg_p0_n440) );
  NAND2_X1 reg_p0_U72 ( .A1(reg_p0_n438), .A2(reg_p0_n437), .ZN(reg_p0_n209)
         );
  NAND2_X1 reg_p0_U71 ( .A1(p0[56]), .A2(reg_p0_n452), .ZN(reg_p0_n437) );
  NAND2_X1 reg_p0_U70 ( .A1(p0_reg[56]), .A2(reg_p0_n451), .ZN(reg_p0_n438) );
  NAND2_X1 reg_p0_U69 ( .A1(reg_p0_n436), .A2(reg_p0_n435), .ZN(reg_p0_n210)
         );
  NAND2_X1 reg_p0_U68 ( .A1(p0[55]), .A2(reg_p0_n452), .ZN(reg_p0_n435) );
  NAND2_X1 reg_p0_U67 ( .A1(p0_reg[55]), .A2(reg_p0_n451), .ZN(reg_p0_n436) );
  NAND2_X1 reg_p0_U66 ( .A1(reg_p0_n434), .A2(reg_p0_n433), .ZN(reg_p0_n211)
         );
  NAND2_X1 reg_p0_U65 ( .A1(p0[54]), .A2(reg_p0_n432), .ZN(reg_p0_n433) );
  NAND2_X1 reg_p0_U64 ( .A1(p0_reg[54]), .A2(reg_p0_n451), .ZN(reg_p0_n434) );
  NAND2_X1 reg_p0_U63 ( .A1(reg_p0_n431), .A2(reg_p0_n430), .ZN(reg_p0_n212)
         );
  NAND2_X1 reg_p0_U62 ( .A1(p0[53]), .A2(reg_p0_n432), .ZN(reg_p0_n430) );
  NAND2_X1 reg_p0_U61 ( .A1(p0_reg[53]), .A2(reg_p0_n451), .ZN(reg_p0_n431) );
  NAND2_X1 reg_p0_U60 ( .A1(reg_p0_n429), .A2(reg_p0_n428), .ZN(reg_p0_n213)
         );
  NAND2_X1 reg_p0_U59 ( .A1(p0[52]), .A2(reg_p0_n432), .ZN(reg_p0_n428) );
  NAND2_X1 reg_p0_U58 ( .A1(p0_reg[52]), .A2(reg_p0_n451), .ZN(reg_p0_n429) );
  NAND2_X1 reg_p0_U57 ( .A1(reg_p0_n427), .A2(reg_p0_n426), .ZN(reg_p0_n214)
         );
  NAND2_X1 reg_p0_U56 ( .A1(p0[51]), .A2(reg_p0_n432), .ZN(reg_p0_n426) );
  NAND2_X1 reg_p0_U55 ( .A1(p0_reg[51]), .A2(reg_p0_n451), .ZN(reg_p0_n427) );
  NAND2_X1 reg_p0_U54 ( .A1(reg_p0_n425), .A2(reg_p0_n424), .ZN(reg_p0_n215)
         );
  NAND2_X1 reg_p0_U53 ( .A1(p0[50]), .A2(reg_p0_n432), .ZN(reg_p0_n424) );
  NAND2_X1 reg_p0_U52 ( .A1(p0_reg[50]), .A2(reg_p0_n451), .ZN(reg_p0_n425) );
  NAND2_X1 reg_p0_U51 ( .A1(reg_p0_n423), .A2(reg_p0_n422), .ZN(reg_p0_n216)
         );
  NAND2_X1 reg_p0_U50 ( .A1(p0[49]), .A2(reg_p0_n432), .ZN(reg_p0_n422) );
  NAND2_X1 reg_p0_U49 ( .A1(p0_reg[49]), .A2(reg_p0_n421), .ZN(reg_p0_n423) );
  NAND2_X1 reg_p0_U48 ( .A1(reg_p0_n420), .A2(reg_p0_n419), .ZN(reg_p0_n217)
         );
  NAND2_X1 reg_p0_U47 ( .A1(p0[48]), .A2(reg_p0_n432), .ZN(reg_p0_n419) );
  NAND2_X1 reg_p0_U46 ( .A1(p0_reg[48]), .A2(reg_p0_n421), .ZN(reg_p0_n420) );
  NAND2_X1 reg_p0_U45 ( .A1(reg_p0_n418), .A2(reg_p0_n417), .ZN(reg_p0_n218)
         );
  NAND2_X1 reg_p0_U44 ( .A1(p0[47]), .A2(reg_p0_n432), .ZN(reg_p0_n417) );
  NAND2_X1 reg_p0_U43 ( .A1(p0_reg[47]), .A2(reg_p0_n421), .ZN(reg_p0_n418) );
  NAND2_X1 reg_p0_U42 ( .A1(reg_p0_n416), .A2(reg_p0_n415), .ZN(reg_p0_n219)
         );
  NAND2_X1 reg_p0_U41 ( .A1(p0[46]), .A2(reg_p0_n432), .ZN(reg_p0_n415) );
  NAND2_X1 reg_p0_U40 ( .A1(p0_reg[46]), .A2(reg_p0_n421), .ZN(reg_p0_n416) );
  NAND2_X1 reg_p0_U39 ( .A1(reg_p0_n414), .A2(reg_p0_n413), .ZN(reg_p0_n220)
         );
  NAND2_X1 reg_p0_U38 ( .A1(p0[45]), .A2(reg_p0_n432), .ZN(reg_p0_n413) );
  NAND2_X1 reg_p0_U37 ( .A1(p0_reg[45]), .A2(reg_p0_n421), .ZN(reg_p0_n414) );
  NAND2_X1 reg_p0_U36 ( .A1(reg_p0_n412), .A2(reg_p0_n411), .ZN(reg_p0_n221)
         );
  NAND2_X1 reg_p0_U35 ( .A1(p0[44]), .A2(reg_p0_n432), .ZN(reg_p0_n411) );
  NAND2_X1 reg_p0_U34 ( .A1(p0_reg[44]), .A2(reg_p0_n421), .ZN(reg_p0_n412) );
  NAND2_X1 reg_p0_U33 ( .A1(reg_p0_n410), .A2(reg_p0_n409), .ZN(reg_p0_n222)
         );
  NAND2_X1 reg_p0_U32 ( .A1(p0[43]), .A2(reg_p0_n432), .ZN(reg_p0_n409) );
  NAND2_X1 reg_p0_U31 ( .A1(p0_reg[43]), .A2(reg_p0_n421), .ZN(reg_p0_n410) );
  NAND2_X1 reg_p0_U30 ( .A1(reg_p0_n408), .A2(reg_p0_n407), .ZN(reg_p0_n223)
         );
  NAND2_X1 reg_p0_U29 ( .A1(p0[42]), .A2(reg_p0_n432), .ZN(reg_p0_n407) );
  NAND2_X1 reg_p0_U28 ( .A1(p0_reg[42]), .A2(reg_p0_n421), .ZN(reg_p0_n408) );
  NAND2_X1 reg_p0_U27 ( .A1(reg_p0_n406), .A2(reg_p0_n405), .ZN(reg_p0_n224)
         );
  NAND2_X1 reg_p0_U26 ( .A1(p0[41]), .A2(reg_p0_n432), .ZN(reg_p0_n405) );
  NAND2_X1 reg_p0_U25 ( .A1(p0_reg[41]), .A2(reg_p0_n421), .ZN(reg_p0_n406) );
  NAND2_X1 reg_p0_U24 ( .A1(reg_p0_n404), .A2(reg_p0_n403), .ZN(reg_p0_n225)
         );
  NAND2_X1 reg_p0_U23 ( .A1(p0[40]), .A2(reg_p0_n432), .ZN(reg_p0_n403) );
  NAND2_X1 reg_p0_U22 ( .A1(p0_reg[40]), .A2(reg_p0_n451), .ZN(reg_p0_n404) );
  NAND2_X1 reg_p0_U21 ( .A1(reg_p0_n402), .A2(reg_p0_n401), .ZN(reg_p0_n226)
         );
  NAND2_X1 reg_p0_U20 ( .A1(p0[39]), .A2(reg_p0_n432), .ZN(reg_p0_n401) );
  NAND2_X1 reg_p0_U19 ( .A1(p0_reg[39]), .A2(reg_p0_n451), .ZN(reg_p0_n402) );
  NAND2_X1 reg_p0_U18 ( .A1(reg_p0_n400), .A2(reg_p0_n399), .ZN(reg_p0_n227)
         );
  NAND2_X1 reg_p0_U17 ( .A1(p0[38]), .A2(reg_p0_n432), .ZN(reg_p0_n399) );
  NAND2_X1 reg_p0_U16 ( .A1(p0_reg[38]), .A2(reg_p0_n451), .ZN(reg_p0_n400) );
  NAND2_X1 reg_p0_U15 ( .A1(reg_p0_n398), .A2(reg_p0_n397), .ZN(reg_p0_n228)
         );
  NAND2_X1 reg_p0_U14 ( .A1(p0[37]), .A2(reg_p0_n432), .ZN(reg_p0_n397) );
  NAND2_X1 reg_p0_U13 ( .A1(p0_reg[37]), .A2(reg_p0_n451), .ZN(reg_p0_n398) );
  NAND2_X1 reg_p0_U12 ( .A1(reg_p0_n396), .A2(reg_p0_n395), .ZN(reg_p0_n229)
         );
  NAND2_X1 reg_p0_U11 ( .A1(reg_p0_n451), .A2(p0_reg[36]), .ZN(reg_p0_n395) );
  INV_X1 reg_p0_U10 ( .A(reg_p0_n457), .ZN(reg_p0_n451) );
  INV_X1 reg_p0_U9 ( .A(reg_p0_n421), .ZN(reg_p0_n457) );
  NAND2_X1 reg_p0_U8 ( .A1(reg_p0_n432), .A2(p0[36]), .ZN(reg_p0_n396) );
  INV_X1 reg_p0_U7 ( .A(reg_p0_n458), .ZN(reg_p0_n432) );
  INV_X1 reg_p0_U6 ( .A(reg_p0_n452), .ZN(reg_p0_n458) );
  NOR2_X4 reg_p0_U5 ( .A1(rst), .A2(reg_p0_n394), .ZN(reg_p0_n452) );
  INV_X1 reg_p0_U4 ( .A(en_sig), .ZN(reg_p0_n394) );
  NOR2_X1 reg_p0_U3 ( .A1(rst), .A2(en_sig), .ZN(reg_p0_n421) );
  DFF_X1 reg_p0_s_current_state_reg_0_ ( .D(reg_p0_n265), .CK(clk), .Q(
        p0_reg[0]) );
  DFF_X1 reg_p0_s_current_state_reg_1_ ( .D(reg_p0_n264), .CK(clk), .Q(
        p0_reg[1]) );
  DFF_X1 reg_p0_s_current_state_reg_2_ ( .D(reg_p0_n263), .CK(clk), .Q(
        p0_reg[2]) );
  DFF_X1 reg_p0_s_current_state_reg_3_ ( .D(reg_p0_n262), .CK(clk), .Q(
        p0_reg[3]) );
  DFF_X1 reg_p0_s_current_state_reg_4_ ( .D(reg_p0_n261), .CK(clk), .Q(
        p0_reg[4]) );
  DFF_X1 reg_p0_s_current_state_reg_5_ ( .D(reg_p0_n260), .CK(clk), .Q(
        p0_reg[5]) );
  DFF_X1 reg_p0_s_current_state_reg_6_ ( .D(reg_p0_n259), .CK(clk), .Q(
        p0_reg[6]) );
  DFF_X1 reg_p0_s_current_state_reg_7_ ( .D(reg_p0_n258), .CK(clk), .Q(
        p0_reg[7]) );
  DFF_X1 reg_p0_s_current_state_reg_8_ ( .D(reg_p0_n257), .CK(clk), .Q(
        p0_reg[8]) );
  DFF_X1 reg_p0_s_current_state_reg_9_ ( .D(reg_p0_n256), .CK(clk), .Q(
        p0_reg[9]) );
  DFF_X1 reg_p0_s_current_state_reg_10_ ( .D(reg_p0_n255), .CK(clk), .Q(
        p0_reg[10]) );
  DFF_X1 reg_p0_s_current_state_reg_11_ ( .D(reg_p0_n254), .CK(clk), .Q(
        p0_reg[11]) );
  DFF_X1 reg_p0_s_current_state_reg_12_ ( .D(reg_p0_n253), .CK(clk), .Q(
        p0_reg[12]) );
  DFF_X1 reg_p0_s_current_state_reg_13_ ( .D(reg_p0_n252), .CK(clk), .Q(
        p0_reg[13]) );
  DFF_X1 reg_p0_s_current_state_reg_14_ ( .D(reg_p0_n251), .CK(clk), .Q(
        p0_reg[14]) );
  DFF_X1 reg_p0_s_current_state_reg_15_ ( .D(reg_p0_n250), .CK(clk), .Q(
        p0_reg[15]) );
  DFF_X1 reg_p0_s_current_state_reg_16_ ( .D(reg_p0_n249), .CK(clk), .Q(
        p0_reg[16]) );
  DFF_X1 reg_p0_s_current_state_reg_17_ ( .D(reg_p0_n248), .CK(clk), .Q(
        p0_reg[17]) );
  DFF_X1 reg_p0_s_current_state_reg_18_ ( .D(reg_p0_n247), .CK(clk), .Q(
        p0_reg[18]) );
  DFF_X1 reg_p0_s_current_state_reg_19_ ( .D(reg_p0_n246), .CK(clk), .Q(
        p0_reg[19]) );
  DFF_X1 reg_p0_s_current_state_reg_20_ ( .D(reg_p0_n245), .CK(clk), .Q(
        p0_reg[20]) );
  DFF_X1 reg_p0_s_current_state_reg_21_ ( .D(reg_p0_n244), .CK(clk), .Q(
        p0_reg[21]) );
  DFF_X1 reg_p0_s_current_state_reg_22_ ( .D(reg_p0_n243), .CK(clk), .Q(
        p0_reg[22]) );
  DFF_X1 reg_p0_s_current_state_reg_23_ ( .D(reg_p0_n242), .CK(clk), .Q(
        p0_reg[23]) );
  DFF_X1 reg_p0_s_current_state_reg_24_ ( .D(reg_p0_n241), .CK(clk), .Q(
        p0_reg[24]) );
  DFF_X1 reg_p0_s_current_state_reg_25_ ( .D(reg_p0_n240), .CK(clk), .Q(
        p0_reg[25]) );
  DFF_X1 reg_p0_s_current_state_reg_26_ ( .D(reg_p0_n239), .CK(clk), .Q(
        p0_reg[26]) );
  DFF_X1 reg_p0_s_current_state_reg_27_ ( .D(reg_p0_n238), .CK(clk), .Q(
        p0_reg[27]) );
  DFF_X1 reg_p0_s_current_state_reg_28_ ( .D(reg_p0_n237), .CK(clk), .Q(
        p0_reg[28]) );
  DFF_X1 reg_p0_s_current_state_reg_29_ ( .D(reg_p0_n236), .CK(clk), .Q(
        p0_reg[29]) );
  DFF_X1 reg_p0_s_current_state_reg_30_ ( .D(reg_p0_n235), .CK(clk), .Q(
        p0_reg[30]) );
  DFF_X1 reg_p0_s_current_state_reg_31_ ( .D(reg_p0_n234), .CK(clk), .Q(
        p0_reg[31]) );
  DFF_X1 reg_p0_s_current_state_reg_32_ ( .D(reg_p0_n233), .CK(clk), .Q(
        p0_reg[32]) );
  DFF_X1 reg_p0_s_current_state_reg_33_ ( .D(reg_p0_n232), .CK(clk), .Q(
        p0_reg[33]) );
  DFF_X1 reg_p0_s_current_state_reg_34_ ( .D(reg_p0_n231), .CK(clk), .Q(
        p0_reg[34]) );
  DFF_X1 reg_p0_s_current_state_reg_35_ ( .D(reg_p0_n230), .CK(clk), .Q(
        p0_reg[35]) );
  DFF_X1 reg_p0_s_current_state_reg_36_ ( .D(reg_p0_n229), .CK(clk), .Q(
        p0_reg[36]) );
  DFF_X1 reg_p0_s_current_state_reg_37_ ( .D(reg_p0_n228), .CK(clk), .Q(
        p0_reg[37]) );
  DFF_X1 reg_p0_s_current_state_reg_38_ ( .D(reg_p0_n227), .CK(clk), .Q(
        p0_reg[38]) );
  DFF_X1 reg_p0_s_current_state_reg_39_ ( .D(reg_p0_n226), .CK(clk), .Q(
        p0_reg[39]) );
  DFF_X1 reg_p0_s_current_state_reg_40_ ( .D(reg_p0_n225), .CK(clk), .Q(
        p0_reg[40]) );
  DFF_X1 reg_p0_s_current_state_reg_41_ ( .D(reg_p0_n224), .CK(clk), .Q(
        p0_reg[41]) );
  DFF_X1 reg_p0_s_current_state_reg_42_ ( .D(reg_p0_n223), .CK(clk), .Q(
        p0_reg[42]) );
  DFF_X1 reg_p0_s_current_state_reg_43_ ( .D(reg_p0_n222), .CK(clk), .Q(
        p0_reg[43]) );
  DFF_X1 reg_p0_s_current_state_reg_44_ ( .D(reg_p0_n221), .CK(clk), .Q(
        p0_reg[44]) );
  DFF_X1 reg_p0_s_current_state_reg_45_ ( .D(reg_p0_n220), .CK(clk), .Q(
        p0_reg[45]) );
  DFF_X1 reg_p0_s_current_state_reg_46_ ( .D(reg_p0_n219), .CK(clk), .Q(
        p0_reg[46]) );
  DFF_X1 reg_p0_s_current_state_reg_47_ ( .D(reg_p0_n218), .CK(clk), .Q(
        p0_reg[47]) );
  DFF_X1 reg_p0_s_current_state_reg_48_ ( .D(reg_p0_n217), .CK(clk), .Q(
        p0_reg[48]) );
  DFF_X1 reg_p0_s_current_state_reg_49_ ( .D(reg_p0_n216), .CK(clk), .Q(
        p0_reg[49]) );
  DFF_X1 reg_p0_s_current_state_reg_50_ ( .D(reg_p0_n215), .CK(clk), .Q(
        p0_reg[50]) );
  DFF_X1 reg_p0_s_current_state_reg_51_ ( .D(reg_p0_n214), .CK(clk), .Q(
        p0_reg[51]) );
  DFF_X1 reg_p0_s_current_state_reg_52_ ( .D(reg_p0_n213), .CK(clk), .Q(
        p0_reg[52]) );
  DFF_X1 reg_p0_s_current_state_reg_53_ ( .D(reg_p0_n212), .CK(clk), .Q(
        p0_reg[53]) );
  DFF_X1 reg_p0_s_current_state_reg_54_ ( .D(reg_p0_n211), .CK(clk), .Q(
        p0_reg[54]) );
  DFF_X1 reg_p0_s_current_state_reg_55_ ( .D(reg_p0_n210), .CK(clk), .Q(
        p0_reg[55]) );
  DFF_X1 reg_p0_s_current_state_reg_56_ ( .D(reg_p0_n209), .CK(clk), .Q(
        p0_reg[56]) );
  DFF_X1 reg_p0_s_current_state_reg_57_ ( .D(reg_p0_n208), .CK(clk), .Q(
        p0_reg[57]) );
  DFF_X1 reg_p0_s_current_state_reg_58_ ( .D(reg_p0_n207), .CK(clk), .Q(
        p0_reg[58]) );
  DFF_X1 reg_p0_s_current_state_reg_59_ ( .D(reg_p0_n206), .CK(clk), .Q(
        p0_reg[59]) );
  DFF_X1 reg_p0_s_current_state_reg_60_ ( .D(reg_p0_n205), .CK(clk), .Q(
        p0_reg[60]) );
  DFF_X1 reg_p0_s_current_state_reg_61_ ( .D(reg_p0_n204), .CK(clk), .Q(
        p0_reg[61]) );
  DFF_X1 reg_p0_s_current_state_reg_62_ ( .D(reg_p0_n203), .CK(clk), .Q(
        p0_reg[62]) );
  DFF_X1 reg_p0_s_current_state_reg_63_ ( .D(reg_p0_n202), .CK(clk), .Q(
        p0_reg[63]) );
  NAND2_X1 reg_p1_U205 ( .A1(reg_p1_n532), .A2(reg_p1_n531), .ZN(reg_p1_n202)
         );
  NAND2_X1 reg_p1_U204 ( .A1(p1[63]), .A2(reg_p1_n530), .ZN(reg_p1_n531) );
  NAND2_X1 reg_p1_U203 ( .A1(init_y[63]), .A2(reg_p1_n529), .ZN(reg_p1_n532)
         );
  NAND2_X1 reg_p1_U202 ( .A1(reg_p1_n528), .A2(reg_p1_n527), .ZN(reg_p1_n203)
         );
  NAND2_X1 reg_p1_U201 ( .A1(p1[62]), .A2(reg_p1_n530), .ZN(reg_p1_n527) );
  NAND2_X1 reg_p1_U200 ( .A1(init_y[62]), .A2(reg_p1_n529), .ZN(reg_p1_n528)
         );
  NAND2_X1 reg_p1_U199 ( .A1(reg_p1_n526), .A2(reg_p1_n525), .ZN(reg_p1_n204)
         );
  NAND2_X1 reg_p1_U198 ( .A1(p1[61]), .A2(reg_p1_n530), .ZN(reg_p1_n525) );
  NAND2_X1 reg_p1_U197 ( .A1(init_y[61]), .A2(reg_p1_n529), .ZN(reg_p1_n526)
         );
  NAND2_X1 reg_p1_U196 ( .A1(reg_p1_n524), .A2(reg_p1_n523), .ZN(reg_p1_n205)
         );
  NAND2_X1 reg_p1_U195 ( .A1(p1[60]), .A2(reg_p1_n530), .ZN(reg_p1_n523) );
  NAND2_X1 reg_p1_U194 ( .A1(init_y[60]), .A2(reg_p1_n529), .ZN(reg_p1_n524)
         );
  NAND2_X1 reg_p1_U193 ( .A1(reg_p1_n522), .A2(reg_p1_n521), .ZN(reg_p1_n230)
         );
  NAND2_X1 reg_p1_U192 ( .A1(p1[35]), .A2(reg_p1_n530), .ZN(reg_p1_n521) );
  NAND2_X1 reg_p1_U191 ( .A1(init_y[51]), .A2(reg_p1_n529), .ZN(reg_p1_n522)
         );
  NAND2_X1 reg_p1_U190 ( .A1(reg_p1_n520), .A2(reg_p1_n519), .ZN(reg_p1_n231)
         );
  NAND2_X1 reg_p1_U189 ( .A1(p1[34]), .A2(reg_p1_n530), .ZN(reg_p1_n519) );
  NAND2_X1 reg_p1_U188 ( .A1(init_y[50]), .A2(reg_p1_n529), .ZN(reg_p1_n520)
         );
  NAND2_X1 reg_p1_U187 ( .A1(reg_p1_n518), .A2(reg_p1_n517), .ZN(reg_p1_n232)
         );
  NAND2_X1 reg_p1_U186 ( .A1(p1[33]), .A2(reg_p1_n530), .ZN(reg_p1_n517) );
  NAND2_X1 reg_p1_U185 ( .A1(init_y[49]), .A2(reg_p1_n529), .ZN(reg_p1_n518)
         );
  NAND2_X1 reg_p1_U184 ( .A1(reg_p1_n516), .A2(reg_p1_n515), .ZN(reg_p1_n233)
         );
  NAND2_X1 reg_p1_U183 ( .A1(p1[32]), .A2(reg_p1_n530), .ZN(reg_p1_n515) );
  NAND2_X1 reg_p1_U182 ( .A1(init_y[48]), .A2(reg_p1_n529), .ZN(reg_p1_n516)
         );
  NAND2_X1 reg_p1_U181 ( .A1(reg_p1_n514), .A2(reg_p1_n513), .ZN(reg_p1_n234)
         );
  NAND2_X1 reg_p1_U180 ( .A1(p1[31]), .A2(reg_p1_n530), .ZN(reg_p1_n513) );
  NAND2_X1 reg_p1_U179 ( .A1(init_y[31]), .A2(reg_p1_n529), .ZN(reg_p1_n514)
         );
  NAND2_X1 reg_p1_U178 ( .A1(reg_p1_n512), .A2(reg_p1_n511), .ZN(reg_p1_n235)
         );
  NAND2_X1 reg_p1_U177 ( .A1(p1[30]), .A2(reg_p1_n530), .ZN(reg_p1_n511) );
  NAND2_X1 reg_p1_U176 ( .A1(init_y[30]), .A2(reg_p1_n529), .ZN(reg_p1_n512)
         );
  NAND2_X1 reg_p1_U175 ( .A1(reg_p1_n510), .A2(reg_p1_n509), .ZN(reg_p1_n236)
         );
  NAND2_X1 reg_p1_U174 ( .A1(p1[29]), .A2(reg_p1_n530), .ZN(reg_p1_n509) );
  NAND2_X1 reg_p1_U173 ( .A1(init_y[29]), .A2(reg_p1_n529), .ZN(reg_p1_n510)
         );
  NAND2_X1 reg_p1_U172 ( .A1(reg_p1_n508), .A2(reg_p1_n507), .ZN(reg_p1_n237)
         );
  NAND2_X1 reg_p1_U171 ( .A1(p1[28]), .A2(reg_p1_n530), .ZN(reg_p1_n507) );
  NAND2_X1 reg_p1_U170 ( .A1(init_y[28]), .A2(reg_p1_n529), .ZN(reg_p1_n508)
         );
  NAND2_X1 reg_p1_U169 ( .A1(reg_p1_n506), .A2(reg_p1_n505), .ZN(reg_p1_n238)
         );
  NAND2_X1 reg_p1_U168 ( .A1(p1[27]), .A2(reg_p1_n504), .ZN(reg_p1_n505) );
  NAND2_X1 reg_p1_U167 ( .A1(init_y[11]), .A2(reg_p1_n503), .ZN(reg_p1_n506)
         );
  NAND2_X1 reg_p1_U166 ( .A1(reg_p1_n502), .A2(reg_p1_n501), .ZN(reg_p1_n239)
         );
  NAND2_X1 reg_p1_U165 ( .A1(p1[26]), .A2(reg_p1_n504), .ZN(reg_p1_n501) );
  NAND2_X1 reg_p1_U164 ( .A1(init_y[10]), .A2(reg_p1_n503), .ZN(reg_p1_n502)
         );
  NAND2_X1 reg_p1_U163 ( .A1(reg_p1_n500), .A2(reg_p1_n499), .ZN(reg_p1_n240)
         );
  NAND2_X1 reg_p1_U162 ( .A1(p1[25]), .A2(reg_p1_n504), .ZN(reg_p1_n499) );
  NAND2_X1 reg_p1_U161 ( .A1(init_y[9]), .A2(reg_p1_n503), .ZN(reg_p1_n500) );
  NAND2_X1 reg_p1_U160 ( .A1(reg_p1_n498), .A2(reg_p1_n497), .ZN(reg_p1_n241)
         );
  NAND2_X1 reg_p1_U159 ( .A1(p1[24]), .A2(reg_p1_n504), .ZN(reg_p1_n497) );
  NAND2_X1 reg_p1_U158 ( .A1(init_y[8]), .A2(reg_p1_n503), .ZN(reg_p1_n498) );
  NAND2_X1 reg_p1_U157 ( .A1(reg_p1_n496), .A2(reg_p1_n495), .ZN(reg_p1_n242)
         );
  NAND2_X1 reg_p1_U156 ( .A1(p1[23]), .A2(reg_p1_n504), .ZN(reg_p1_n495) );
  NAND2_X1 reg_p1_U155 ( .A1(init_y[55]), .A2(reg_p1_n503), .ZN(reg_p1_n496)
         );
  NAND2_X1 reg_p1_U154 ( .A1(reg_p1_n494), .A2(reg_p1_n493), .ZN(reg_p1_n243)
         );
  NAND2_X1 reg_p1_U153 ( .A1(p1[22]), .A2(reg_p1_n504), .ZN(reg_p1_n493) );
  NAND2_X1 reg_p1_U152 ( .A1(init_y[54]), .A2(reg_p1_n503), .ZN(reg_p1_n494)
         );
  NAND2_X1 reg_p1_U151 ( .A1(reg_p1_n492), .A2(reg_p1_n491), .ZN(reg_p1_n244)
         );
  NAND2_X1 reg_p1_U150 ( .A1(p1[21]), .A2(reg_p1_n504), .ZN(reg_p1_n491) );
  NAND2_X1 reg_p1_U149 ( .A1(init_y[53]), .A2(reg_p1_n503), .ZN(reg_p1_n492)
         );
  NAND2_X1 reg_p1_U148 ( .A1(reg_p1_n490), .A2(reg_p1_n489), .ZN(reg_p1_n245)
         );
  NAND2_X1 reg_p1_U147 ( .A1(p1[20]), .A2(reg_p1_n504), .ZN(reg_p1_n489) );
  NAND2_X1 reg_p1_U146 ( .A1(init_y[52]), .A2(reg_p1_n503), .ZN(reg_p1_n490)
         );
  NAND2_X1 reg_p1_U145 ( .A1(reg_p1_n488), .A2(reg_p1_n487), .ZN(reg_p1_n246)
         );
  NAND2_X1 reg_p1_U144 ( .A1(p1[19]), .A2(reg_p1_n504), .ZN(reg_p1_n487) );
  NAND2_X1 reg_p1_U143 ( .A1(init_y[35]), .A2(reg_p1_n503), .ZN(reg_p1_n488)
         );
  NAND2_X1 reg_p1_U142 ( .A1(reg_p1_n486), .A2(reg_p1_n485), .ZN(reg_p1_n247)
         );
  NAND2_X1 reg_p1_U141 ( .A1(p1[18]), .A2(reg_p1_n504), .ZN(reg_p1_n485) );
  NAND2_X1 reg_p1_U140 ( .A1(init_y[34]), .A2(reg_p1_n503), .ZN(reg_p1_n486)
         );
  NAND2_X1 reg_p1_U139 ( .A1(reg_p1_n484), .A2(reg_p1_n483), .ZN(reg_p1_n248)
         );
  NAND2_X1 reg_p1_U138 ( .A1(p1[17]), .A2(reg_p1_n504), .ZN(reg_p1_n483) );
  NAND2_X1 reg_p1_U137 ( .A1(init_y[33]), .A2(reg_p1_n503), .ZN(reg_p1_n484)
         );
  NAND2_X1 reg_p1_U136 ( .A1(reg_p1_n482), .A2(reg_p1_n481), .ZN(reg_p1_n249)
         );
  NAND2_X1 reg_p1_U135 ( .A1(p1[16]), .A2(reg_p1_n504), .ZN(reg_p1_n481) );
  NAND2_X1 reg_p1_U134 ( .A1(init_y[32]), .A2(reg_p1_n503), .ZN(reg_p1_n482)
         );
  NAND2_X1 reg_p1_U133 ( .A1(reg_p1_n480), .A2(reg_p1_n479), .ZN(reg_p1_n250)
         );
  NAND2_X1 reg_p1_U132 ( .A1(p1[15]), .A2(reg_p1_n504), .ZN(reg_p1_n479) );
  NAND2_X1 reg_p1_U131 ( .A1(init_y[15]), .A2(reg_p1_n503), .ZN(reg_p1_n480)
         );
  NAND2_X1 reg_p1_U130 ( .A1(reg_p1_n478), .A2(reg_p1_n477), .ZN(reg_p1_n251)
         );
  NAND2_X1 reg_p1_U129 ( .A1(p1[14]), .A2(reg_p1_n530), .ZN(reg_p1_n477) );
  NAND2_X1 reg_p1_U128 ( .A1(init_y[14]), .A2(reg_p1_n529), .ZN(reg_p1_n478)
         );
  NAND2_X1 reg_p1_U127 ( .A1(reg_p1_n476), .A2(reg_p1_n475), .ZN(reg_p1_n252)
         );
  NAND2_X1 reg_p1_U126 ( .A1(p1[13]), .A2(reg_p1_n504), .ZN(reg_p1_n475) );
  NAND2_X1 reg_p1_U125 ( .A1(init_y[13]), .A2(reg_p1_n503), .ZN(reg_p1_n476)
         );
  NAND2_X1 reg_p1_U124 ( .A1(reg_p1_n474), .A2(reg_p1_n473), .ZN(reg_p1_n253)
         );
  NAND2_X1 reg_p1_U123 ( .A1(p1[12]), .A2(reg_p1_n530), .ZN(reg_p1_n473) );
  NAND2_X1 reg_p1_U122 ( .A1(init_y[12]), .A2(reg_p1_n529), .ZN(reg_p1_n474)
         );
  NAND2_X1 reg_p1_U121 ( .A1(reg_p1_n472), .A2(reg_p1_n471), .ZN(reg_p1_n254)
         );
  NAND2_X1 reg_p1_U120 ( .A1(p1[11]), .A2(reg_p1_n504), .ZN(reg_p1_n471) );
  NAND2_X1 reg_p1_U119 ( .A1(init_y[59]), .A2(reg_p1_n503), .ZN(reg_p1_n472)
         );
  NAND2_X1 reg_p1_U118 ( .A1(reg_p1_n470), .A2(reg_p1_n469), .ZN(reg_p1_n255)
         );
  NAND2_X1 reg_p1_U117 ( .A1(p1[10]), .A2(reg_p1_n530), .ZN(reg_p1_n469) );
  NAND2_X1 reg_p1_U116 ( .A1(init_y[58]), .A2(reg_p1_n529), .ZN(reg_p1_n470)
         );
  NAND2_X1 reg_p1_U115 ( .A1(reg_p1_n468), .A2(reg_p1_n467), .ZN(reg_p1_n256)
         );
  NAND2_X1 reg_p1_U114 ( .A1(p1[9]), .A2(reg_p1_n504), .ZN(reg_p1_n467) );
  NAND2_X1 reg_p1_U113 ( .A1(init_y[57]), .A2(reg_p1_n503), .ZN(reg_p1_n468)
         );
  NAND2_X1 reg_p1_U112 ( .A1(reg_p1_n466), .A2(reg_p1_n465), .ZN(reg_p1_n257)
         );
  NAND2_X1 reg_p1_U111 ( .A1(p1[8]), .A2(reg_p1_n530), .ZN(reg_p1_n465) );
  NAND2_X1 reg_p1_U110 ( .A1(init_y[56]), .A2(reg_p1_n529), .ZN(reg_p1_n466)
         );
  NAND2_X1 reg_p1_U109 ( .A1(reg_p1_n464), .A2(reg_p1_n463), .ZN(reg_p1_n258)
         );
  NAND2_X1 reg_p1_U108 ( .A1(p1[7]), .A2(reg_p1_n504), .ZN(reg_p1_n463) );
  NAND2_X1 reg_p1_U107 ( .A1(init_y[39]), .A2(reg_p1_n503), .ZN(reg_p1_n464)
         );
  NAND2_X1 reg_p1_U106 ( .A1(reg_p1_n462), .A2(reg_p1_n461), .ZN(reg_p1_n259)
         );
  NAND2_X1 reg_p1_U105 ( .A1(p1[6]), .A2(reg_p1_n530), .ZN(reg_p1_n461) );
  NAND2_X1 reg_p1_U104 ( .A1(init_y[38]), .A2(reg_p1_n529), .ZN(reg_p1_n462)
         );
  NAND2_X1 reg_p1_U103 ( .A1(reg_p1_n460), .A2(reg_p1_n459), .ZN(reg_p1_n260)
         );
  NAND2_X1 reg_p1_U102 ( .A1(p1[5]), .A2(reg_p1_n504), .ZN(reg_p1_n459) );
  INV_X1 reg_p1_U101 ( .A(reg_p1_n458), .ZN(reg_p1_n504) );
  NAND2_X1 reg_p1_U100 ( .A1(init_y[37]), .A2(reg_p1_n503), .ZN(reg_p1_n460)
         );
  INV_X1 reg_p1_U99 ( .A(reg_p1_n457), .ZN(reg_p1_n503) );
  NAND2_X1 reg_p1_U98 ( .A1(reg_p1_n456), .A2(reg_p1_n455), .ZN(reg_p1_n261)
         );
  NAND2_X1 reg_p1_U97 ( .A1(p1[4]), .A2(reg_p1_n530), .ZN(reg_p1_n455) );
  INV_X1 reg_p1_U96 ( .A(reg_p1_n458), .ZN(reg_p1_n530) );
  NAND2_X1 reg_p1_U95 ( .A1(init_y[36]), .A2(reg_p1_n529), .ZN(reg_p1_n456) );
  INV_X1 reg_p1_U94 ( .A(reg_p1_n457), .ZN(reg_p1_n529) );
  NAND2_X1 reg_p1_U93 ( .A1(reg_p1_n454), .A2(reg_p1_n453), .ZN(reg_p1_n262)
         );
  NAND2_X1 reg_p1_U92 ( .A1(p1[3]), .A2(reg_p1_n452), .ZN(reg_p1_n453) );
  NAND2_X1 reg_p1_U91 ( .A1(init_y[19]), .A2(reg_p1_n451), .ZN(reg_p1_n454) );
  NAND2_X1 reg_p1_U90 ( .A1(reg_p1_n450), .A2(reg_p1_n449), .ZN(reg_p1_n263)
         );
  NAND2_X1 reg_p1_U89 ( .A1(p1[2]), .A2(reg_p1_n452), .ZN(reg_p1_n449) );
  NAND2_X1 reg_p1_U88 ( .A1(init_y[18]), .A2(reg_p1_n451), .ZN(reg_p1_n450) );
  NAND2_X1 reg_p1_U87 ( .A1(reg_p1_n448), .A2(reg_p1_n447), .ZN(reg_p1_n264)
         );
  NAND2_X1 reg_p1_U86 ( .A1(p1[1]), .A2(reg_p1_n452), .ZN(reg_p1_n447) );
  NAND2_X1 reg_p1_U85 ( .A1(init_y[17]), .A2(reg_p1_n451), .ZN(reg_p1_n448) );
  NAND2_X1 reg_p1_U84 ( .A1(reg_p1_n446), .A2(reg_p1_n445), .ZN(reg_p1_n265)
         );
  NAND2_X1 reg_p1_U83 ( .A1(p1[0]), .A2(reg_p1_n452), .ZN(reg_p1_n445) );
  NAND2_X1 reg_p1_U82 ( .A1(init_y[16]), .A2(reg_p1_n451), .ZN(reg_p1_n446) );
  NAND2_X1 reg_p1_U81 ( .A1(reg_p1_n444), .A2(reg_p1_n443), .ZN(reg_p1_n206)
         );
  NAND2_X1 reg_p1_U80 ( .A1(p1[59]), .A2(reg_p1_n452), .ZN(reg_p1_n443) );
  NAND2_X1 reg_p1_U79 ( .A1(init_y[43]), .A2(reg_p1_n451), .ZN(reg_p1_n444) );
  NAND2_X1 reg_p1_U78 ( .A1(reg_p1_n442), .A2(reg_p1_n441), .ZN(reg_p1_n207)
         );
  NAND2_X1 reg_p1_U77 ( .A1(p1[58]), .A2(reg_p1_n452), .ZN(reg_p1_n441) );
  NAND2_X1 reg_p1_U76 ( .A1(init_y[42]), .A2(reg_p1_n451), .ZN(reg_p1_n442) );
  NAND2_X1 reg_p1_U75 ( .A1(reg_p1_n440), .A2(reg_p1_n439), .ZN(reg_p1_n208)
         );
  NAND2_X1 reg_p1_U74 ( .A1(p1[57]), .A2(reg_p1_n452), .ZN(reg_p1_n439) );
  NAND2_X1 reg_p1_U73 ( .A1(init_y[41]), .A2(reg_p1_n451), .ZN(reg_p1_n440) );
  NAND2_X1 reg_p1_U72 ( .A1(reg_p1_n438), .A2(reg_p1_n437), .ZN(reg_p1_n209)
         );
  NAND2_X1 reg_p1_U71 ( .A1(p1[56]), .A2(reg_p1_n452), .ZN(reg_p1_n437) );
  NAND2_X1 reg_p1_U70 ( .A1(init_y[40]), .A2(reg_p1_n451), .ZN(reg_p1_n438) );
  NAND2_X1 reg_p1_U69 ( .A1(reg_p1_n436), .A2(reg_p1_n435), .ZN(reg_p1_n210)
         );
  NAND2_X1 reg_p1_U68 ( .A1(p1[55]), .A2(reg_p1_n452), .ZN(reg_p1_n435) );
  NAND2_X1 reg_p1_U67 ( .A1(init_y[23]), .A2(reg_p1_n451), .ZN(reg_p1_n436) );
  NAND2_X1 reg_p1_U66 ( .A1(reg_p1_n434), .A2(reg_p1_n433), .ZN(reg_p1_n211)
         );
  NAND2_X1 reg_p1_U65 ( .A1(p1[54]), .A2(reg_p1_n432), .ZN(reg_p1_n433) );
  NAND2_X1 reg_p1_U64 ( .A1(init_y[22]), .A2(reg_p1_n451), .ZN(reg_p1_n434) );
  NAND2_X1 reg_p1_U63 ( .A1(reg_p1_n431), .A2(reg_p1_n430), .ZN(reg_p1_n212)
         );
  NAND2_X1 reg_p1_U62 ( .A1(p1[53]), .A2(reg_p1_n432), .ZN(reg_p1_n430) );
  NAND2_X1 reg_p1_U61 ( .A1(init_y[21]), .A2(reg_p1_n451), .ZN(reg_p1_n431) );
  NAND2_X1 reg_p1_U60 ( .A1(reg_p1_n429), .A2(reg_p1_n428), .ZN(reg_p1_n213)
         );
  NAND2_X1 reg_p1_U59 ( .A1(p1[52]), .A2(reg_p1_n432), .ZN(reg_p1_n428) );
  NAND2_X1 reg_p1_U58 ( .A1(init_y[20]), .A2(reg_p1_n451), .ZN(reg_p1_n429) );
  NAND2_X1 reg_p1_U57 ( .A1(reg_p1_n427), .A2(reg_p1_n426), .ZN(reg_p1_n214)
         );
  NAND2_X1 reg_p1_U56 ( .A1(p1[51]), .A2(reg_p1_n432), .ZN(reg_p1_n426) );
  NAND2_X1 reg_p1_U55 ( .A1(init_y[3]), .A2(reg_p1_n451), .ZN(reg_p1_n427) );
  NAND2_X1 reg_p1_U54 ( .A1(reg_p1_n425), .A2(reg_p1_n424), .ZN(reg_p1_n215)
         );
  NAND2_X1 reg_p1_U53 ( .A1(p1[50]), .A2(reg_p1_n432), .ZN(reg_p1_n424) );
  NAND2_X1 reg_p1_U52 ( .A1(init_y[2]), .A2(reg_p1_n451), .ZN(reg_p1_n425) );
  NAND2_X1 reg_p1_U51 ( .A1(reg_p1_n423), .A2(reg_p1_n422), .ZN(reg_p1_n216)
         );
  NAND2_X1 reg_p1_U50 ( .A1(p1[49]), .A2(reg_p1_n432), .ZN(reg_p1_n422) );
  NAND2_X1 reg_p1_U49 ( .A1(init_y[1]), .A2(reg_p1_n421), .ZN(reg_p1_n423) );
  NAND2_X1 reg_p1_U48 ( .A1(reg_p1_n420), .A2(reg_p1_n419), .ZN(reg_p1_n217)
         );
  NAND2_X1 reg_p1_U47 ( .A1(p1[48]), .A2(reg_p1_n432), .ZN(reg_p1_n419) );
  NAND2_X1 reg_p1_U46 ( .A1(init_y[0]), .A2(reg_p1_n421), .ZN(reg_p1_n420) );
  NAND2_X1 reg_p1_U45 ( .A1(reg_p1_n418), .A2(reg_p1_n417), .ZN(reg_p1_n218)
         );
  NAND2_X1 reg_p1_U44 ( .A1(p1[47]), .A2(reg_p1_n432), .ZN(reg_p1_n417) );
  NAND2_X1 reg_p1_U43 ( .A1(init_y[47]), .A2(reg_p1_n421), .ZN(reg_p1_n418) );
  NAND2_X1 reg_p1_U42 ( .A1(reg_p1_n416), .A2(reg_p1_n415), .ZN(reg_p1_n219)
         );
  NAND2_X1 reg_p1_U41 ( .A1(p1[46]), .A2(reg_p1_n432), .ZN(reg_p1_n415) );
  NAND2_X1 reg_p1_U40 ( .A1(init_y[46]), .A2(reg_p1_n421), .ZN(reg_p1_n416) );
  NAND2_X1 reg_p1_U39 ( .A1(reg_p1_n414), .A2(reg_p1_n413), .ZN(reg_p1_n220)
         );
  NAND2_X1 reg_p1_U38 ( .A1(p1[45]), .A2(reg_p1_n432), .ZN(reg_p1_n413) );
  NAND2_X1 reg_p1_U37 ( .A1(init_y[45]), .A2(reg_p1_n421), .ZN(reg_p1_n414) );
  NAND2_X1 reg_p1_U36 ( .A1(reg_p1_n412), .A2(reg_p1_n411), .ZN(reg_p1_n221)
         );
  NAND2_X1 reg_p1_U35 ( .A1(p1[44]), .A2(reg_p1_n432), .ZN(reg_p1_n411) );
  NAND2_X1 reg_p1_U34 ( .A1(init_y[44]), .A2(reg_p1_n421), .ZN(reg_p1_n412) );
  NAND2_X1 reg_p1_U33 ( .A1(reg_p1_n410), .A2(reg_p1_n409), .ZN(reg_p1_n222)
         );
  NAND2_X1 reg_p1_U32 ( .A1(p1[43]), .A2(reg_p1_n432), .ZN(reg_p1_n409) );
  NAND2_X1 reg_p1_U31 ( .A1(init_y[27]), .A2(reg_p1_n421), .ZN(reg_p1_n410) );
  NAND2_X1 reg_p1_U30 ( .A1(reg_p1_n408), .A2(reg_p1_n407), .ZN(reg_p1_n223)
         );
  NAND2_X1 reg_p1_U29 ( .A1(p1[42]), .A2(reg_p1_n432), .ZN(reg_p1_n407) );
  NAND2_X1 reg_p1_U28 ( .A1(init_y[26]), .A2(reg_p1_n421), .ZN(reg_p1_n408) );
  NAND2_X1 reg_p1_U27 ( .A1(reg_p1_n406), .A2(reg_p1_n405), .ZN(reg_p1_n224)
         );
  NAND2_X1 reg_p1_U26 ( .A1(p1[41]), .A2(reg_p1_n432), .ZN(reg_p1_n405) );
  NAND2_X1 reg_p1_U25 ( .A1(init_y[25]), .A2(reg_p1_n421), .ZN(reg_p1_n406) );
  NAND2_X1 reg_p1_U24 ( .A1(reg_p1_n404), .A2(reg_p1_n403), .ZN(reg_p1_n225)
         );
  NAND2_X1 reg_p1_U23 ( .A1(p1[40]), .A2(reg_p1_n432), .ZN(reg_p1_n403) );
  NAND2_X1 reg_p1_U22 ( .A1(init_y[24]), .A2(reg_p1_n451), .ZN(reg_p1_n404) );
  NAND2_X1 reg_p1_U21 ( .A1(reg_p1_n402), .A2(reg_p1_n401), .ZN(reg_p1_n226)
         );
  NAND2_X1 reg_p1_U20 ( .A1(p1[39]), .A2(reg_p1_n432), .ZN(reg_p1_n401) );
  NAND2_X1 reg_p1_U19 ( .A1(init_y[7]), .A2(reg_p1_n451), .ZN(reg_p1_n402) );
  NAND2_X1 reg_p1_U18 ( .A1(reg_p1_n400), .A2(reg_p1_n399), .ZN(reg_p1_n227)
         );
  NAND2_X1 reg_p1_U17 ( .A1(p1[38]), .A2(reg_p1_n432), .ZN(reg_p1_n399) );
  NAND2_X1 reg_p1_U16 ( .A1(init_y[6]), .A2(reg_p1_n451), .ZN(reg_p1_n400) );
  NAND2_X1 reg_p1_U15 ( .A1(reg_p1_n398), .A2(reg_p1_n397), .ZN(reg_p1_n228)
         );
  NAND2_X1 reg_p1_U14 ( .A1(p1[37]), .A2(reg_p1_n432), .ZN(reg_p1_n397) );
  NAND2_X1 reg_p1_U13 ( .A1(init_y[5]), .A2(reg_p1_n451), .ZN(reg_p1_n398) );
  NAND2_X1 reg_p1_U12 ( .A1(reg_p1_n396), .A2(reg_p1_n395), .ZN(reg_p1_n229)
         );
  NAND2_X1 reg_p1_U11 ( .A1(reg_p1_n451), .A2(init_y[4]), .ZN(reg_p1_n395) );
  INV_X1 reg_p1_U10 ( .A(reg_p1_n457), .ZN(reg_p1_n451) );
  INV_X1 reg_p1_U9 ( .A(reg_p1_n421), .ZN(reg_p1_n457) );
  NAND2_X1 reg_p1_U8 ( .A1(reg_p1_n432), .A2(p1[36]), .ZN(reg_p1_n396) );
  INV_X1 reg_p1_U7 ( .A(reg_p1_n458), .ZN(reg_p1_n432) );
  INV_X1 reg_p1_U6 ( .A(reg_p1_n452), .ZN(reg_p1_n458) );
  NOR2_X1 reg_p1_U5 ( .A1(rst), .A2(reg_p1_n394), .ZN(reg_p1_n452) );
  NOR2_X1 reg_p1_U4 ( .A1(rst), .A2(en_sig), .ZN(reg_p1_n421) );
  INV_X1 reg_p1_U3 ( .A(en_sig), .ZN(reg_p1_n394) );
  DFF_X1 reg_p1_s_current_state_reg_0_ ( .D(reg_p1_n265), .CK(clk), .Q(
        init_y[16]) );
  DFF_X1 reg_p1_s_current_state_reg_1_ ( .D(reg_p1_n264), .CK(clk), .Q(
        init_y[17]) );
  DFF_X1 reg_p1_s_current_state_reg_2_ ( .D(reg_p1_n263), .CK(clk), .Q(
        init_y[18]) );
  DFF_X1 reg_p1_s_current_state_reg_3_ ( .D(reg_p1_n262), .CK(clk), .Q(
        init_y[19]) );
  DFF_X1 reg_p1_s_current_state_reg_4_ ( .D(reg_p1_n261), .CK(clk), .Q(
        init_y[36]) );
  DFF_X1 reg_p1_s_current_state_reg_5_ ( .D(reg_p1_n260), .CK(clk), .Q(
        init_y[37]) );
  DFF_X1 reg_p1_s_current_state_reg_6_ ( .D(reg_p1_n259), .CK(clk), .Q(
        init_y[38]) );
  DFF_X1 reg_p1_s_current_state_reg_7_ ( .D(reg_p1_n258), .CK(clk), .Q(
        init_y[39]) );
  DFF_X1 reg_p1_s_current_state_reg_8_ ( .D(reg_p1_n257), .CK(clk), .Q(
        init_y[56]) );
  DFF_X1 reg_p1_s_current_state_reg_9_ ( .D(reg_p1_n256), .CK(clk), .Q(
        init_y[57]) );
  DFF_X1 reg_p1_s_current_state_reg_10_ ( .D(reg_p1_n255), .CK(clk), .Q(
        init_y[58]) );
  DFF_X1 reg_p1_s_current_state_reg_11_ ( .D(reg_p1_n254), .CK(clk), .Q(
        init_y[59]) );
  DFF_X1 reg_p1_s_current_state_reg_12_ ( .D(reg_p1_n253), .CK(clk), .Q(
        init_y[12]) );
  DFF_X1 reg_p1_s_current_state_reg_13_ ( .D(reg_p1_n252), .CK(clk), .Q(
        init_y[13]) );
  DFF_X1 reg_p1_s_current_state_reg_14_ ( .D(reg_p1_n251), .CK(clk), .Q(
        init_y[14]) );
  DFF_X1 reg_p1_s_current_state_reg_15_ ( .D(reg_p1_n250), .CK(clk), .Q(
        init_y[15]) );
  DFF_X1 reg_p1_s_current_state_reg_16_ ( .D(reg_p1_n249), .CK(clk), .Q(
        init_y[32]) );
  DFF_X1 reg_p1_s_current_state_reg_17_ ( .D(reg_p1_n248), .CK(clk), .Q(
        init_y[33]) );
  DFF_X1 reg_p1_s_current_state_reg_18_ ( .D(reg_p1_n247), .CK(clk), .Q(
        init_y[34]) );
  DFF_X1 reg_p1_s_current_state_reg_19_ ( .D(reg_p1_n246), .CK(clk), .Q(
        init_y[35]) );
  DFF_X1 reg_p1_s_current_state_reg_20_ ( .D(reg_p1_n245), .CK(clk), .Q(
        init_y[52]) );
  DFF_X1 reg_p1_s_current_state_reg_21_ ( .D(reg_p1_n244), .CK(clk), .Q(
        init_y[53]) );
  DFF_X1 reg_p1_s_current_state_reg_22_ ( .D(reg_p1_n243), .CK(clk), .Q(
        init_y[54]) );
  DFF_X1 reg_p1_s_current_state_reg_23_ ( .D(reg_p1_n242), .CK(clk), .Q(
        init_y[55]) );
  DFF_X1 reg_p1_s_current_state_reg_24_ ( .D(reg_p1_n241), .CK(clk), .Q(
        init_y[8]) );
  DFF_X1 reg_p1_s_current_state_reg_25_ ( .D(reg_p1_n240), .CK(clk), .Q(
        init_y[9]) );
  DFF_X1 reg_p1_s_current_state_reg_26_ ( .D(reg_p1_n239), .CK(clk), .Q(
        init_y[10]) );
  DFF_X1 reg_p1_s_current_state_reg_27_ ( .D(reg_p1_n238), .CK(clk), .Q(
        init_y[11]) );
  DFF_X1 reg_p1_s_current_state_reg_28_ ( .D(reg_p1_n237), .CK(clk), .Q(
        init_y[28]) );
  DFF_X1 reg_p1_s_current_state_reg_29_ ( .D(reg_p1_n236), .CK(clk), .Q(
        init_y[29]) );
  DFF_X1 reg_p1_s_current_state_reg_30_ ( .D(reg_p1_n235), .CK(clk), .Q(
        init_y[30]) );
  DFF_X1 reg_p1_s_current_state_reg_31_ ( .D(reg_p1_n234), .CK(clk), .Q(
        init_y[31]) );
  DFF_X1 reg_p1_s_current_state_reg_32_ ( .D(reg_p1_n233), .CK(clk), .Q(
        init_y[48]) );
  DFF_X1 reg_p1_s_current_state_reg_33_ ( .D(reg_p1_n232), .CK(clk), .Q(
        init_y[49]) );
  DFF_X1 reg_p1_s_current_state_reg_34_ ( .D(reg_p1_n231), .CK(clk), .Q(
        init_y[50]) );
  DFF_X1 reg_p1_s_current_state_reg_35_ ( .D(reg_p1_n230), .CK(clk), .Q(
        init_y[51]) );
  DFF_X1 reg_p1_s_current_state_reg_36_ ( .D(reg_p1_n229), .CK(clk), .Q(
        init_y[4]) );
  DFF_X1 reg_p1_s_current_state_reg_37_ ( .D(reg_p1_n228), .CK(clk), .Q(
        init_y[5]) );
  DFF_X1 reg_p1_s_current_state_reg_38_ ( .D(reg_p1_n227), .CK(clk), .Q(
        init_y[6]) );
  DFF_X1 reg_p1_s_current_state_reg_39_ ( .D(reg_p1_n226), .CK(clk), .Q(
        init_y[7]) );
  DFF_X1 reg_p1_s_current_state_reg_40_ ( .D(reg_p1_n225), .CK(clk), .Q(
        init_y[24]) );
  DFF_X1 reg_p1_s_current_state_reg_41_ ( .D(reg_p1_n224), .CK(clk), .Q(
        init_y[25]) );
  DFF_X1 reg_p1_s_current_state_reg_42_ ( .D(reg_p1_n223), .CK(clk), .Q(
        init_y[26]) );
  DFF_X1 reg_p1_s_current_state_reg_43_ ( .D(reg_p1_n222), .CK(clk), .Q(
        init_y[27]) );
  DFF_X1 reg_p1_s_current_state_reg_44_ ( .D(reg_p1_n221), .CK(clk), .Q(
        init_y[44]) );
  DFF_X1 reg_p1_s_current_state_reg_45_ ( .D(reg_p1_n220), .CK(clk), .Q(
        init_y[45]) );
  DFF_X1 reg_p1_s_current_state_reg_46_ ( .D(reg_p1_n219), .CK(clk), .Q(
        init_y[46]) );
  DFF_X1 reg_p1_s_current_state_reg_47_ ( .D(reg_p1_n218), .CK(clk), .Q(
        init_y[47]) );
  DFF_X1 reg_p1_s_current_state_reg_48_ ( .D(reg_p1_n217), .CK(clk), .Q(
        init_y[0]) );
  DFF_X1 reg_p1_s_current_state_reg_49_ ( .D(reg_p1_n216), .CK(clk), .Q(
        init_y[1]) );
  DFF_X1 reg_p1_s_current_state_reg_50_ ( .D(reg_p1_n215), .CK(clk), .Q(
        init_y[2]) );
  DFF_X1 reg_p1_s_current_state_reg_51_ ( .D(reg_p1_n214), .CK(clk), .Q(
        init_y[3]) );
  DFF_X1 reg_p1_s_current_state_reg_52_ ( .D(reg_p1_n213), .CK(clk), .Q(
        init_y[20]) );
  DFF_X1 reg_p1_s_current_state_reg_53_ ( .D(reg_p1_n212), .CK(clk), .Q(
        init_y[21]) );
  DFF_X1 reg_p1_s_current_state_reg_54_ ( .D(reg_p1_n211), .CK(clk), .Q(
        init_y[22]) );
  DFF_X1 reg_p1_s_current_state_reg_55_ ( .D(reg_p1_n210), .CK(clk), .Q(
        init_y[23]) );
  DFF_X1 reg_p1_s_current_state_reg_56_ ( .D(reg_p1_n209), .CK(clk), .Q(
        init_y[40]) );
  DFF_X1 reg_p1_s_current_state_reg_57_ ( .D(reg_p1_n208), .CK(clk), .Q(
        init_y[41]) );
  DFF_X1 reg_p1_s_current_state_reg_58_ ( .D(reg_p1_n207), .CK(clk), .Q(
        init_y[42]) );
  DFF_X1 reg_p1_s_current_state_reg_59_ ( .D(reg_p1_n206), .CK(clk), .Q(
        init_y[43]) );
  DFF_X1 reg_p1_s_current_state_reg_60_ ( .D(reg_p1_n205), .CK(clk), .Q(
        init_y[60]) );
  DFF_X1 reg_p1_s_current_state_reg_61_ ( .D(reg_p1_n204), .CK(clk), .Q(
        init_y[61]) );
  DFF_X1 reg_p1_s_current_state_reg_62_ ( .D(reg_p1_n203), .CK(clk), .Q(
        init_y[62]) );
  DFF_X1 reg_p1_s_current_state_reg_63_ ( .D(reg_p1_n202), .CK(clk), .Q(
        init_y[63]) );
  MUX2_X1 mux_x_U68 ( .A(rout_x[9]), .B(init_x[9]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[57]) );
  MUX2_X1 mux_x_U67 ( .A(rout_x[6]), .B(init_x[6]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[38]) );
  MUX2_X1 mux_x_U66 ( .A(rout_x[7]), .B(init_x[7]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[39]) );
  MUX2_X1 mux_x_U65 ( .A(rout_x[8]), .B(init_x[8]), .S(start_sig), .Z(
        prince_inst_srin_x[56]) );
  MUX2_X1 mux_x_U64 ( .A(rout_x[62]), .B(init_x[62]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[62]) );
  MUX2_X1 mux_x_U63 ( .A(rout_x[61]), .B(init_x[61]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[61]) );
  MUX2_X1 mux_x_U62 ( .A(rout_x[63]), .B(init_x[63]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[63]) );
  MUX2_X1 mux_x_U61 ( .A(rout_x[10]), .B(init_x[10]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[58]) );
  MUX2_X1 mux_x_U60 ( .A(rout_x[11]), .B(init_x[11]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[59]) );
  MUX2_X1 mux_x_U59 ( .A(rout_x[22]), .B(init_x[22]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[54]) );
  MUX2_X1 mux_x_U58 ( .A(rout_x[21]), .B(init_x[21]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[53]) );
  MUX2_X1 mux_x_U57 ( .A(rout_x[23]), .B(init_x[23]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[55]) );
  MUX2_X1 mux_x_U56 ( .A(rout_x[34]), .B(init_x[34]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[50]) );
  MUX2_X1 mux_x_U55 ( .A(rout_x[33]), .B(init_x[33]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[49]) );
  MUX2_X1 mux_x_U54 ( .A(rout_x[35]), .B(init_x[35]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[51]) );
  MUX2_X1 mux_x_U53 ( .A(rout_x[46]), .B(init_x[46]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[46]) );
  MUX2_X1 mux_x_U52 ( .A(rout_x[45]), .B(init_x[45]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[45]) );
  MUX2_X1 mux_x_U51 ( .A(rout_x[47]), .B(init_x[47]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[47]) );
  MUX2_X1 mux_x_U50 ( .A(rout_x[58]), .B(init_x[58]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[42]) );
  MUX2_X1 mux_x_U49 ( .A(rout_x[57]), .B(init_x[57]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[41]) );
  MUX2_X1 mux_x_U48 ( .A(rout_x[59]), .B(init_x[59]), .S(start_sig), .Z(
        prince_inst_srin_x[43]) );
  MUX2_X1 mux_x_U47 ( .A(rout_x[5]), .B(init_x[5]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[37]) );
  MUX2_X1 mux_x_U46 ( .A(rout_x[18]), .B(init_x[18]), .S(start_sig), .Z(
        prince_inst_srin_x[34]) );
  MUX2_X1 mux_x_U45 ( .A(rout_x[17]), .B(init_x[17]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[33]) );
  MUX2_X1 mux_x_U44 ( .A(rout_x[19]), .B(init_x[19]), .S(start_sig), .Z(
        prince_inst_srin_x[35]) );
  MUX2_X1 mux_x_U43 ( .A(rout_x[30]), .B(init_x[30]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[30]) );
  MUX2_X1 mux_x_U42 ( .A(rout_x[29]), .B(init_x[29]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[29]) );
  MUX2_X1 mux_x_U41 ( .A(rout_x[31]), .B(init_x[31]), .S(start_sig), .Z(
        prince_inst_srin_x[31]) );
  MUX2_X1 mux_x_U40 ( .A(rout_x[42]), .B(init_x[42]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[26]) );
  MUX2_X1 mux_x_U39 ( .A(rout_x[41]), .B(init_x[41]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[25]) );
  MUX2_X1 mux_x_U38 ( .A(rout_x[43]), .B(init_x[43]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[27]) );
  MUX2_X1 mux_x_U37 ( .A(rout_x[54]), .B(init_x[54]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[22]) );
  MUX2_X1 mux_x_U36 ( .A(rout_x[53]), .B(init_x[53]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[21]) );
  MUX2_X1 mux_x_U35 ( .A(rout_x[55]), .B(init_x[55]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[23]) );
  MUX2_X1 mux_x_U34 ( .A(rout_x[2]), .B(init_x[2]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[18]) );
  MUX2_X1 mux_x_U33 ( .A(rout_x[1]), .B(init_x[1]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[17]) );
  MUX2_X1 mux_x_U32 ( .A(rout_x[3]), .B(init_x[3]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[19]) );
  MUX2_X1 mux_x_U31 ( .A(rout_x[14]), .B(init_x[14]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[14]) );
  MUX2_X1 mux_x_U30 ( .A(rout_x[13]), .B(init_x[13]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[13]) );
  MUX2_X1 mux_x_U29 ( .A(rout_x[15]), .B(init_x[15]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[15]) );
  MUX2_X1 mux_x_U28 ( .A(rout_x[26]), .B(init_x[26]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[10]) );
  MUX2_X1 mux_x_U27 ( .A(rout_x[25]), .B(init_x[25]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[9]) );
  MUX2_X1 mux_x_U26 ( .A(rout_x[27]), .B(init_x[27]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[11]) );
  MUX2_X1 mux_x_U25 ( .A(rout_x[38]), .B(init_x[38]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[6]) );
  MUX2_X1 mux_x_U24 ( .A(rout_x[37]), .B(init_x[37]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[5]) );
  MUX2_X1 mux_x_U23 ( .A(rout_x[39]), .B(init_x[39]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[7]) );
  MUX2_X1 mux_x_U22 ( .A(rout_x[50]), .B(init_x[50]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[2]) );
  MUX2_X1 mux_x_U21 ( .A(rout_x[51]), .B(init_x[51]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[3]) );
  MUX2_X1 mux_x_U20 ( .A(rout_x[49]), .B(init_x[49]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[1]) );
  MUX2_X1 mux_x_U19 ( .A(rout_x[60]), .B(init_x[60]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[60]) );
  MUX2_X1 mux_x_U18 ( .A(rout_x[20]), .B(init_x[20]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[52]) );
  MUX2_X1 mux_x_U17 ( .A(rout_x[32]), .B(init_x[32]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[48]) );
  MUX2_X1 mux_x_U16 ( .A(rout_x[44]), .B(init_x[44]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[44]) );
  MUX2_X1 mux_x_U15 ( .A(rout_x[56]), .B(init_x[56]), .S(start_sig), .Z(
        prince_inst_srin_x[40]) );
  MUX2_X1 mux_x_U14 ( .A(rout_x[4]), .B(init_x[4]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[36]) );
  MUX2_X1 mux_x_U13 ( .A(rout_x[16]), .B(init_x[16]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[32]) );
  MUX2_X1 mux_x_U12 ( .A(rout_x[28]), .B(init_x[28]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[28]) );
  MUX2_X1 mux_x_U11 ( .A(rout_x[40]), .B(init_x[40]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[24]) );
  MUX2_X1 mux_x_U10 ( .A(rout_x[52]), .B(init_x[52]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[20]) );
  MUX2_X1 mux_x_U9 ( .A(rout_x[0]), .B(init_x[0]), .S(start_sig), .Z(
        prince_inst_srin_x[16]) );
  MUX2_X1 mux_x_U8 ( .A(rout_x[12]), .B(init_x[12]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[12]) );
  MUX2_X1 mux_x_U7 ( .A(rout_x[24]), .B(init_x[24]), .S(mux_x_n136), .Z(
        prince_inst_srin_x[8]) );
  INV_X1 mux_x_U6 ( .A(mux_x_n135), .ZN(mux_x_n136) );
  MUX2_X1 mux_x_U5 ( .A(rout_x[36]), .B(init_x[36]), .S(mux_x_n137), .Z(
        prince_inst_srin_x[4]) );
  INV_X1 mux_x_U4 ( .A(mux_x_n135), .ZN(mux_x_n137) );
  MUX2_X1 mux_x_U3 ( .A(rout_x[48]), .B(init_x[48]), .S(mux_x_n138), .Z(
        prince_inst_srin_x[0]) );
  INV_X1 mux_x_U2 ( .A(mux_x_n135), .ZN(mux_x_n138) );
  INV_X1 mux_x_U1 ( .A(start_sig), .ZN(mux_x_n135) );
  MUX2_X1 mux_y_U69 ( .A(rout_y[9]), .B(init_y[9]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[57]) );
  MUX2_X1 mux_y_U68 ( .A(rout_y[6]), .B(init_y[6]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[38]) );
  MUX2_X1 mux_y_U67 ( .A(rout_y[7]), .B(init_y[7]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[39]) );
  MUX2_X1 mux_y_U66 ( .A(rout_y[51]), .B(init_y[51]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[3]) );
  MUX2_X1 mux_y_U65 ( .A(rout_y[19]), .B(init_y[19]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[35]) );
  MUX2_X1 mux_y_U64 ( .A(rout_y[61]), .B(init_y[61]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[61]) );
  MUX2_X1 mux_y_U63 ( .A(rout_y[41]), .B(init_y[41]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[25]) );
  MUX2_X1 mux_y_U62 ( .A(rout_y[21]), .B(init_y[21]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[53]) );
  MUX2_X1 mux_y_U61 ( .A(rout_y[33]), .B(init_y[33]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[49]) );
  MUX2_X1 mux_y_U60 ( .A(rout_y[1]), .B(init_y[1]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[17]) );
  MUX2_X1 mux_y_U59 ( .A(rout_y[45]), .B(init_y[45]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[45]) );
  MUX2_X1 mux_y_U58 ( .A(rout_y[57]), .B(init_y[57]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[41]) );
  MUX2_X1 mux_y_U57 ( .A(rout_y[25]), .B(init_y[25]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[9]) );
  MUX2_X1 mux_y_U56 ( .A(rout_y[5]), .B(init_y[5]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[37]) );
  MUX2_X1 mux_y_U55 ( .A(rout_y[17]), .B(init_y[17]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[33]) );
  MUX2_X1 mux_y_U54 ( .A(rout_y[49]), .B(init_y[49]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[1]) );
  MUX2_X1 mux_y_U53 ( .A(rout_y[29]), .B(init_y[29]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[29]) );
  MUX2_X1 mux_y_U52 ( .A(rout_y[53]), .B(init_y[53]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[21]) );
  MUX2_X1 mux_y_U51 ( .A(rout_y[13]), .B(init_y[13]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[13]) );
  MUX2_X1 mux_y_U50 ( .A(rout_y[37]), .B(init_y[37]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[5]) );
  MUX2_X1 mux_y_U49 ( .A(rout_y[62]), .B(init_y[62]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[62]) );
  MUX2_X1 mux_y_U48 ( .A(rout_y[10]), .B(init_y[10]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[58]) );
  MUX2_X1 mux_y_U47 ( .A(rout_y[42]), .B(init_y[42]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[26]) );
  MUX2_X1 mux_y_U46 ( .A(rout_y[22]), .B(init_y[22]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[54]) );
  MUX2_X1 mux_y_U45 ( .A(rout_y[34]), .B(init_y[34]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[50]) );
  MUX2_X1 mux_y_U44 ( .A(rout_y[2]), .B(init_y[2]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[18]) );
  MUX2_X1 mux_y_U43 ( .A(rout_y[46]), .B(init_y[46]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[46]) );
  MUX2_X1 mux_y_U42 ( .A(rout_y[58]), .B(init_y[58]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[42]) );
  MUX2_X1 mux_y_U41 ( .A(rout_y[26]), .B(init_y[26]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[10]) );
  MUX2_X1 mux_y_U40 ( .A(rout_y[18]), .B(init_y[18]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[34]) );
  MUX2_X1 mux_y_U39 ( .A(rout_y[50]), .B(init_y[50]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[2]) );
  MUX2_X1 mux_y_U38 ( .A(rout_y[30]), .B(init_y[30]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[30]) );
  MUX2_X1 mux_y_U37 ( .A(rout_y[54]), .B(init_y[54]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[22]) );
  MUX2_X1 mux_y_U36 ( .A(rout_y[14]), .B(init_y[14]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[14]) );
  MUX2_X1 mux_y_U35 ( .A(rout_y[38]), .B(init_y[38]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[6]) );
  MUX2_X1 mux_y_U34 ( .A(rout_y[63]), .B(init_y[63]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[63]) );
  MUX2_X1 mux_y_U33 ( .A(rout_y[11]), .B(init_y[11]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[59]) );
  MUX2_X1 mux_y_U32 ( .A(rout_y[43]), .B(init_y[43]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[27]) );
  MUX2_X1 mux_y_U31 ( .A(rout_y[23]), .B(init_y[23]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[55]) );
  MUX2_X1 mux_y_U30 ( .A(rout_y[35]), .B(init_y[35]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[51]) );
  MUX2_X1 mux_y_U29 ( .A(rout_y[3]), .B(init_y[3]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[19]) );
  MUX2_X1 mux_y_U28 ( .A(rout_y[47]), .B(init_y[47]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[47]) );
  MUX2_X1 mux_y_U27 ( .A(rout_y[59]), .B(init_y[59]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[43]) );
  MUX2_X1 mux_y_U26 ( .A(rout_y[27]), .B(init_y[27]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[11]) );
  MUX2_X1 mux_y_U25 ( .A(rout_y[31]), .B(init_y[31]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[31]) );
  MUX2_X1 mux_y_U24 ( .A(rout_y[55]), .B(init_y[55]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[23]) );
  MUX2_X1 mux_y_U23 ( .A(rout_y[15]), .B(init_y[15]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[15]) );
  MUX2_X1 mux_y_U22 ( .A(rout_y[39]), .B(init_y[39]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[7]) );
  MUX2_X1 mux_y_U21 ( .A(rout_y[8]), .B(init_y[8]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[56]) );
  MUX2_X1 mux_y_U20 ( .A(rout_y[60]), .B(init_y[60]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[60]) );
  MUX2_X1 mux_y_U19 ( .A(rout_y[40]), .B(init_y[40]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[24]) );
  MUX2_X1 mux_y_U18 ( .A(rout_y[20]), .B(init_y[20]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[52]) );
  MUX2_X1 mux_y_U17 ( .A(rout_y[32]), .B(init_y[32]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[48]) );
  MUX2_X1 mux_y_U16 ( .A(rout_y[0]), .B(init_y[0]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[16]) );
  MUX2_X1 mux_y_U15 ( .A(rout_y[44]), .B(init_y[44]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[44]) );
  MUX2_X1 mux_y_U14 ( .A(rout_y[56]), .B(init_y[56]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[40]) );
  MUX2_X1 mux_y_U13 ( .A(rout_y[24]), .B(init_y[24]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[8]) );
  MUX2_X1 mux_y_U12 ( .A(rout_y[4]), .B(init_y[4]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[36]) );
  MUX2_X1 mux_y_U11 ( .A(rout_y[16]), .B(init_y[16]), .S(mux_y_n267), .Z(
        prince_inst_srin_y[32]) );
  INV_X1 mux_y_U10 ( .A(mux_y_n263), .ZN(mux_y_n267) );
  MUX2_X1 mux_y_U9 ( .A(rout_y[48]), .B(init_y[48]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[0]) );
  MUX2_X1 mux_y_U8 ( .A(rout_y[28]), .B(init_y[28]), .S(mux_y_n264), .Z(
        prince_inst_srin_y[28]) );
  INV_X1 mux_y_U7 ( .A(mux_y_n263), .ZN(mux_y_n264) );
  MUX2_X1 mux_y_U6 ( .A(rout_y[52]), .B(init_y[52]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[20]) );
  MUX2_X1 mux_y_U5 ( .A(rout_y[12]), .B(init_y[12]), .S(mux_y_n265), .Z(
        prince_inst_srin_y[12]) );
  INV_X1 mux_y_U4 ( .A(mux_y_n263), .ZN(mux_y_n265) );
  MUX2_X1 mux_y_U3 ( .A(rout_y[36]), .B(init_y[36]), .S(mux_y_n266), .Z(
        prince_inst_srin_y[4]) );
  INV_X1 mux_y_U2 ( .A(mux_y_n263), .ZN(mux_y_n266) );
  INV_X1 mux_y_U1 ( .A(start_sig), .ZN(mux_y_n263) );
  NOR3_X1 cntrl_inst_U296 ( .A1(cntrl_inst_n164), .A2(rst), .A3(
        cntrl_inst_n163), .ZN(cntrl_inst_n207) );
  NOR2_X1 cntrl_inst_U295 ( .A1(cntrl_inst_n168), .A2(cntrl_inst_counter_0_), 
        .ZN(cntrl_inst_n164) );
  MUX2_X1 cntrl_inst_U294 ( .A(cntrl_inst_n162), .B(cntrl_inst_n36), .S(
        cntrl_inst_n163), .Z(cntrl_inst_n208) );
  NOR2_X1 cntrl_inst_U293 ( .A1(cntrl_inst_n36), .A2(rst), .ZN(cntrl_inst_n162) );
  NAND2_X1 cntrl_inst_U292 ( .A1(cntrl_inst_n161), .A2(cntrl_inst_n160), .ZN(
        cntrl_inst_n209) );
  NAND2_X1 cntrl_inst_U291 ( .A1(cntrl_inst_n165), .A2(cntrl_inst_n3), .ZN(
        cntrl_inst_n160) );
  NAND2_X1 cntrl_inst_U290 ( .A1(cntrl_inst_n163), .A2(cntrl_inst_n166), .ZN(
        cntrl_inst_n161) );
  NOR2_X1 cntrl_inst_U289 ( .A1(cntrl_inst_n40), .A2(cntrl_inst_n159), .ZN(
        cntrl_inst_n163) );
  NAND2_X1 cntrl_inst_U288 ( .A1(cntrl_inst_n3), .A2(cntrl_inst_n158), .ZN(
        cntrl_inst_n210) );
  NAND2_X1 cntrl_inst_U287 ( .A1(cntrl_inst_n159), .A2(en_sig), .ZN(
        cntrl_inst_n158) );
  NAND3_X1 cntrl_inst_U286 ( .A1(cntrl_inst_counter_0_), .A2(cntrl_inst_n157), 
        .A3(cntrl_inst_n3), .ZN(cntrl_inst_n159) );
  NAND2_X1 cntrl_inst_U285 ( .A1(cntrl_inst_n156), .A2(cntrl_inst_n165), .ZN(
        inv_sig2) );
  NAND3_X1 cntrl_inst_U284 ( .A1(cntrl_inst_n167), .A2(cntrl_inst_n40), .A3(
        cntrl_inst_n36), .ZN(cntrl_inst_n156) );
  XOR2_X1 cntrl_inst_U283 ( .A(cntrl_inst_n155), .B(kext[176]), .Z(
        prince_inst_rc2_inv[0]) );
  XNOR2_X1 cntrl_inst_U282 ( .A(kext[179]), .B(cntrl_inst_n154), .ZN(
        prince_inst_rc2_inv[3]) );
  NOR3_X1 cntrl_inst_U281 ( .A1(cntrl_inst_n153), .A2(cntrl_inst_n152), .A3(
        cntrl_inst_n151), .ZN(cntrl_inst_n154) );
  XNOR2_X1 cntrl_inst_U280 ( .A(kext[171]), .B(cntrl_inst_n150), .ZN(
        prince_inst_rc2_inv[27]) );
  NOR3_X1 cntrl_inst_U279 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n148), .A3(
        cntrl_inst_n147), .ZN(cntrl_inst_n150) );
  XNOR2_X1 cntrl_inst_U278 ( .A(cntrl_inst_n146), .B(kext[152]), .ZN(
        prince_inst_rc2_inv[8]) );
  NOR2_X1 cntrl_inst_U277 ( .A1(cntrl_inst_n147), .A2(cntrl_inst_n145), .ZN(
        cntrl_inst_n146) );
  INV_X1 cntrl_inst_U276 ( .A(cntrl_inst_n144), .ZN(cntrl_inst_n145) );
  XNOR2_X1 cntrl_inst_U275 ( .A(cntrl_inst_n143), .B(kext[146]), .ZN(
        prince_inst_rc2_inv[34]) );
  XNOR2_X1 cntrl_inst_U274 ( .A(cntrl_inst_n143), .B(kext[135]), .ZN(
        prince_inst_rc2_inv[39]) );
  NOR3_X1 cntrl_inst_U273 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n142), .A3(
        cntrl_inst_n141), .ZN(cntrl_inst_n143) );
  XNOR2_X1 cntrl_inst_U272 ( .A(kext[178]), .B(cntrl_inst_n140), .ZN(
        prince_inst_rc2_inv[2]) );
  XNOR2_X1 cntrl_inst_U271 ( .A(kext[131]), .B(cntrl_inst_n140), .ZN(
        prince_inst_rc2_inv[19]) );
  NOR2_X1 cntrl_inst_U270 ( .A1(cntrl_inst_n139), .A2(cntrl_inst_n138), .ZN(
        cntrl_inst_n140) );
  INV_X1 cntrl_inst_U269 ( .A(cntrl_inst_n137), .ZN(cntrl_inst_n139) );
  XOR2_X1 cntrl_inst_U268 ( .A(kext[155]), .B(cntrl_inst_n136), .Z(
        prince_inst_rc2_inv[11]) );
  NAND2_X1 cntrl_inst_U267 ( .A1(cntrl_inst_n135), .A2(cntrl_inst_n134), .ZN(
        cntrl_inst_n136) );
  XNOR2_X1 cntrl_inst_U266 ( .A(cntrl_inst_n133), .B(kext[173]), .ZN(
        prince_inst_rc2_inv[45]) );
  NOR2_X1 cntrl_inst_U265 ( .A1(cntrl_inst_n138), .A2(cntrl_inst_n132), .ZN(
        cntrl_inst_n133) );
  XNOR2_X1 cntrl_inst_U264 ( .A(kext[167]), .B(cntrl_inst_n131), .ZN(
        prince_inst_rc2_inv[7]) );
  NOR2_X1 cntrl_inst_U263 ( .A1(cntrl_inst_n130), .A2(cntrl_inst_n138), .ZN(
        cntrl_inst_n131) );
  INV_X1 cntrl_inst_U262 ( .A(cntrl_inst_n129), .ZN(cntrl_inst_n130) );
  XNOR2_X1 cntrl_inst_U261 ( .A(kext[147]), .B(cntrl_inst_n128), .ZN(
        prince_inst_rc2_inv[35]) );
  NOR3_X1 cntrl_inst_U260 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n142), .A3(
        cntrl_inst_n138), .ZN(cntrl_inst_n128) );
  NAND3_X1 cntrl_inst_U259 ( .A1(cntrl_inst_n127), .A2(cntrl_inst_n126), .A3(
        cntrl_inst_n125), .ZN(cntrl_inst_n138) );
  INV_X1 cntrl_inst_U258 ( .A(cntrl_inst_n124), .ZN(cntrl_inst_n126) );
  XOR2_X1 cntrl_inst_U257 ( .A(kext[183]), .B(cntrl_inst_n123), .Z(
        prince_inst_rc2_inv[23]) );
  NAND2_X1 cntrl_inst_U256 ( .A1(cntrl_inst_n122), .A2(cntrl_inst_n137), .ZN(
        cntrl_inst_n123) );
  XOR2_X1 cntrl_inst_U255 ( .A(kext[190]), .B(cntrl_inst_n121), .Z(rc[62]) );
  XOR2_X1 cntrl_inst_U254 ( .A(kext[189]), .B(cntrl_inst_n120), .Z(rc[61]) );
  XOR2_X1 cntrl_inst_U253 ( .A(kext[191]), .B(cntrl_inst_n119), .Z(rc[63]) );
  NAND3_X1 cntrl_inst_U252 ( .A1(cntrl_inst_n118), .A2(cntrl_inst_n117), .A3(
        cntrl_inst_n116), .ZN(cntrl_inst_n119) );
  NAND2_X1 cntrl_inst_U251 ( .A1(cntrl_inst_n115), .A2(cntrl_inst_n114), .ZN(
        cntrl_inst_n118) );
  XOR2_X1 cntrl_inst_U250 ( .A(kext[186]), .B(cntrl_inst_n113), .Z(rc[58]) );
  XOR2_X1 cntrl_inst_U249 ( .A(kext[185]), .B(cntrl_inst_n112), .Z(rc[57]) );
  XNOR2_X1 cntrl_inst_U248 ( .A(kext[181]), .B(cntrl_inst_n111), .ZN(rc[53])
         );
  XOR2_X1 cntrl_inst_U247 ( .A(kext[183]), .B(cntrl_inst_n110), .Z(rc[55]) );
  NOR2_X1 cntrl_inst_U246 ( .A1(cntrl_inst_n109), .A2(cntrl_inst_n108), .ZN(
        cntrl_inst_n110) );
  XNOR2_X1 cntrl_inst_U245 ( .A(cntrl_inst_n107), .B(kext[178]), .ZN(rc[50])
         );
  XNOR2_X1 cntrl_inst_U244 ( .A(cntrl_inst_n106), .B(kext[177]), .ZN(rc[49])
         );
  XNOR2_X1 cntrl_inst_U243 ( .A(cntrl_inst_n105), .B(kext[179]), .ZN(rc[51])
         );
  NOR2_X1 cntrl_inst_U242 ( .A1(cntrl_inst_n104), .A2(cntrl_inst_n103), .ZN(
        cntrl_inst_n105) );
  XNOR2_X1 cntrl_inst_U241 ( .A(kext[173]), .B(cntrl_inst_n102), .ZN(rc[45])
         );
  NOR2_X1 cntrl_inst_U240 ( .A1(cntrl_inst_n101), .A2(cntrl_inst_n100), .ZN(
        cntrl_inst_n102) );
  XOR2_X1 cntrl_inst_U239 ( .A(kext[175]), .B(cntrl_inst_n99), .Z(rc[47]) );
  NAND2_X1 cntrl_inst_U238 ( .A1(cntrl_inst_n98), .A2(cntrl_inst_n106), .ZN(
        cntrl_inst_n99) );
  NOR2_X1 cntrl_inst_U237 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n103), .ZN(
        cntrl_inst_n106) );
  XOR2_X1 cntrl_inst_U236 ( .A(kext[169]), .B(cntrl_inst_n97), .Z(rc[41]) );
  XNOR2_X1 cntrl_inst_U235 ( .A(cntrl_inst_n96), .B(kext[171]), .ZN(rc[43]) );
  NOR2_X1 cntrl_inst_U234 ( .A1(cntrl_inst_n95), .A2(cntrl_inst_n103), .ZN(
        cntrl_inst_n96) );
  XOR2_X1 cntrl_inst_U233 ( .A(kext[166]), .B(cntrl_inst_n94), .Z(rc[38]) );
  XNOR2_X1 cntrl_inst_U232 ( .A(cntrl_inst_n93), .B(kext[165]), .ZN(rc[37]) );
  XNOR2_X1 cntrl_inst_U231 ( .A(cntrl_inst_n92), .B(kext[167]), .ZN(rc[39]) );
  NOR2_X1 cntrl_inst_U230 ( .A1(cntrl_inst_n100), .A2(cntrl_inst_n91), .ZN(
        cntrl_inst_n92) );
  XOR2_X1 cntrl_inst_U229 ( .A(kext[163]), .B(cntrl_inst_n97), .Z(rc[35]) );
  NAND2_X1 cntrl_inst_U228 ( .A1(cntrl_inst_n98), .A2(cntrl_inst_n90), .ZN(
        cntrl_inst_n97) );
  XNOR2_X1 cntrl_inst_U227 ( .A(kext[158]), .B(cntrl_inst_n89), .ZN(rc[30]) );
  XNOR2_X1 cntrl_inst_U226 ( .A(kext[159]), .B(cntrl_inst_n89), .ZN(rc[31]) );
  XNOR2_X1 cntrl_inst_U225 ( .A(cntrl_inst_n88), .B(kext[155]), .ZN(rc[27]) );
  NOR2_X1 cntrl_inst_U224 ( .A1(cntrl_inst_n87), .A2(cntrl_inst_n101), .ZN(
        cntrl_inst_n88) );
  INV_X1 cntrl_inst_U223 ( .A(cntrl_inst_n86), .ZN(cntrl_inst_n101) );
  XOR2_X1 cntrl_inst_U222 ( .A(kext[151]), .B(cntrl_inst_n113), .Z(rc[23]) );
  NAND3_X1 cntrl_inst_U221 ( .A1(cntrl_inst_n85), .A2(cntrl_inst_n86), .A3(
        cntrl_inst_n84), .ZN(cntrl_inst_n113) );
  XNOR2_X1 cntrl_inst_U220 ( .A(kext[146]), .B(cntrl_inst_n83), .ZN(rc[18]) );
  XNOR2_X1 cntrl_inst_U219 ( .A(kext[147]), .B(cntrl_inst_n82), .ZN(rc[19]) );
  NOR3_X1 cntrl_inst_U218 ( .A1(cntrl_inst_n81), .A2(cntrl_inst_n151), .A3(
        cntrl_inst_n100), .ZN(cntrl_inst_n82) );
  INV_X1 cntrl_inst_U217 ( .A(cntrl_inst_n80), .ZN(cntrl_inst_n151) );
  XOR2_X1 cntrl_inst_U216 ( .A(kext[141]), .B(cntrl_inst_n79), .Z(rc[13]) );
  NAND3_X1 cntrl_inst_U215 ( .A1(cntrl_inst_n98), .A2(cntrl_inst_n144), .A3(
        cntrl_inst_n78), .ZN(cntrl_inst_n79) );
  XOR2_X1 cntrl_inst_U214 ( .A(kext[137]), .B(cntrl_inst_n77), .Z(rc[9]) );
  XOR2_X1 cntrl_inst_U213 ( .A(kext[133]), .B(cntrl_inst_n94), .Z(rc[5]) );
  XNOR2_X1 cntrl_inst_U212 ( .A(kext[135]), .B(cntrl_inst_n83), .ZN(rc[7]) );
  NOR2_X1 cntrl_inst_U211 ( .A1(cntrl_inst_n115), .A2(cntrl_inst_n155), .ZN(
        cntrl_inst_n83) );
  XNOR2_X1 cntrl_inst_U210 ( .A(kext[131]), .B(cntrl_inst_n107), .ZN(rc[3]) );
  NOR2_X1 cntrl_inst_U209 ( .A1(cntrl_inst_n76), .A2(cntrl_inst_n100), .ZN(
        cntrl_inst_n107) );
  NAND2_X1 cntrl_inst_U208 ( .A1(cntrl_inst_n129), .A2(cntrl_inst_n75), .ZN(
        cntrl_inst_n100) );
  XOR2_X1 cntrl_inst_U207 ( .A(kext[188]), .B(cntrl_inst_n112), .Z(rc[60]) );
  XOR2_X1 cntrl_inst_U206 ( .A(kext[184]), .B(cntrl_inst_n77), .Z(rc[56]) );
  NAND3_X1 cntrl_inst_U205 ( .A1(cntrl_inst_n98), .A2(cntrl_inst_n74), .A3(
        cntrl_inst_n80), .ZN(cntrl_inst_n77) );
  XOR2_X1 cntrl_inst_U204 ( .A(kext[180]), .B(cntrl_inst_n112), .Z(rc[52]) );
  NAND2_X1 cntrl_inst_U203 ( .A1(cntrl_inst_n73), .A2(cntrl_inst_n72), .ZN(
        cntrl_inst_n112) );
  XOR2_X1 cntrl_inst_U202 ( .A(kext[176]), .B(cntrl_inst_n71), .Z(rc[48]) );
  NAND2_X1 cntrl_inst_U201 ( .A1(cntrl_inst_n98), .A2(cntrl_inst_n70), .ZN(
        cntrl_inst_n71) );
  XOR2_X1 cntrl_inst_U200 ( .A(kext[168]), .B(cntrl_inst_n121), .Z(rc[40]) );
  NAND3_X1 cntrl_inst_U199 ( .A1(cntrl_inst_n69), .A2(cntrl_inst_n68), .A3(
        cntrl_inst_n73), .ZN(cntrl_inst_n121) );
  XNOR2_X1 cntrl_inst_U198 ( .A(kext[164]), .B(cntrl_inst_n89), .ZN(rc[36]) );
  NOR2_X1 cntrl_inst_U197 ( .A1(cntrl_inst_n76), .A2(cntrl_inst_n87), .ZN(
        cntrl_inst_n89) );
  XOR2_X1 cntrl_inst_U196 ( .A(kext[160]), .B(cntrl_inst_n67), .Z(rc[32]) );
  NAND3_X1 cntrl_inst_U195 ( .A1(cntrl_inst_n68), .A2(cntrl_inst_n129), .A3(
        cntrl_inst_n84), .ZN(cntrl_inst_n67) );
  XOR2_X1 cntrl_inst_U194 ( .A(kext[156]), .B(cntrl_inst_n94), .Z(rc[28]) );
  NAND3_X1 cntrl_inst_U193 ( .A1(cntrl_inst_n85), .A2(cntrl_inst_n74), .A3(
        cntrl_inst_n80), .ZN(cntrl_inst_n94) );
  XNOR2_X1 cntrl_inst_U192 ( .A(kext[152]), .B(cntrl_inst_n66), .ZN(rc[24]) );
  NOR2_X1 cntrl_inst_U191 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n95), .ZN(
        cntrl_inst_n66) );
  NAND2_X1 cntrl_inst_U190 ( .A1(cntrl_inst_n65), .A2(cntrl_inst_n80), .ZN(
        cntrl_inst_n95) );
  XNOR2_X1 cntrl_inst_U189 ( .A(cntrl_inst_n93), .B(kext[148]), .ZN(rc[20]) );
  XOR2_X1 cntrl_inst_U188 ( .A(kext[144]), .B(cntrl_inst_n120), .Z(rc[16]) );
  NAND2_X1 cntrl_inst_U187 ( .A1(cntrl_inst_n70), .A2(cntrl_inst_n85), .ZN(
        cntrl_inst_n120) );
  NOR2_X1 cntrl_inst_U186 ( .A1(cntrl_inst_n81), .A2(cntrl_inst_n64), .ZN(
        cntrl_inst_n70) );
  XNOR2_X1 cntrl_inst_U185 ( .A(cntrl_inst_n93), .B(kext[140]), .ZN(rc[12]) );
  NOR2_X1 cntrl_inst_U184 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n104), .ZN(
        cntrl_inst_n93) );
  NAND2_X1 cntrl_inst_U183 ( .A1(cntrl_inst_n65), .A2(cntrl_inst_n74), .ZN(
        cntrl_inst_n104) );
  NOR3_X1 cntrl_inst_U182 ( .A1(cntrl_inst_n124), .A2(cntrl_inst_n63), .A3(
        cntrl_inst_n62), .ZN(cntrl_inst_n65) );
  XOR2_X1 cntrl_inst_U181 ( .A(kext[132]), .B(cntrl_inst_n61), .Z(rc[4]) );
  NAND3_X1 cntrl_inst_U180 ( .A1(cntrl_inst_n68), .A2(cntrl_inst_n86), .A3(
        cntrl_inst_n73), .ZN(cntrl_inst_n61) );
  NOR2_X1 cntrl_inst_U179 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n60), .ZN(
        cntrl_inst_n68) );
  XNOR2_X1 cntrl_inst_U178 ( .A(kext[128]), .B(cntrl_inst_n111), .ZN(rc[0]) );
  NOR2_X1 cntrl_inst_U177 ( .A1(cntrl_inst_n91), .A2(cntrl_inst_n87), .ZN(
        cntrl_inst_n111) );
  NAND2_X1 cntrl_inst_U176 ( .A1(cntrl_inst_n73), .A2(cntrl_inst_n75), .ZN(
        cntrl_inst_n87) );
  XOR2_X1 cntrl_inst_U175 ( .A(kext[191]), .B(cntrl_inst_n59), .Z(
        prince_inst_rc2_inv[63]) );
  NAND3_X1 cntrl_inst_U174 ( .A1(cntrl_inst_n58), .A2(cntrl_inst_n57), .A3(
        cntrl_inst_n75), .ZN(cntrl_inst_n59) );
  XNOR2_X1 cntrl_inst_U173 ( .A(kext[160]), .B(cntrl_inst_n56), .ZN(
        prince_inst_rc2_inv[48]) );
  NOR2_X1 cntrl_inst_U172 ( .A1(cntrl_inst_n60), .A2(cntrl_inst_n55), .ZN(
        cntrl_inst_n56) );
  XOR2_X1 cntrl_inst_U171 ( .A(kext[164]), .B(cntrl_inst_n54), .Z(
        prince_inst_rc2_inv[4]) );
  XOR2_X1 cntrl_inst_U170 ( .A(kext[159]), .B(cntrl_inst_n54), .Z(
        prince_inst_rc2_inv[31]) );
  XOR2_X1 cntrl_inst_U169 ( .A(kext[158]), .B(cntrl_inst_n54), .Z(
        prince_inst_rc2_inv[30]) );
  NAND2_X1 cntrl_inst_U168 ( .A1(cntrl_inst_n137), .A2(cntrl_inst_n134), .ZN(
        cntrl_inst_n54) );
  XOR2_X1 cntrl_inst_U167 ( .A(kext[184]), .B(cntrl_inst_n53), .Z(
        prince_inst_rc2_inv[40]) );
  XOR2_X1 cntrl_inst_U166 ( .A(kext[137]), .B(cntrl_inst_n53), .Z(
        prince_inst_rc2_inv[57]) );
  XNOR2_X1 cntrl_inst_U165 ( .A(cntrl_inst_n52), .B(kext[172]), .ZN(
        prince_inst_rc2_inv[44]) );
  XNOR2_X1 cntrl_inst_U164 ( .A(cntrl_inst_n52), .B(kext[145]), .ZN(
        prince_inst_rc2_inv[33]) );
  NOR2_X1 cntrl_inst_U163 ( .A1(cntrl_inst_n91), .A2(cntrl_inst_n51), .ZN(
        cntrl_inst_n52) );
  XOR2_X1 cntrl_inst_U162 ( .A(kext[187]), .B(cntrl_inst_n50), .Z(
        prince_inst_rc2_inv[43]) );
  XOR2_X1 cntrl_inst_U161 ( .A(kext[174]), .B(cntrl_inst_n50), .Z(
        prince_inst_rc2_inv[46]) );
  XOR2_X1 cntrl_inst_U160 ( .A(kext[154]), .B(cntrl_inst_n50), .Z(
        prince_inst_rc2_inv[10]) );
  XOR2_X1 cntrl_inst_U159 ( .A(kext[139]), .B(cntrl_inst_n50), .Z(
        prince_inst_rc2_inv[59]) );
  XOR2_X1 cntrl_inst_U158 ( .A(kext[138]), .B(cntrl_inst_n50), .Z(
        prince_inst_rc2_inv[58]) );
  XNOR2_X1 cntrl_inst_U157 ( .A(cntrl_inst_n69), .B(kext[177]), .ZN(
        prince_inst_rc2_inv[1]) );
  XOR2_X1 cntrl_inst_U156 ( .A(kext[190]), .B(cntrl_inst_n49), .Z(
        prince_inst_rc2_inv[62]) );
  XOR2_X1 cntrl_inst_U155 ( .A(kext[181]), .B(cntrl_inst_n48), .Z(
        prince_inst_rc2_inv[21]) );
  XOR2_X1 cntrl_inst_U154 ( .A(kext[168]), .B(cntrl_inst_n49), .Z(
        prince_inst_rc2_inv[24]) );
  NAND2_X1 cntrl_inst_U153 ( .A1(cntrl_inst_n129), .A2(cntrl_inst_n122), .ZN(
        cntrl_inst_n49) );
  XOR2_X1 cntrl_inst_U152 ( .A(kext[128]), .B(cntrl_inst_n48), .Z(
        prince_inst_rc2_inv[16]) );
  NAND2_X1 cntrl_inst_U151 ( .A1(cntrl_inst_n129), .A2(cntrl_inst_n134), .ZN(
        cntrl_inst_n48) );
  NOR2_X1 cntrl_inst_U150 ( .A1(cntrl_inst_n60), .A2(cntrl_inst_n141), .ZN(
        cntrl_inst_n134) );
  NAND2_X1 cntrl_inst_U149 ( .A1(cntrl_inst_n127), .A2(cntrl_inst_n80), .ZN(
        cntrl_inst_n141) );
  XNOR2_X1 cntrl_inst_U148 ( .A(kext[165]), .B(cntrl_inst_n47), .ZN(
        prince_inst_rc2_inv[5]) );
  XNOR2_X1 cntrl_inst_U147 ( .A(kext[148]), .B(cntrl_inst_n47), .ZN(
        prince_inst_rc2_inv[52]) );
  XNOR2_X1 cntrl_inst_U146 ( .A(kext[140]), .B(cntrl_inst_n47), .ZN(
        prince_inst_rc2_inv[12]) );
  NOR3_X1 cntrl_inst_U145 ( .A1(cntrl_inst_n64), .A2(cntrl_inst_n46), .A3(
        cntrl_inst_n147), .ZN(cntrl_inst_n47) );
  NAND3_X1 cntrl_inst_U144 ( .A1(cntrl_inst_n45), .A2(cntrl_inst_n80), .A3(
        cntrl_inst_n78), .ZN(cntrl_inst_n147) );
  INV_X1 cntrl_inst_U143 ( .A(cntrl_inst_n152), .ZN(cntrl_inst_n45) );
  XNOR2_X1 cntrl_inst_U142 ( .A(cntrl_inst_n44), .B(kext[153]), .ZN(
        prince_inst_rc2_inv[9]) );
  XNOR2_X1 cntrl_inst_U141 ( .A(cntrl_inst_n116), .B(kext[129]), .ZN(
        prince_inst_rc2_inv[17]) );
  XNOR2_X1 cntrl_inst_U140 ( .A(cntrl_inst_n43), .B(kext[188]), .ZN(
        prince_inst_rc2_inv[60]) );
  XNOR2_X1 cntrl_inst_U139 ( .A(cntrl_inst_n43), .B(kext[185]), .ZN(
        prince_inst_rc2_inv[41]) );
  XNOR2_X1 cntrl_inst_U138 ( .A(kext[180]), .B(cntrl_inst_n43), .ZN(
        prince_inst_rc2_inv[20]) );
  NOR2_X1 cntrl_inst_U137 ( .A1(cntrl_inst_n42), .A2(cntrl_inst_n62), .ZN(
        cntrl_inst_n43) );
  XOR2_X1 cntrl_inst_U136 ( .A(kext[166]), .B(cntrl_inst_n41), .Z(
        prince_inst_rc2_inv[6]) );
  XOR2_X1 cntrl_inst_U135 ( .A(kext[156]), .B(cntrl_inst_n41), .Z(
        prince_inst_rc2_inv[28]) );
  XOR2_X1 cntrl_inst_U134 ( .A(kext[133]), .B(cntrl_inst_n41), .Z(
        prince_inst_rc2_inv[37]) );
  XOR2_X1 cntrl_inst_U133 ( .A(kext[132]), .B(cntrl_inst_n39), .Z(
        prince_inst_rc2_inv[36]) );
  NAND2_X1 cntrl_inst_U132 ( .A1(cntrl_inst_n135), .A2(cntrl_inst_n122), .ZN(
        cntrl_inst_n39) );
  NOR3_X1 cntrl_inst_U131 ( .A1(cntrl_inst_n152), .A2(cntrl_inst_n76), .A3(
        cntrl_inst_n60), .ZN(cntrl_inst_n122) );
  XNOR2_X1 cntrl_inst_U130 ( .A(kext[182]), .B(cntrl_inst_n38), .ZN(
        prince_inst_rc2_inv[22]) );
  XNOR2_X1 cntrl_inst_U129 ( .A(kext[170]), .B(cntrl_inst_n38), .ZN(
        prince_inst_rc2_inv[26]) );
  XOR2_X1 cntrl_inst_U128 ( .A(kext[157]), .B(cntrl_inst_n37), .Z(
        prince_inst_rc2_inv[29]) );
  NAND2_X1 cntrl_inst_U127 ( .A1(cntrl_inst_n69), .A2(cntrl_inst_n35), .ZN(
        cntrl_inst_n37) );
  XNOR2_X1 cntrl_inst_U126 ( .A(kext[141]), .B(cntrl_inst_n34), .ZN(
        prince_inst_rc2_inv[13]) );
  NOR3_X1 cntrl_inst_U125 ( .A1(cntrl_inst_n91), .A2(cntrl_inst_n51), .A3(
        cntrl_inst_n62), .ZN(cntrl_inst_n34) );
  XOR2_X1 cntrl_inst_U124 ( .A(kext[142]), .B(cntrl_inst_n33), .Z(
        prince_inst_rc2_inv[14]) );
  NAND4_X1 cntrl_inst_U123 ( .A1(cntrl_inst_n57), .A2(cntrl_inst_n127), .A3(
        cntrl_inst_n80), .A4(cntrl_inst_n117), .ZN(cntrl_inst_n33) );
  NAND2_X1 cntrl_inst_U122 ( .A1(cntrl_inst_n32), .A2(cntrl_inst_n155), .ZN(
        cntrl_inst_n117) );
  XNOR2_X1 cntrl_inst_U121 ( .A(cntrl_inst_n31), .B(kext[144]), .ZN(
        prince_inst_rc2_inv[32]) );
  XNOR2_X1 cntrl_inst_U120 ( .A(cntrl_inst_n30), .B(kext[149]), .ZN(
        prince_inst_rc2_inv[53]) );
  NOR2_X1 cntrl_inst_U119 ( .A1(cntrl_inst_n55), .A2(cntrl_inst_n81), .ZN(
        cntrl_inst_n30) );
  NAND2_X1 cntrl_inst_U118 ( .A1(cntrl_inst_n137), .A2(cntrl_inst_n58), .ZN(
        cntrl_inst_n55) );
  NOR2_X1 cntrl_inst_U117 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n29), .ZN(
        cntrl_inst_n137) );
  XOR2_X1 cntrl_inst_U116 ( .A(kext[150]), .B(cntrl_inst_n28), .Z(
        prince_inst_rc2_inv[54]) );
  NAND4_X1 cntrl_inst_U115 ( .A1(cntrl_inst_n27), .A2(cntrl_inst_n73), .A3(
        cntrl_inst_n127), .A4(cntrl_inst_n26), .ZN(cntrl_inst_n28) );
  INV_X1 cntrl_inst_U114 ( .A(cntrl_inst_n46), .ZN(cntrl_inst_n26) );
  XNOR2_X1 cntrl_inst_U113 ( .A(cntrl_inst_n35), .B(kext[151]), .ZN(
        prince_inst_rc2_inv[55]) );
  XOR2_X1 cntrl_inst_U112 ( .A(kext[130]), .B(cntrl_inst_n25), .Z(
        prince_inst_rc2_inv[18]) );
  XOR2_X1 cntrl_inst_U111 ( .A(kext[161]), .B(cntrl_inst_n24), .Z(
        prince_inst_rc2_inv[49]) );
  XOR2_X1 cntrl_inst_U110 ( .A(kext[162]), .B(cntrl_inst_n25), .Z(
        prince_inst_rc2_inv[50]) );
  NAND3_X1 cntrl_inst_U109 ( .A1(cntrl_inst_n58), .A2(cntrl_inst_n129), .A3(
        cntrl_inst_n27), .ZN(cntrl_inst_n25) );
  NOR2_X1 cntrl_inst_U108 ( .A1(cntrl_inst_n29), .A2(cntrl_inst_n46), .ZN(
        cntrl_inst_n129) );
  XNOR2_X1 cntrl_inst_U107 ( .A(cntrl_inst_n23), .B(kext[163]), .ZN(
        prince_inst_rc2_inv[51]) );
  XNOR2_X1 cntrl_inst_U106 ( .A(kext[169]), .B(cntrl_inst_n23), .ZN(
        prince_inst_rc2_inv[25]) );
  NOR2_X1 cntrl_inst_U105 ( .A1(cntrl_inst_n62), .A2(cntrl_inst_n50), .ZN(
        cntrl_inst_n23) );
  NAND2_X1 cntrl_inst_U104 ( .A1(cntrl_inst_n69), .A2(cntrl_inst_n38), .ZN(
        cntrl_inst_n50) );
  XNOR2_X1 cntrl_inst_U103 ( .A(cntrl_inst_n22), .B(kext[175]), .ZN(
        prince_inst_rc2_inv[47]) );
  NOR2_X1 cntrl_inst_U102 ( .A1(cntrl_inst_n62), .A2(cntrl_inst_n91), .ZN(
        cntrl_inst_n22) );
  XNOR2_X1 cntrl_inst_U101 ( .A(cntrl_inst_n35), .B(kext[186]), .ZN(
        prince_inst_rc2_inv[42]) );
  NOR2_X1 cntrl_inst_U100 ( .A1(cntrl_inst_n51), .A2(cntrl_inst_n41), .ZN(
        cntrl_inst_n35) );
  NAND2_X1 cntrl_inst_U99 ( .A1(cntrl_inst_n116), .A2(cntrl_inst_n38), .ZN(
        cntrl_inst_n41) );
  XNOR2_X1 cntrl_inst_U98 ( .A(kext[189]), .B(cntrl_inst_n31), .ZN(
        prince_inst_rc2_inv[61]) );
  NOR2_X1 cntrl_inst_U97 ( .A1(cntrl_inst_n42), .A2(cntrl_inst_n51), .ZN(
        cntrl_inst_n31) );
  INV_X1 cntrl_inst_U96 ( .A(cntrl_inst_n38), .ZN(cntrl_inst_n42) );
  NAND2_X1 cntrl_inst_U95 ( .A1(cntrl_inst_n21), .A2(cntrl_inst_n20), .ZN(
        cntrl_inst_n38) );
  XOR2_X1 cntrl_inst_U94 ( .A(kext[134]), .B(cntrl_inst_n24), .Z(
        prince_inst_rc2_inv[38]) );
  NAND3_X1 cntrl_inst_U93 ( .A1(cntrl_inst_n58), .A2(cntrl_inst_n27), .A3(
        cntrl_inst_n135), .ZN(cntrl_inst_n24) );
  NOR3_X1 cntrl_inst_U92 ( .A1(cntrl_inst_n152), .A2(cntrl_inst_n124), .A3(
        cntrl_inst_n64), .ZN(cntrl_inst_n58) );
  NOR2_X1 cntrl_inst_U91 ( .A1(cntrl_inst_n108), .A2(cntrl_inst_n127), .ZN(
        cntrl_inst_n152) );
  NAND2_X1 cntrl_inst_U90 ( .A1(cntrl_inst_n32), .A2(cntrl_inst_n109), .ZN(
        cntrl_inst_n127) );
  NOR2_X1 cntrl_inst_U89 ( .A1(cntrl_inst_n20), .A2(cntrl_inst_n19), .ZN(
        cntrl_inst_n109) );
  XNOR2_X1 cntrl_inst_U88 ( .A(cntrl_inst_n18), .B(kext[136]), .ZN(
        prince_inst_rc2_inv[56]) );
  NOR2_X1 cntrl_inst_U87 ( .A1(cntrl_inst_n53), .A2(cntrl_inst_n51), .ZN(
        cntrl_inst_n18) );
  OR2_X1 cntrl_inst_U86 ( .A1(cntrl_inst_n29), .A2(cntrl_inst_n103), .ZN(
        cntrl_inst_n51) );
  NOR2_X1 cntrl_inst_U85 ( .A1(cntrl_inst_n135), .A2(cntrl_inst_n17), .ZN(
        cntrl_inst_n103) );
  NAND2_X1 cntrl_inst_U84 ( .A1(cntrl_inst_n116), .A2(cntrl_inst_n44), .ZN(
        cntrl_inst_n53) );
  INV_X1 cntrl_inst_U83 ( .A(cntrl_inst_n62), .ZN(cntrl_inst_n44) );
  NAND2_X1 cntrl_inst_U82 ( .A1(cntrl_inst_n27), .A2(cntrl_inst_n125), .ZN(
        cntrl_inst_n62) );
  INV_X1 cntrl_inst_U81 ( .A(cntrl_inst_n81), .ZN(cntrl_inst_n27) );
  NOR2_X1 cntrl_inst_U80 ( .A1(cntrl_inst_n17), .A2(cntrl_inst_n86), .ZN(
        cntrl_inst_n81) );
  NOR2_X1 cntrl_inst_U79 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n46), .ZN(
        cntrl_inst_n116) );
  XNOR2_X1 cntrl_inst_U78 ( .A(cntrl_inst_n90), .B(kext[138]), .ZN(rc[10]) );
  XNOR2_X1 cntrl_inst_U77 ( .A(cntrl_inst_n90), .B(kext[139]), .ZN(rc[11]) );
  XNOR2_X1 cntrl_inst_U76 ( .A(kext[142]), .B(cntrl_inst_n16), .ZN(rc[14]) );
  NOR4_X1 cntrl_inst_U75 ( .A1(cntrl_inst_n124), .A2(cntrl_inst_n76), .A3(
        cntrl_inst_n142), .A4(cntrl_inst_n63), .ZN(cntrl_inst_n16) );
  XOR2_X1 cntrl_inst_U74 ( .A(kext[145]), .B(cntrl_inst_n15), .Z(rc[17]) );
  XOR2_X1 cntrl_inst_U73 ( .A(kext[129]), .B(cntrl_inst_n14), .Z(rc[1]) );
  NAND2_X1 cntrl_inst_U72 ( .A1(cntrl_inst_n74), .A2(cntrl_inst_n80), .ZN(
        cntrl_inst_n14) );
  NAND2_X1 cntrl_inst_U71 ( .A1(cntrl_inst_n76), .A2(cntrl_inst_n20), .ZN(
        cntrl_inst_n80) );
  INV_X1 cntrl_inst_U70 ( .A(cntrl_inst_n84), .ZN(cntrl_inst_n76) );
  INV_X1 cntrl_inst_U69 ( .A(cntrl_inst_n148), .ZN(cntrl_inst_n74) );
  XOR2_X1 cntrl_inst_U68 ( .A(kext[149]), .B(cntrl_inst_n13), .Z(rc[21]) );
  NAND2_X1 cntrl_inst_U67 ( .A1(cntrl_inst_n84), .A2(cntrl_inst_n12), .ZN(
        cntrl_inst_n13) );
  XNOR2_X1 cntrl_inst_U66 ( .A(kext[150]), .B(cntrl_inst_n11), .ZN(rc[22]) );
  NOR4_X1 cntrl_inst_U65 ( .A1(cntrl_inst_n142), .A2(cntrl_inst_n46), .A3(
        cntrl_inst_n63), .A4(cntrl_inst_n91), .ZN(cntrl_inst_n11) );
  INV_X1 cntrl_inst_U64 ( .A(cntrl_inst_n69), .ZN(cntrl_inst_n91) );
  INV_X1 cntrl_inst_U63 ( .A(cntrl_inst_n75), .ZN(cntrl_inst_n142) );
  XNOR2_X1 cntrl_inst_U62 ( .A(cntrl_inst_n98), .B(kext[153]), .ZN(rc[25]) );
  XNOR2_X1 cntrl_inst_U61 ( .A(cntrl_inst_n90), .B(kext[154]), .ZN(rc[26]) );
  XNOR2_X1 cntrl_inst_U60 ( .A(cntrl_inst_n10), .B(kext[157]), .ZN(rc[29]) );
  NOR2_X1 cntrl_inst_U59 ( .A1(cntrl_inst_n21), .A2(cntrl_inst_n153), .ZN(
        cntrl_inst_n10) );
  XOR2_X1 cntrl_inst_U58 ( .A(kext[130]), .B(cntrl_inst_n9), .Z(rc[2]) );
  XOR2_X1 cntrl_inst_U57 ( .A(kext[161]), .B(cntrl_inst_n8), .Z(rc[33]) );
  XOR2_X1 cntrl_inst_U56 ( .A(kext[162]), .B(cntrl_inst_n9), .Z(rc[34]) );
  NAND2_X1 cntrl_inst_U55 ( .A1(cntrl_inst_n69), .A2(cntrl_inst_n12), .ZN(
        cntrl_inst_n9) );
  NOR2_X1 cntrl_inst_U54 ( .A1(cntrl_inst_n64), .A2(cntrl_inst_n148), .ZN(
        cntrl_inst_n69) );
  NOR2_X1 cntrl_inst_U53 ( .A1(cntrl_inst_n20), .A2(cntrl_inst_n86), .ZN(
        cntrl_inst_n148) );
  NOR2_X1 cntrl_inst_U52 ( .A1(cntrl_inst_n20), .A2(cntrl_inst_n84), .ZN(
        cntrl_inst_n64) );
  XNOR2_X1 cntrl_inst_U51 ( .A(cntrl_inst_n85), .B(kext[170]), .ZN(rc[42]) );
  XOR2_X1 cntrl_inst_U50 ( .A(kext[172]), .B(cntrl_inst_n15), .Z(rc[44]) );
  NAND2_X1 cntrl_inst_U49 ( .A1(cntrl_inst_n144), .A2(cntrl_inst_n78), .ZN(
        cntrl_inst_n15) );
  NAND2_X1 cntrl_inst_U48 ( .A1(cntrl_inst_n153), .A2(cntrl_inst_n20), .ZN(
        cntrl_inst_n78) );
  XNOR2_X1 cntrl_inst_U47 ( .A(cntrl_inst_n90), .B(kext[174]), .ZN(rc[46]) );
  XNOR2_X1 cntrl_inst_U46 ( .A(cntrl_inst_n85), .B(kext[182]), .ZN(rc[54]) );
  NOR2_X1 cntrl_inst_U45 ( .A1(cntrl_inst_n124), .A2(cntrl_inst_n46), .ZN(
        cntrl_inst_n85) );
  NOR2_X1 cntrl_inst_U44 ( .A1(cntrl_inst_n20), .A2(cntrl_inst_n135), .ZN(
        cntrl_inst_n46) );
  INV_X1 cntrl_inst_U43 ( .A(cntrl_inst_n132), .ZN(cntrl_inst_n135) );
  INV_X1 cntrl_inst_U42 ( .A(cntrl_inst_n17), .ZN(cntrl_inst_n20) );
  XNOR2_X1 cntrl_inst_U41 ( .A(cntrl_inst_n90), .B(kext[187]), .ZN(rc[59]) );
  NOR2_X1 cntrl_inst_U40 ( .A1(cntrl_inst_n32), .A2(cntrl_inst_n7), .ZN(
        cntrl_inst_n132) );
  NOR2_X1 cntrl_inst_U39 ( .A1(cntrl_inst_n6), .A2(cntrl_inst_n73), .ZN(
        cntrl_inst_n124) );
  XOR2_X1 cntrl_inst_U38 ( .A(kext[134]), .B(cntrl_inst_n8), .Z(rc[6]) );
  NAND2_X1 cntrl_inst_U37 ( .A1(cntrl_inst_n12), .A2(cntrl_inst_n86), .ZN(
        cntrl_inst_n8) );
  AND3_X1 cntrl_inst_U36 ( .A1(cntrl_inst_n57), .A2(cntrl_inst_n125), .A3(
        cntrl_inst_n72), .ZN(cntrl_inst_n12) );
  INV_X1 cntrl_inst_U35 ( .A(cntrl_inst_n60), .ZN(cntrl_inst_n125) );
  NOR2_X1 cntrl_inst_U34 ( .A1(cntrl_inst_n108), .A2(cntrl_inst_n75), .ZN(
        cntrl_inst_n60) );
  NAND2_X1 cntrl_inst_U33 ( .A1(cntrl_inst_n155), .A2(cntrl_inst_n114), .ZN(
        cntrl_inst_n75) );
  NOR2_X1 cntrl_inst_U32 ( .A1(cntrl_inst_n17), .A2(cntrl_inst_n19), .ZN(
        cntrl_inst_n155) );
  INV_X1 cntrl_inst_U31 ( .A(cntrl_inst_n149), .ZN(cntrl_inst_n57) );
  NAND2_X1 cntrl_inst_U30 ( .A1(cntrl_inst_n17), .A2(cntrl_inst_n21), .ZN(
        cntrl_inst_n144) );
  XOR2_X1 cntrl_inst_U29 ( .A(kext[136]), .B(cntrl_inst_n5), .Z(rc[8]) );
  NAND3_X1 cntrl_inst_U28 ( .A1(cntrl_inst_n98), .A2(cntrl_inst_n86), .A3(
        cntrl_inst_n84), .ZN(cntrl_inst_n5) );
  NAND2_X1 cntrl_inst_U27 ( .A1(cntrl_inst_n21), .A2(cntrl_inst_n114), .ZN(
        cntrl_inst_n84) );
  NOR2_X1 cntrl_inst_U26 ( .A1(cntrl_inst_n6), .A2(cntrl_inst_n108), .ZN(
        cntrl_inst_n21) );
  NAND2_X1 cntrl_inst_U25 ( .A1(cntrl_inst_n153), .A2(cntrl_inst_n32), .ZN(
        cntrl_inst_n86) );
  INV_X1 cntrl_inst_U24 ( .A(cntrl_inst_n7), .ZN(cntrl_inst_n153) );
  NAND2_X1 cntrl_inst_U23 ( .A1(cntrl_inst_n108), .A2(cntrl_inst_n6), .ZN(
        cntrl_inst_n7) );
  NOR2_X1 cntrl_inst_U22 ( .A1(cntrl_inst_n29), .A2(cntrl_inst_n63), .ZN(
        cntrl_inst_n98) );
  NOR2_X1 cntrl_inst_U21 ( .A1(cntrl_inst_n6), .A2(cntrl_inst_n72), .ZN(
        cntrl_inst_n63) );
  NAND3_X1 cntrl_inst_U20 ( .A1(cntrl_inst_n17), .A2(cntrl_inst_n108), .A3(
        cntrl_inst_n114), .ZN(cntrl_inst_n72) );
  INV_X1 cntrl_inst_U19 ( .A(cntrl_inst_n32), .ZN(cntrl_inst_n114) );
  NOR2_X1 cntrl_inst_U18 ( .A1(cntrl_inst_n19), .A2(cntrl_inst_n73), .ZN(
        cntrl_inst_n29) );
  NAND2_X1 cntrl_inst_U17 ( .A1(cntrl_inst_n32), .A2(cntrl_inst_n115), .ZN(
        cntrl_inst_n73) );
  NOR2_X1 cntrl_inst_U16 ( .A1(cntrl_inst_n17), .A2(cntrl_inst_n108), .ZN(
        cntrl_inst_n115) );
  XNOR2_X1 cntrl_inst_U15 ( .A(enc), .B(inv_sig), .ZN(cntrl_inst_n108) );
  XOR2_X1 cntrl_inst_U14 ( .A(cntrl_inst_n40), .B(enc), .Z(cntrl_inst_n17) );
  XOR2_X1 cntrl_inst_U13 ( .A(enc), .B(cntrl_inst_counter_0_), .Z(
        cntrl_inst_n32) );
  INV_X1 cntrl_inst_U12 ( .A(cntrl_inst_n6), .ZN(cntrl_inst_n19) );
  XOR2_X1 cntrl_inst_U11 ( .A(enc), .B(cntrl_inst_n36), .Z(cntrl_inst_n6) );
  INV_X4 cntrl_inst_U10 ( .A(done), .ZN(en_sig) );
  NAND4_X1 cntrl_inst_U9 ( .A1(inv_sig), .A2(cntrl_inst_n36), .A3(en), .A4(
        cntrl_inst_n167), .ZN(cntrl_inst_n4) );
  NOR2_X2 cntrl_inst_U8 ( .A1(cntrl_inst_counter_0_), .A2(cntrl_inst_n157), 
        .ZN(done) );
  NAND3_X1 cntrl_inst_U7 ( .A1(cntrl_inst_n168), .A2(cntrl_inst_n166), .A3(
        cntrl_inst_n165), .ZN(cntrl_inst_n157) );
  NOR2_X1 cntrl_inst_U6 ( .A1(cntrl_inst_n40), .A2(cntrl_inst_n4), .ZN(
        start_sig) );
  NOR2_X2 cntrl_inst_U5 ( .A1(cntrl_inst_n114), .A2(cntrl_inst_n144), .ZN(
        cntrl_inst_n149) );
  NOR3_X2 cntrl_inst_U4 ( .A1(cntrl_inst_n149), .A2(cntrl_inst_n124), .A3(
        cntrl_inst_n132), .ZN(cntrl_inst_n90) );
  INV_X1 cntrl_inst_U3 ( .A(rst), .ZN(cntrl_inst_n3) );
  DFF_X1 cntrl_inst_counter_reg_2_ ( .D(cntrl_inst_n208), .CK(clk), .Q(
        cntrl_inst_n166), .QN(cntrl_inst_n36) );
  DFF_X1 cntrl_inst_counter_reg_1_ ( .D(cntrl_inst_n207), .CK(clk), .Q(
        cntrl_inst_n168), .QN(cntrl_inst_n40) );
  DFF_X1 cntrl_inst_counter_reg_3_ ( .D(cntrl_inst_n209), .CK(clk), .Q(
        cntrl_inst_n165), .QN(inv_sig) );
  DFF_X1 cntrl_inst_counter_reg_0_ ( .D(cntrl_inst_n210), .CK(clk), .Q(
        cntrl_inst_counter_0_), .QN(cntrl_inst_n167) );
  INV_X1 prince_inst_U16 ( .A(inv_sig2), .ZN(prince_inst_n25) );
  INV_X1 prince_inst_U15 ( .A(prince_inst_n25), .ZN(prince_inst_n20) );
  INV_X1 prince_inst_U14 ( .A(prince_inst_n25), .ZN(prince_inst_n21) );
  INV_X1 prince_inst_U13 ( .A(prince_inst_n34), .ZN(prince_inst_n26) );
  INV_X1 prince_inst_U12 ( .A(prince_inst_n25), .ZN(prince_inst_n22) );
  INV_X1 prince_inst_U11 ( .A(prince_inst_n25), .ZN(prince_inst_n23) );
  INV_X1 prince_inst_U10 ( .A(prince_inst_n25), .ZN(prince_inst_n19) );
  INV_X1 prince_inst_U9 ( .A(prince_inst_n34), .ZN(prince_inst_n27) );
  INV_X1 prince_inst_U8 ( .A(prince_inst_n34), .ZN(prince_inst_n28) );
  INV_X1 prince_inst_U7 ( .A(prince_inst_n25), .ZN(prince_inst_n24) );
  INV_X1 prince_inst_U6 ( .A(prince_inst_n34), .ZN(prince_inst_n29) );
  INV_X1 prince_inst_U5 ( .A(prince_inst_n34), .ZN(prince_inst_n32) );
  INV_X1 prince_inst_U4 ( .A(prince_inst_n34), .ZN(prince_inst_n31) );
  INV_X1 prince_inst_U3 ( .A(prince_inst_n34), .ZN(prince_inst_n30) );
  INV_X1 prince_inst_U2 ( .A(prince_inst_n34), .ZN(prince_inst_n33) );
  INV_X1 prince_inst_U1 ( .A(inv_sig), .ZN(prince_inst_n34) );
  XOR2_X1 prince_inst_S_0__x_U1 ( .A(rc[0]), .B(prince_inst_srin_x[32]), .Z(
        prince_inst_xout_x[0]) );
  XOR2_X1 prince_inst_S_0__srx_U1 ( .A(prince_inst_rc2_inv[0]), .B(
        prince_inst_sout_x[0]), .Z(final_x[48]) );
  MUX2_X1 prince_inst_S_0__mux_inv_x1_U1 ( .A(prince_inst_srin_x[0]), .B(
        prince_inst_xout_x[0]), .S(prince_inst_n30), .Z(prince_inst_sin_x[0])
         );
  MUX2_X1 prince_inst_S_0__mux_inv_y1_U1 ( .A(prince_inst_srin_y[0]), .B(
        prince_inst_srin_y[32]), .S(prince_inst_n30), .Z(prince_inst_sin_y[0])
         );
  MUX2_X1 prince_inst_S_0__mux_inv_x2_U1 ( .A(final_x[48]), .B(
        prince_inst_sout_x[0]), .S(prince_inst_n23), .Z(prince_inst_min_x[0])
         );
  MUX2_X1 prince_inst_S_0__mux_inv_y2_U1 ( .A(final_y[48]), .B(final_y[48]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[0]) );
  XOR2_X1 prince_inst_S_1__x_U1 ( .A(rc[1]), .B(prince_inst_srin_x[33]), .Z(
        prince_inst_xout_x[1]) );
  XOR2_X1 prince_inst_S_1__srx_U1 ( .A(prince_inst_rc2_inv[1]), .B(
        prince_inst_sout_x[1]), .Z(final_x[49]) );
  MUX2_X1 prince_inst_S_1__mux_inv_x1_U1 ( .A(prince_inst_srin_x[1]), .B(
        prince_inst_xout_x[1]), .S(prince_inst_n32), .Z(prince_inst_sin_x[1])
         );
  MUX2_X1 prince_inst_S_1__mux_inv_y1_U1 ( .A(prince_inst_srin_y[1]), .B(
        prince_inst_srin_y[33]), .S(prince_inst_n33), .Z(prince_inst_sin_y[1])
         );
  MUX2_X1 prince_inst_S_1__mux_inv_x2_U1 ( .A(final_x[49]), .B(
        prince_inst_sout_x[1]), .S(prince_inst_n19), .Z(prince_inst_min_x[1])
         );
  MUX2_X1 prince_inst_S_1__mux_inv_y2_U1 ( .A(final_y[49]), .B(final_y[49]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[1]) );
  XOR2_X1 prince_inst_S_2__x_U1 ( .A(rc[2]), .B(prince_inst_srin_x[34]), .Z(
        prince_inst_xout_x[2]) );
  XOR2_X1 prince_inst_S_2__srx_U1 ( .A(prince_inst_rc2_inv[2]), .B(
        prince_inst_sout_x[2]), .Z(final_x[50]) );
  MUX2_X1 prince_inst_S_2__mux_inv_x1_U1 ( .A(prince_inst_srin_x[2]), .B(
        prince_inst_xout_x[2]), .S(prince_inst_n33), .Z(prince_inst_sin_x[2])
         );
  MUX2_X1 prince_inst_S_2__mux_inv_y1_U1 ( .A(prince_inst_srin_y[2]), .B(
        prince_inst_srin_y[34]), .S(prince_inst_n33), .Z(prince_inst_sin_y[2])
         );
  MUX2_X1 prince_inst_S_2__mux_inv_x2_U1 ( .A(final_x[50]), .B(
        prince_inst_sout_x[2]), .S(prince_inst_n19), .Z(prince_inst_min_x[2])
         );
  MUX2_X1 prince_inst_S_2__mux_inv_y2_U1 ( .A(final_y[50]), .B(final_y[50]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[2]) );
  XOR2_X1 prince_inst_S_3__x_U1 ( .A(rc[3]), .B(prince_inst_srin_x[35]), .Z(
        prince_inst_xout_x[3]) );
  XOR2_X1 prince_inst_S_3__srx_U1 ( .A(prince_inst_rc2_inv[3]), .B(
        prince_inst_sout_x[3]), .Z(final_x[51]) );
  MUX2_X1 prince_inst_S_3__mux_inv_x1_U1 ( .A(prince_inst_srin_x[3]), .B(
        prince_inst_xout_x[3]), .S(prince_inst_n33), .Z(prince_inst_sin_x[3])
         );
  MUX2_X1 prince_inst_S_3__mux_inv_y1_U1 ( .A(prince_inst_srin_y[3]), .B(
        prince_inst_srin_y[35]), .S(prince_inst_n33), .Z(prince_inst_sin_y[3])
         );
  MUX2_X1 prince_inst_S_3__mux_inv_x2_U1 ( .A(final_x[51]), .B(
        prince_inst_sout_x[3]), .S(prince_inst_n19), .Z(prince_inst_min_x[3])
         );
  MUX2_X1 prince_inst_S_3__mux_inv_y2_U1 ( .A(final_y[51]), .B(final_y[51]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[3]) );
  XOR2_X1 prince_inst_S_4__x_U1 ( .A(rc[4]), .B(prince_inst_srin_x[4]), .Z(
        prince_inst_xout_x[4]) );
  XOR2_X1 prince_inst_S_4__srx_U1 ( .A(prince_inst_rc2_inv[4]), .B(
        prince_inst_sout_x[4]), .Z(final_x[36]) );
  MUX2_X1 prince_inst_S_4__mux_inv_x1_U1 ( .A(prince_inst_srin_x[4]), .B(
        prince_inst_xout_x[4]), .S(prince_inst_n33), .Z(prince_inst_sin_x[4])
         );
  MUX2_X1 prince_inst_S_4__mux_inv_y1_U1 ( .A(prince_inst_srin_y[4]), .B(
        prince_inst_srin_y[4]), .S(prince_inst_n33), .Z(prince_inst_sin_y[4])
         );
  MUX2_X1 prince_inst_S_4__mux_inv_x2_U1 ( .A(final_x[36]), .B(
        prince_inst_sout_x[4]), .S(prince_inst_n19), .Z(prince_inst_min_x[4])
         );
  MUX2_X1 prince_inst_S_4__mux_inv_y2_U1 ( .A(final_y[36]), .B(final_y[36]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[4]) );
  XOR2_X1 prince_inst_S_5__x_U1 ( .A(rc[5]), .B(prince_inst_srin_x[5]), .Z(
        prince_inst_xout_x[5]) );
  XOR2_X1 prince_inst_S_5__srx_U1 ( .A(prince_inst_rc2_inv[5]), .B(
        prince_inst_sout_x[5]), .Z(final_x[37]) );
  MUX2_X1 prince_inst_S_5__mux_inv_x1_U1 ( .A(prince_inst_srin_x[5]), .B(
        prince_inst_xout_x[5]), .S(prince_inst_n33), .Z(prince_inst_sin_x[5])
         );
  MUX2_X1 prince_inst_S_5__mux_inv_y1_U1 ( .A(prince_inst_srin_y[5]), .B(
        prince_inst_srin_y[5]), .S(prince_inst_n28), .Z(prince_inst_sin_y[5])
         );
  MUX2_X1 prince_inst_S_5__mux_inv_x2_U1 ( .A(final_x[37]), .B(
        prince_inst_sout_x[5]), .S(prince_inst_n19), .Z(prince_inst_min_x[5])
         );
  MUX2_X1 prince_inst_S_5__mux_inv_y2_U1 ( .A(final_y[37]), .B(final_y[37]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[5]) );
  XOR2_X1 prince_inst_S_6__x_U1 ( .A(rc[6]), .B(prince_inst_srin_x[6]), .Z(
        prince_inst_xout_x[6]) );
  XOR2_X1 prince_inst_S_6__srx_U1 ( .A(prince_inst_rc2_inv[6]), .B(
        prince_inst_sout_x[6]), .Z(final_x[38]) );
  MUX2_X1 prince_inst_S_6__mux_inv_x1_U1 ( .A(prince_inst_srin_x[6]), .B(
        prince_inst_xout_x[6]), .S(prince_inst_n27), .Z(prince_inst_sin_x[6])
         );
  MUX2_X1 prince_inst_S_6__mux_inv_y1_U1 ( .A(prince_inst_srin_y[6]), .B(
        prince_inst_srin_y[6]), .S(prince_inst_n31), .Z(prince_inst_sin_y[6])
         );
  MUX2_X1 prince_inst_S_6__mux_inv_x2_U1 ( .A(final_x[38]), .B(
        prince_inst_sout_x[6]), .S(prince_inst_n19), .Z(prince_inst_min_x[6])
         );
  MUX2_X1 prince_inst_S_6__mux_inv_y2_U1 ( .A(final_y[38]), .B(final_y[38]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[6]) );
  XOR2_X1 prince_inst_S_7__x_U1 ( .A(rc[7]), .B(prince_inst_srin_x[7]), .Z(
        prince_inst_xout_x[7]) );
  XOR2_X1 prince_inst_S_7__srx_U1 ( .A(prince_inst_rc2_inv[7]), .B(
        prince_inst_sout_x[7]), .Z(final_x[39]) );
  MUX2_X1 prince_inst_S_7__mux_inv_x1_U1 ( .A(prince_inst_srin_x[7]), .B(
        prince_inst_xout_x[7]), .S(prince_inst_n32), .Z(prince_inst_sin_x[7])
         );
  MUX2_X1 prince_inst_S_7__mux_inv_y1_U1 ( .A(prince_inst_srin_y[7]), .B(
        prince_inst_srin_y[7]), .S(prince_inst_n30), .Z(prince_inst_sin_y[7])
         );
  MUX2_X1 prince_inst_S_7__mux_inv_x2_U1 ( .A(final_x[39]), .B(
        prince_inst_sout_x[7]), .S(prince_inst_n19), .Z(prince_inst_min_x[7])
         );
  MUX2_X1 prince_inst_S_7__mux_inv_y2_U1 ( .A(final_y[39]), .B(final_y[39]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[7]) );
  XOR2_X1 prince_inst_S_8__x_U1 ( .A(rc[8]), .B(prince_inst_srin_x[40]), .Z(
        prince_inst_xout_x[8]) );
  XOR2_X1 prince_inst_S_8__srx_U1 ( .A(prince_inst_rc2_inv[8]), .B(
        prince_inst_sout_x[8]), .Z(final_x[24]) );
  MUX2_X1 prince_inst_S_8__mux_inv_x1_U1 ( .A(prince_inst_srin_x[8]), .B(
        prince_inst_xout_x[8]), .S(prince_inst_n26), .Z(prince_inst_sin_x[8])
         );
  MUX2_X1 prince_inst_S_8__mux_inv_y1_U1 ( .A(prince_inst_srin_y[8]), .B(
        prince_inst_srin_y[40]), .S(prince_inst_n29), .Z(prince_inst_sin_y[8])
         );
  MUX2_X1 prince_inst_S_8__mux_inv_x2_U1 ( .A(final_x[24]), .B(
        prince_inst_sout_x[8]), .S(prince_inst_n19), .Z(prince_inst_min_x[8])
         );
  MUX2_X1 prince_inst_S_8__mux_inv_y2_U1 ( .A(final_y[24]), .B(final_y[24]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[8]) );
  XOR2_X1 prince_inst_S_9__x_U1 ( .A(rc[9]), .B(prince_inst_srin_x[41]), .Z(
        prince_inst_xout_x[9]) );
  XOR2_X1 prince_inst_S_9__srx_U1 ( .A(prince_inst_rc2_inv[9]), .B(
        prince_inst_sout_x[9]), .Z(final_x[25]) );
  MUX2_X1 prince_inst_S_9__mux_inv_x1_U1 ( .A(prince_inst_srin_x[9]), .B(
        prince_inst_xout_x[9]), .S(prince_inst_n30), .Z(prince_inst_sin_x[9])
         );
  MUX2_X1 prince_inst_S_9__mux_inv_y1_U1 ( .A(prince_inst_srin_y[9]), .B(
        prince_inst_srin_y[41]), .S(prince_inst_n27), .Z(prince_inst_sin_y[9])
         );
  MUX2_X1 prince_inst_S_9__mux_inv_x2_U1 ( .A(final_x[25]), .B(
        prince_inst_sout_x[9]), .S(prince_inst_n19), .Z(prince_inst_min_x[9])
         );
  MUX2_X1 prince_inst_S_9__mux_inv_y2_U1 ( .A(final_y[25]), .B(final_y[25]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[9]) );
  XOR2_X1 prince_inst_S_10__x_U1 ( .A(rc[10]), .B(prince_inst_srin_x[42]), .Z(
        prince_inst_xout_x[10]) );
  XOR2_X1 prince_inst_S_10__srx_U1 ( .A(prince_inst_rc2_inv[10]), .B(
        prince_inst_sout_x[10]), .Z(final_x[26]) );
  MUX2_X1 prince_inst_S_10__mux_inv_x1_U1 ( .A(prince_inst_srin_x[10]), .B(
        prince_inst_xout_x[10]), .S(prince_inst_n28), .Z(prince_inst_sin_x[10]) );
  MUX2_X1 prince_inst_S_10__mux_inv_y1_U1 ( .A(prince_inst_srin_y[10]), .B(
        prince_inst_srin_y[42]), .S(prince_inst_n32), .Z(prince_inst_sin_y[10]) );
  MUX2_X1 prince_inst_S_10__mux_inv_x2_U1 ( .A(final_x[26]), .B(
        prince_inst_sout_x[10]), .S(prince_inst_n19), .Z(prince_inst_min_x[10]) );
  MUX2_X1 prince_inst_S_10__mux_inv_y2_U1 ( .A(final_y[26]), .B(final_y[26]), 
        .S(prince_inst_n22), .Z(prince_inst_min_y[10]) );
  XOR2_X1 prince_inst_S_11__x_U1 ( .A(rc[11]), .B(prince_inst_srin_x[43]), .Z(
        prince_inst_xout_x[11]) );
  XOR2_X1 prince_inst_S_11__srx_U1 ( .A(prince_inst_rc2_inv[11]), .B(
        prince_inst_sout_x[11]), .Z(final_x[27]) );
  MUX2_X1 prince_inst_S_11__mux_inv_x1_U1 ( .A(prince_inst_srin_x[11]), .B(
        prince_inst_xout_x[11]), .S(prince_inst_n31), .Z(prince_inst_sin_x[11]) );
  MUX2_X1 prince_inst_S_11__mux_inv_y1_U1 ( .A(prince_inst_srin_y[11]), .B(
        prince_inst_srin_y[43]), .S(prince_inst_n26), .Z(prince_inst_sin_y[11]) );
  MUX2_X1 prince_inst_S_11__mux_inv_x2_U1 ( .A(final_x[27]), .B(
        prince_inst_sout_x[11]), .S(prince_inst_n19), .Z(prince_inst_min_x[11]) );
  MUX2_X1 prince_inst_S_11__mux_inv_y2_U1 ( .A(final_y[27]), .B(final_y[27]), 
        .S(prince_inst_n20), .Z(prince_inst_min_y[11]) );
  XOR2_X1 prince_inst_S_12__x_U1 ( .A(rc[12]), .B(prince_inst_srin_x[12]), .Z(
        prince_inst_xout_x[12]) );
  XOR2_X1 prince_inst_S_12__srx_U1 ( .A(prince_inst_rc2_inv[12]), .B(
        prince_inst_sout_x[12]), .Z(final_x[12]) );
  MUX2_X1 prince_inst_S_12__mux_inv_x1_U1 ( .A(prince_inst_srin_x[12]), .B(
        prince_inst_xout_x[12]), .S(prince_inst_n30), .Z(prince_inst_sin_x[12]) );
  MUX2_X1 prince_inst_S_12__mux_inv_y1_U1 ( .A(prince_inst_srin_y[12]), .B(
        prince_inst_srin_y[12]), .S(prince_inst_n30), .Z(prince_inst_sin_y[12]) );
  MUX2_X1 prince_inst_S_12__mux_inv_x2_U1 ( .A(final_x[12]), .B(
        prince_inst_sout_x[12]), .S(prince_inst_n19), .Z(prince_inst_min_x[12]) );
  MUX2_X1 prince_inst_S_12__mux_inv_y2_U1 ( .A(final_y[12]), .B(final_y[12]), 
        .S(prince_inst_n21), .Z(prince_inst_min_y[12]) );
  XOR2_X1 prince_inst_S_13__x_U1 ( .A(rc[13]), .B(prince_inst_srin_x[13]), .Z(
        prince_inst_xout_x[13]) );
  XOR2_X1 prince_inst_S_13__srx_U1 ( .A(prince_inst_rc2_inv[13]), .B(
        prince_inst_sout_x[13]), .Z(final_x[13]) );
  MUX2_X1 prince_inst_S_13__mux_inv_x1_U1 ( .A(prince_inst_srin_x[13]), .B(
        prince_inst_xout_x[13]), .S(prince_inst_n32), .Z(prince_inst_sin_x[13]) );
  MUX2_X1 prince_inst_S_13__mux_inv_y1_U1 ( .A(prince_inst_srin_y[13]), .B(
        prince_inst_srin_y[13]), .S(prince_inst_n29), .Z(prince_inst_sin_y[13]) );
  MUX2_X1 prince_inst_S_13__mux_inv_x2_U1 ( .A(final_x[13]), .B(
        prince_inst_sout_x[13]), .S(prince_inst_n20), .Z(prince_inst_min_x[13]) );
  MUX2_X1 prince_inst_S_13__mux_inv_y2_U1 ( .A(final_y[13]), .B(final_y[13]), 
        .S(prince_inst_n20), .Z(prince_inst_min_y[13]) );
  XOR2_X1 prince_inst_S_14__x_U1 ( .A(rc[14]), .B(prince_inst_srin_x[14]), .Z(
        prince_inst_xout_x[14]) );
  XOR2_X1 prince_inst_S_14__srx_U1 ( .A(prince_inst_rc2_inv[14]), .B(
        prince_inst_sout_x[14]), .Z(final_x[14]) );
  MUX2_X1 prince_inst_S_14__mux_inv_x1_U1 ( .A(prince_inst_srin_x[14]), .B(
        prince_inst_xout_x[14]), .S(prince_inst_n32), .Z(prince_inst_sin_x[14]) );
  MUX2_X1 prince_inst_S_14__mux_inv_y1_U1 ( .A(prince_inst_srin_y[14]), .B(
        prince_inst_srin_y[14]), .S(prince_inst_n27), .Z(prince_inst_sin_y[14]) );
  MUX2_X1 prince_inst_S_14__mux_inv_x2_U1 ( .A(final_x[14]), .B(
        prince_inst_sout_x[14]), .S(prince_inst_n20), .Z(prince_inst_min_x[14]) );
  MUX2_X1 prince_inst_S_14__mux_inv_y2_U1 ( .A(final_y[14]), .B(final_y[14]), 
        .S(prince_inst_n21), .Z(prince_inst_min_y[14]) );
  XOR2_X1 prince_inst_S_15__x_U1 ( .A(prince_inst_rc2_inv[15]), .B(
        prince_inst_srin_x[15]), .Z(prince_inst_xout_x[15]) );
  XOR2_X1 prince_inst_S_15__srx_U1 ( .A(prince_inst_rc2_inv[15]), .B(
        prince_inst_sout_x[15]), .Z(final_x[15]) );
  MUX2_X1 prince_inst_S_15__mux_inv_x1_U1 ( .A(prince_inst_srin_x[15]), .B(
        prince_inst_xout_x[15]), .S(prince_inst_n28), .Z(prince_inst_sin_x[15]) );
  MUX2_X1 prince_inst_S_15__mux_inv_y1_U1 ( .A(prince_inst_srin_y[15]), .B(
        prince_inst_srin_y[15]), .S(prince_inst_n27), .Z(prince_inst_sin_y[15]) );
  MUX2_X1 prince_inst_S_15__mux_inv_x2_U1 ( .A(final_x[15]), .B(
        prince_inst_sout_x[15]), .S(prince_inst_n19), .Z(prince_inst_min_x[15]) );
  MUX2_X1 prince_inst_S_15__mux_inv_y2_U1 ( .A(final_y[15]), .B(final_y[15]), 
        .S(prince_inst_n19), .Z(prince_inst_min_y[15]) );
  XOR2_X1 prince_inst_S_16__x_U1 ( .A(rc[16]), .B(prince_inst_srin_x[48]), .Z(
        prince_inst_xout_x[16]) );
  XOR2_X1 prince_inst_S_16__srx_U1 ( .A(prince_inst_rc2_inv[16]), .B(
        prince_inst_sout_x[16]), .Z(final_x[0]) );
  MUX2_X1 prince_inst_S_16__mux_inv_x1_U1 ( .A(prince_inst_srin_x[16]), .B(
        prince_inst_xout_x[16]), .S(prince_inst_n31), .Z(prince_inst_sin_x[16]) );
  MUX2_X1 prince_inst_S_16__mux_inv_y1_U1 ( .A(prince_inst_srin_y[16]), .B(
        prince_inst_srin_y[48]), .S(prince_inst_n31), .Z(prince_inst_sin_y[16]) );
  MUX2_X1 prince_inst_S_16__mux_inv_x2_U1 ( .A(final_x[0]), .B(
        prince_inst_sout_x[16]), .S(prince_inst_n20), .Z(prince_inst_min_x[16]) );
  MUX2_X1 prince_inst_S_16__mux_inv_y2_U1 ( .A(final_y[0]), .B(final_y[0]), 
        .S(prince_inst_n23), .Z(prince_inst_min_y[16]) );
  XOR2_X1 prince_inst_S_17__x_U1 ( .A(rc[17]), .B(prince_inst_srin_x[49]), .Z(
        prince_inst_xout_x[17]) );
  XOR2_X1 prince_inst_S_17__srx_U1 ( .A(prince_inst_rc2_inv[17]), .B(
        prince_inst_sout_x[17]), .Z(final_x[1]) );
  MUX2_X1 prince_inst_S_17__mux_inv_x1_U1 ( .A(prince_inst_srin_x[17]), .B(
        prince_inst_xout_x[17]), .S(prince_inst_n31), .Z(prince_inst_sin_x[17]) );
  MUX2_X1 prince_inst_S_17__mux_inv_y1_U1 ( .A(prince_inst_srin_y[17]), .B(
        prince_inst_srin_y[49]), .S(prince_inst_n32), .Z(prince_inst_sin_y[17]) );
  MUX2_X1 prince_inst_S_17__mux_inv_x2_U1 ( .A(final_x[1]), .B(
        prince_inst_sout_x[17]), .S(prince_inst_n20), .Z(prince_inst_min_x[17]) );
  MUX2_X1 prince_inst_S_17__mux_inv_y2_U1 ( .A(final_y[1]), .B(final_y[1]), 
        .S(prince_inst_n20), .Z(prince_inst_min_y[17]) );
  XOR2_X1 prince_inst_S_18__x_U1 ( .A(rc[18]), .B(prince_inst_srin_x[50]), .Z(
        prince_inst_xout_x[18]) );
  XOR2_X1 prince_inst_S_18__srx_U1 ( .A(prince_inst_rc2_inv[18]), .B(
        prince_inst_sout_x[18]), .Z(final_x[2]) );
  MUX2_X1 prince_inst_S_18__mux_inv_x1_U1 ( .A(prince_inst_srin_x[18]), .B(
        prince_inst_xout_x[18]), .S(prince_inst_n32), .Z(prince_inst_sin_x[18]) );
  MUX2_X1 prince_inst_S_18__mux_inv_y1_U1 ( .A(prince_inst_srin_y[18]), .B(
        prince_inst_srin_y[50]), .S(prince_inst_n32), .Z(prince_inst_sin_y[18]) );
  MUX2_X1 prince_inst_S_18__mux_inv_x2_U1 ( .A(final_x[2]), .B(
        prince_inst_sout_x[18]), .S(prince_inst_n20), .Z(prince_inst_min_x[18]) );
  MUX2_X1 prince_inst_S_18__mux_inv_y2_U1 ( .A(final_y[2]), .B(final_y[2]), 
        .S(prince_inst_n21), .Z(prince_inst_min_y[18]) );
  XOR2_X1 prince_inst_S_19__x_U1 ( .A(rc[19]), .B(prince_inst_srin_x[51]), .Z(
        prince_inst_xout_x[19]) );
  XOR2_X1 prince_inst_S_19__srx_U1 ( .A(prince_inst_rc2_inv[19]), .B(
        prince_inst_sout_x[19]), .Z(final_x[3]) );
  MUX2_X1 prince_inst_S_19__mux_inv_x1_U1 ( .A(prince_inst_srin_x[19]), .B(
        prince_inst_xout_x[19]), .S(prince_inst_n32), .Z(prince_inst_sin_x[19]) );
  MUX2_X1 prince_inst_S_19__mux_inv_y1_U1 ( .A(prince_inst_srin_y[19]), .B(
        prince_inst_srin_y[51]), .S(prince_inst_n32), .Z(prince_inst_sin_y[19]) );
  MUX2_X1 prince_inst_S_19__mux_inv_x2_U1 ( .A(final_x[3]), .B(
        prince_inst_sout_x[19]), .S(prince_inst_n20), .Z(prince_inst_min_x[19]) );
  MUX2_X1 prince_inst_S_19__mux_inv_y2_U1 ( .A(final_y[3]), .B(final_y[3]), 
        .S(prince_inst_n22), .Z(prince_inst_min_y[19]) );
  XOR2_X1 prince_inst_S_20__x_U1 ( .A(rc[20]), .B(prince_inst_srin_x[20]), .Z(
        prince_inst_xout_x[20]) );
  XOR2_X1 prince_inst_S_20__srx_U1 ( .A(prince_inst_rc2_inv[20]), .B(
        prince_inst_sout_x[20]), .Z(final_x[52]) );
  MUX2_X1 prince_inst_S_20__mux_inv_x1_U1 ( .A(prince_inst_srin_x[20]), .B(
        prince_inst_xout_x[20]), .S(prince_inst_n32), .Z(prince_inst_sin_x[20]) );
  MUX2_X1 prince_inst_S_20__mux_inv_y1_U1 ( .A(prince_inst_srin_y[20]), .B(
        prince_inst_srin_y[20]), .S(prince_inst_n32), .Z(prince_inst_sin_y[20]) );
  MUX2_X1 prince_inst_S_20__mux_inv_x2_U1 ( .A(final_x[52]), .B(
        prince_inst_sout_x[20]), .S(prince_inst_n20), .Z(prince_inst_min_x[20]) );
  MUX2_X1 prince_inst_S_20__mux_inv_y2_U1 ( .A(final_y[52]), .B(final_y[52]), 
        .S(prince_inst_n19), .Z(prince_inst_min_y[20]) );
  XOR2_X1 prince_inst_S_21__x_U1 ( .A(rc[21]), .B(prince_inst_srin_x[21]), .Z(
        prince_inst_xout_x[21]) );
  XOR2_X1 prince_inst_S_21__srx_U1 ( .A(prince_inst_rc2_inv[21]), .B(
        prince_inst_sout_x[21]), .Z(final_x[53]) );
  MUX2_X1 prince_inst_S_21__mux_inv_x1_U1 ( .A(prince_inst_srin_x[21]), .B(
        prince_inst_xout_x[21]), .S(prince_inst_n32), .Z(prince_inst_sin_x[21]) );
  MUX2_X1 prince_inst_S_21__mux_inv_y1_U1 ( .A(prince_inst_srin_y[21]), .B(
        prince_inst_srin_y[21]), .S(prince_inst_n32), .Z(prince_inst_sin_y[21]) );
  MUX2_X1 prince_inst_S_21__mux_inv_x2_U1 ( .A(final_x[53]), .B(
        prince_inst_sout_x[21]), .S(prince_inst_n20), .Z(prince_inst_min_x[21]) );
  MUX2_X1 prince_inst_S_21__mux_inv_y2_U1 ( .A(final_y[53]), .B(final_y[53]), 
        .S(inv_sig2), .Z(prince_inst_min_y[21]) );
  XOR2_X1 prince_inst_S_22__x_U1 ( .A(rc[22]), .B(prince_inst_srin_x[22]), .Z(
        prince_inst_xout_x[22]) );
  XOR2_X1 prince_inst_S_22__srx_U1 ( .A(prince_inst_rc2_inv[22]), .B(
        prince_inst_sout_x[22]), .Z(final_x[54]) );
  MUX2_X1 prince_inst_S_22__mux_inv_x1_U1 ( .A(prince_inst_srin_x[22]), .B(
        prince_inst_xout_x[22]), .S(prince_inst_n32), .Z(prince_inst_sin_x[22]) );
  MUX2_X1 prince_inst_S_22__mux_inv_y1_U1 ( .A(prince_inst_srin_y[22]), .B(
        prince_inst_srin_y[22]), .S(prince_inst_n32), .Z(prince_inst_sin_y[22]) );
  MUX2_X1 prince_inst_S_22__mux_inv_x2_U1 ( .A(final_x[54]), .B(
        prince_inst_sout_x[22]), .S(prince_inst_n20), .Z(prince_inst_min_x[22]) );
  MUX2_X1 prince_inst_S_22__mux_inv_y2_U1 ( .A(final_y[54]), .B(final_y[54]), 
        .S(inv_sig2), .Z(prince_inst_min_y[22]) );
  XOR2_X1 prince_inst_S_23__x_U1 ( .A(rc[23]), .B(prince_inst_srin_x[23]), .Z(
        prince_inst_xout_x[23]) );
  XOR2_X1 prince_inst_S_23__srx_U1 ( .A(prince_inst_rc2_inv[23]), .B(
        prince_inst_sout_x[23]), .Z(final_x[55]) );
  MUX2_X1 prince_inst_S_23__mux_inv_x1_U1 ( .A(prince_inst_srin_x[23]), .B(
        prince_inst_xout_x[23]), .S(prince_inst_n32), .Z(prince_inst_sin_x[23]) );
  MUX2_X1 prince_inst_S_23__mux_inv_y1_U1 ( .A(prince_inst_srin_y[23]), .B(
        prince_inst_srin_y[23]), .S(prince_inst_n31), .Z(prince_inst_sin_y[23]) );
  MUX2_X1 prince_inst_S_23__mux_inv_x2_U1 ( .A(final_x[55]), .B(
        prince_inst_sout_x[23]), .S(prince_inst_n20), .Z(prince_inst_min_x[23]) );
  MUX2_X1 prince_inst_S_23__mux_inv_y2_U1 ( .A(final_y[55]), .B(final_y[55]), 
        .S(prince_inst_n21), .Z(prince_inst_min_y[23]) );
  XOR2_X1 prince_inst_S_24__x_U1 ( .A(rc[24]), .B(prince_inst_srin_x[56]), .Z(
        prince_inst_xout_x[24]) );
  XOR2_X1 prince_inst_S_24__srx_U1 ( .A(prince_inst_rc2_inv[24]), .B(
        prince_inst_sout_x[24]), .Z(final_x[40]) );
  MUX2_X1 prince_inst_S_24__mux_inv_x1_U1 ( .A(prince_inst_srin_x[24]), .B(
        prince_inst_xout_x[24]), .S(prince_inst_n31), .Z(prince_inst_sin_x[24]) );
  MUX2_X1 prince_inst_S_24__mux_inv_y1_U1 ( .A(prince_inst_srin_y[24]), .B(
        prince_inst_srin_y[56]), .S(prince_inst_n31), .Z(prince_inst_sin_y[24]) );
  MUX2_X1 prince_inst_S_24__mux_inv_x2_U1 ( .A(final_x[40]), .B(
        prince_inst_sout_x[24]), .S(prince_inst_n20), .Z(prince_inst_min_x[24]) );
  MUX2_X1 prince_inst_S_24__mux_inv_y2_U1 ( .A(final_y[40]), .B(final_y[40]), 
        .S(prince_inst_n20), .Z(prince_inst_min_y[24]) );
  XOR2_X1 prince_inst_S_25__x_U1 ( .A(rc[25]), .B(prince_inst_srin_x[57]), .Z(
        prince_inst_xout_x[25]) );
  XOR2_X1 prince_inst_S_25__srx_U1 ( .A(prince_inst_rc2_inv[25]), .B(
        prince_inst_sout_x[25]), .Z(final_x[41]) );
  MUX2_X1 prince_inst_S_25__mux_inv_x1_U1 ( .A(prince_inst_srin_x[25]), .B(
        prince_inst_xout_x[25]), .S(prince_inst_n31), .Z(prince_inst_sin_x[25]) );
  MUX2_X1 prince_inst_S_25__mux_inv_y1_U1 ( .A(prince_inst_srin_y[25]), .B(
        prince_inst_srin_y[57]), .S(prince_inst_n31), .Z(prince_inst_sin_y[25]) );
  MUX2_X1 prince_inst_S_25__mux_inv_x2_U1 ( .A(final_x[41]), .B(
        prince_inst_sout_x[25]), .S(prince_inst_n20), .Z(prince_inst_min_x[25]) );
  MUX2_X1 prince_inst_S_25__mux_inv_y2_U1 ( .A(final_y[41]), .B(final_y[41]), 
        .S(inv_sig2), .Z(prince_inst_min_y[25]) );
  XOR2_X1 prince_inst_S_26__x_U1 ( .A(rc[26]), .B(prince_inst_srin_x[58]), .Z(
        prince_inst_xout_x[26]) );
  XOR2_X1 prince_inst_S_26__srx_U1 ( .A(prince_inst_rc2_inv[26]), .B(
        prince_inst_sout_x[26]), .Z(final_x[42]) );
  MUX2_X1 prince_inst_S_26__mux_inv_x1_U1 ( .A(prince_inst_srin_x[26]), .B(
        prince_inst_xout_x[26]), .S(prince_inst_n31), .Z(prince_inst_sin_x[26]) );
  MUX2_X1 prince_inst_S_26__mux_inv_y1_U1 ( .A(prince_inst_srin_y[26]), .B(
        prince_inst_srin_y[58]), .S(prince_inst_n31), .Z(prince_inst_sin_y[26]) );
  MUX2_X1 prince_inst_S_26__mux_inv_x2_U1 ( .A(final_x[42]), .B(
        prince_inst_sout_x[26]), .S(prince_inst_n21), .Z(prince_inst_min_x[26]) );
  MUX2_X1 prince_inst_S_26__mux_inv_y2_U1 ( .A(final_y[42]), .B(final_y[42]), 
        .S(inv_sig2), .Z(prince_inst_min_y[26]) );
  XOR2_X1 prince_inst_S_27__x_U1 ( .A(rc[27]), .B(prince_inst_srin_x[59]), .Z(
        prince_inst_xout_x[27]) );
  XOR2_X1 prince_inst_S_27__srx_U1 ( .A(prince_inst_rc2_inv[27]), .B(
        prince_inst_sout_x[27]), .Z(final_x[43]) );
  MUX2_X1 prince_inst_S_27__mux_inv_x1_U1 ( .A(prince_inst_srin_x[27]), .B(
        prince_inst_xout_x[27]), .S(prince_inst_n31), .Z(prince_inst_sin_x[27]) );
  MUX2_X1 prince_inst_S_27__mux_inv_y1_U1 ( .A(prince_inst_srin_y[27]), .B(
        prince_inst_srin_y[59]), .S(prince_inst_n31), .Z(prince_inst_sin_y[27]) );
  MUX2_X1 prince_inst_S_27__mux_inv_x2_U1 ( .A(final_x[43]), .B(
        prince_inst_sout_x[27]), .S(prince_inst_n21), .Z(prince_inst_min_x[27]) );
  MUX2_X1 prince_inst_S_27__mux_inv_y2_U1 ( .A(final_y[43]), .B(final_y[43]), 
        .S(prince_inst_n19), .Z(prince_inst_min_y[27]) );
  XOR2_X1 prince_inst_S_28__x_U1 ( .A(rc[28]), .B(prince_inst_srin_x[28]), .Z(
        prince_inst_xout_x[28]) );
  XOR2_X1 prince_inst_S_28__srx_U1 ( .A(prince_inst_rc2_inv[28]), .B(
        prince_inst_sout_x[28]), .Z(final_x[28]) );
  MUX2_X1 prince_inst_S_28__mux_inv_x1_U1 ( .A(prince_inst_srin_x[28]), .B(
        prince_inst_xout_x[28]), .S(prince_inst_n31), .Z(prince_inst_sin_x[28]) );
  MUX2_X1 prince_inst_S_28__mux_inv_y1_U1 ( .A(prince_inst_srin_y[28]), .B(
        prince_inst_srin_y[28]), .S(prince_inst_n31), .Z(prince_inst_sin_y[28]) );
  MUX2_X1 prince_inst_S_28__mux_inv_x2_U1 ( .A(final_x[28]), .B(
        prince_inst_sout_x[28]), .S(prince_inst_n21), .Z(prince_inst_min_x[28]) );
  MUX2_X1 prince_inst_S_28__mux_inv_y2_U1 ( .A(final_y[28]), .B(final_y[28]), 
        .S(inv_sig2), .Z(prince_inst_min_y[28]) );
  XOR2_X1 prince_inst_S_29__x_U1 ( .A(rc[29]), .B(prince_inst_srin_x[29]), .Z(
        prince_inst_xout_x[29]) );
  XOR2_X1 prince_inst_S_29__srx_U1 ( .A(prince_inst_rc2_inv[29]), .B(
        prince_inst_sout_x[29]), .Z(final_x[29]) );
  MUX2_X1 prince_inst_S_29__mux_inv_x1_U1 ( .A(prince_inst_srin_x[29]), .B(
        prince_inst_xout_x[29]), .S(prince_inst_n31), .Z(prince_inst_sin_x[29]) );
  MUX2_X1 prince_inst_S_29__mux_inv_y1_U1 ( .A(prince_inst_srin_y[29]), .B(
        prince_inst_srin_y[29]), .S(prince_inst_n30), .Z(prince_inst_sin_y[29]) );
  MUX2_X1 prince_inst_S_29__mux_inv_x2_U1 ( .A(final_x[29]), .B(
        prince_inst_sout_x[29]), .S(prince_inst_n21), .Z(prince_inst_min_x[29]) );
  MUX2_X1 prince_inst_S_29__mux_inv_y2_U1 ( .A(final_y[29]), .B(final_y[29]), 
        .S(inv_sig2), .Z(prince_inst_min_y[29]) );
  XOR2_X1 prince_inst_S_30__x_U1 ( .A(rc[30]), .B(prince_inst_srin_x[30]), .Z(
        prince_inst_xout_x[30]) );
  XOR2_X1 prince_inst_S_30__srx_U1 ( .A(prince_inst_rc2_inv[30]), .B(
        prince_inst_sout_x[30]), .Z(final_x[30]) );
  MUX2_X1 prince_inst_S_30__mux_inv_x1_U1 ( .A(prince_inst_srin_x[30]), .B(
        prince_inst_xout_x[30]), .S(prince_inst_n30), .Z(prince_inst_sin_x[30]) );
  MUX2_X1 prince_inst_S_30__mux_inv_y1_U1 ( .A(prince_inst_srin_y[30]), .B(
        prince_inst_srin_y[30]), .S(prince_inst_n30), .Z(prince_inst_sin_y[30]) );
  MUX2_X1 prince_inst_S_30__mux_inv_x2_U1 ( .A(final_x[30]), .B(
        prince_inst_sout_x[30]), .S(prince_inst_n21), .Z(prince_inst_min_x[30]) );
  MUX2_X1 prince_inst_S_30__mux_inv_y2_U1 ( .A(final_y[30]), .B(final_y[30]), 
        .S(inv_sig2), .Z(prince_inst_min_y[30]) );
  XOR2_X1 prince_inst_S_31__x_U1 ( .A(rc[31]), .B(prince_inst_srin_x[31]), .Z(
        prince_inst_xout_x[31]) );
  XOR2_X1 prince_inst_S_31__srx_U1 ( .A(prince_inst_rc2_inv[31]), .B(
        prince_inst_sout_x[31]), .Z(final_x[31]) );
  MUX2_X1 prince_inst_S_31__mux_inv_x1_U1 ( .A(prince_inst_srin_x[31]), .B(
        prince_inst_xout_x[31]), .S(prince_inst_n30), .Z(prince_inst_sin_x[31]) );
  MUX2_X1 prince_inst_S_31__mux_inv_y1_U1 ( .A(prince_inst_srin_y[31]), .B(
        prince_inst_srin_y[31]), .S(prince_inst_n30), .Z(prince_inst_sin_y[31]) );
  MUX2_X1 prince_inst_S_31__mux_inv_x2_U1 ( .A(final_x[31]), .B(
        prince_inst_sout_x[31]), .S(prince_inst_n21), .Z(prince_inst_min_x[31]) );
  MUX2_X1 prince_inst_S_31__mux_inv_y2_U1 ( .A(final_y[31]), .B(final_y[31]), 
        .S(prince_inst_n23), .Z(prince_inst_min_y[31]) );
  XOR2_X1 prince_inst_S_32__x_U1 ( .A(rc[32]), .B(prince_inst_srin_x[0]), .Z(
        prince_inst_xout_x[32]) );
  XOR2_X1 prince_inst_S_32__srx_U1 ( .A(prince_inst_rc2_inv[32]), .B(
        prince_inst_sout_x[32]), .Z(final_x[16]) );
  MUX2_X1 prince_inst_S_32__mux_inv_x1_U1 ( .A(prince_inst_srin_x[32]), .B(
        prince_inst_xout_x[32]), .S(prince_inst_n30), .Z(prince_inst_sin_x[32]) );
  MUX2_X1 prince_inst_S_32__mux_inv_y1_U1 ( .A(prince_inst_srin_y[32]), .B(
        prince_inst_srin_y[0]), .S(prince_inst_n30), .Z(prince_inst_sin_y[32])
         );
  MUX2_X1 prince_inst_S_32__mux_inv_x2_U1 ( .A(final_x[16]), .B(
        prince_inst_sout_x[32]), .S(prince_inst_n21), .Z(prince_inst_min_x[32]) );
  MUX2_X1 prince_inst_S_32__mux_inv_y2_U1 ( .A(final_y[16]), .B(final_y[16]), 
        .S(prince_inst_n21), .Z(prince_inst_min_y[32]) );
  XOR2_X1 prince_inst_S_33__x_U1 ( .A(rc[33]), .B(prince_inst_srin_x[1]), .Z(
        prince_inst_xout_x[33]) );
  XOR2_X1 prince_inst_S_33__srx_U1 ( .A(prince_inst_rc2_inv[33]), .B(
        prince_inst_sout_x[33]), .Z(final_x[17]) );
  MUX2_X1 prince_inst_S_33__mux_inv_x1_U1 ( .A(prince_inst_srin_x[33]), .B(
        prince_inst_xout_x[33]), .S(prince_inst_n30), .Z(prince_inst_sin_x[33]) );
  MUX2_X1 prince_inst_S_33__mux_inv_y1_U1 ( .A(prince_inst_srin_y[33]), .B(
        prince_inst_srin_y[1]), .S(prince_inst_n30), .Z(prince_inst_sin_y[33])
         );
  MUX2_X1 prince_inst_S_33__mux_inv_x2_U1 ( .A(final_x[17]), .B(
        prince_inst_sout_x[33]), .S(prince_inst_n21), .Z(prince_inst_min_x[33]) );
  MUX2_X1 prince_inst_S_33__mux_inv_y2_U1 ( .A(final_y[17]), .B(final_y[17]), 
        .S(inv_sig2), .Z(prince_inst_min_y[33]) );
  XOR2_X1 prince_inst_S_34__x_U1 ( .A(rc[34]), .B(prince_inst_srin_x[2]), .Z(
        prince_inst_xout_x[34]) );
  XOR2_X1 prince_inst_S_34__srx_U1 ( .A(prince_inst_rc2_inv[34]), .B(
        prince_inst_sout_x[34]), .Z(final_x[18]) );
  MUX2_X1 prince_inst_S_34__mux_inv_x1_U1 ( .A(prince_inst_srin_x[34]), .B(
        prince_inst_xout_x[34]), .S(prince_inst_n30), .Z(prince_inst_sin_x[34]) );
  MUX2_X1 prince_inst_S_34__mux_inv_y1_U1 ( .A(prince_inst_srin_y[34]), .B(
        prince_inst_srin_y[2]), .S(prince_inst_n30), .Z(prince_inst_sin_y[34])
         );
  MUX2_X1 prince_inst_S_34__mux_inv_x2_U1 ( .A(final_x[18]), .B(
        prince_inst_sout_x[34]), .S(prince_inst_n21), .Z(prince_inst_min_x[34]) );
  MUX2_X1 prince_inst_S_34__mux_inv_y2_U1 ( .A(final_y[18]), .B(final_y[18]), 
        .S(prince_inst_n23), .Z(prince_inst_min_y[34]) );
  XOR2_X1 prince_inst_S_35__x_U1 ( .A(rc[35]), .B(prince_inst_srin_x[3]), .Z(
        prince_inst_xout_x[35]) );
  XOR2_X1 prince_inst_S_35__srx_U1 ( .A(prince_inst_rc2_inv[35]), .B(
        prince_inst_sout_x[35]), .Z(final_x[19]) );
  MUX2_X1 prince_inst_S_35__mux_inv_x1_U1 ( .A(prince_inst_srin_x[35]), .B(
        prince_inst_xout_x[35]), .S(prince_inst_n29), .Z(prince_inst_sin_x[35]) );
  MUX2_X1 prince_inst_S_35__mux_inv_y1_U1 ( .A(prince_inst_srin_y[35]), .B(
        prince_inst_srin_y[3]), .S(prince_inst_n29), .Z(prince_inst_sin_y[35])
         );
  MUX2_X1 prince_inst_S_35__mux_inv_x2_U1 ( .A(final_x[19]), .B(
        prince_inst_sout_x[35]), .S(prince_inst_n21), .Z(prince_inst_min_x[35]) );
  MUX2_X1 prince_inst_S_35__mux_inv_y2_U1 ( .A(final_y[19]), .B(final_y[19]), 
        .S(prince_inst_n22), .Z(prince_inst_min_y[35]) );
  XOR2_X1 prince_inst_S_36__x_U1 ( .A(rc[36]), .B(prince_inst_srin_x[36]), .Z(
        prince_inst_xout_x[36]) );
  XOR2_X1 prince_inst_S_36__srx_U1 ( .A(prince_inst_rc2_inv[36]), .B(
        prince_inst_sout_x[36]), .Z(final_x[4]) );
  MUX2_X1 prince_inst_S_36__mux_inv_x1_U1 ( .A(prince_inst_srin_x[36]), .B(
        prince_inst_xout_x[36]), .S(prince_inst_n29), .Z(prince_inst_sin_x[36]) );
  MUX2_X1 prince_inst_S_36__mux_inv_y1_U1 ( .A(prince_inst_srin_y[36]), .B(
        prince_inst_srin_y[36]), .S(prince_inst_n29), .Z(prince_inst_sin_y[36]) );
  MUX2_X1 prince_inst_S_36__mux_inv_x2_U1 ( .A(final_x[4]), .B(
        prince_inst_sout_x[36]), .S(prince_inst_n21), .Z(prince_inst_min_x[36]) );
  MUX2_X1 prince_inst_S_36__mux_inv_y2_U1 ( .A(final_y[4]), .B(final_y[4]), 
        .S(prince_inst_n22), .Z(prince_inst_min_y[36]) );
  XOR2_X1 prince_inst_S_37__x_U1 ( .A(rc[37]), .B(prince_inst_srin_x[37]), .Z(
        prince_inst_xout_x[37]) );
  XOR2_X1 prince_inst_S_37__srx_U1 ( .A(prince_inst_rc2_inv[37]), .B(
        prince_inst_sout_x[37]), .Z(final_x[5]) );
  MUX2_X1 prince_inst_S_37__mux_inv_x1_U1 ( .A(prince_inst_srin_x[37]), .B(
        prince_inst_xout_x[37]), .S(prince_inst_n29), .Z(prince_inst_sin_x[37]) );
  MUX2_X1 prince_inst_S_37__mux_inv_y1_U1 ( .A(prince_inst_srin_y[37]), .B(
        prince_inst_srin_y[37]), .S(prince_inst_n29), .Z(prince_inst_sin_y[37]) );
  MUX2_X1 prince_inst_S_37__mux_inv_x2_U1 ( .A(final_x[5]), .B(
        prince_inst_sout_x[37]), .S(prince_inst_n21), .Z(prince_inst_min_x[37]) );
  MUX2_X1 prince_inst_S_37__mux_inv_y2_U1 ( .A(final_y[5]), .B(final_y[5]), 
        .S(inv_sig2), .Z(prince_inst_min_y[37]) );
  XOR2_X1 prince_inst_S_38__x_U1 ( .A(rc[38]), .B(prince_inst_srin_x[38]), .Z(
        prince_inst_xout_x[38]) );
  XOR2_X1 prince_inst_S_38__srx_U1 ( .A(prince_inst_rc2_inv[38]), .B(
        prince_inst_sout_x[38]), .Z(final_x[6]) );
  MUX2_X1 prince_inst_S_38__mux_inv_x1_U1 ( .A(prince_inst_srin_x[38]), .B(
        prince_inst_xout_x[38]), .S(prince_inst_n29), .Z(prince_inst_sin_x[38]) );
  MUX2_X1 prince_inst_S_38__mux_inv_y1_U1 ( .A(prince_inst_srin_y[38]), .B(
        prince_inst_srin_y[38]), .S(prince_inst_n29), .Z(prince_inst_sin_y[38]) );
  MUX2_X1 prince_inst_S_38__mux_inv_x2_U1 ( .A(final_x[6]), .B(
        prince_inst_sout_x[38]), .S(prince_inst_n22), .Z(prince_inst_min_x[38]) );
  MUX2_X1 prince_inst_S_38__mux_inv_y2_U1 ( .A(final_y[6]), .B(final_y[6]), 
        .S(inv_sig2), .Z(prince_inst_min_y[38]) );
  XOR2_X1 prince_inst_S_39__x_U1 ( .A(rc[39]), .B(prince_inst_srin_x[39]), .Z(
        prince_inst_xout_x[39]) );
  XOR2_X1 prince_inst_S_39__srx_U1 ( .A(prince_inst_rc2_inv[39]), .B(
        prince_inst_sout_x[39]), .Z(final_x[7]) );
  MUX2_X1 prince_inst_S_39__mux_inv_x1_U1 ( .A(prince_inst_srin_x[39]), .B(
        prince_inst_xout_x[39]), .S(prince_inst_n29), .Z(prince_inst_sin_x[39]) );
  MUX2_X1 prince_inst_S_39__mux_inv_y1_U1 ( .A(prince_inst_srin_y[39]), .B(
        prince_inst_srin_y[39]), .S(prince_inst_n29), .Z(prince_inst_sin_y[39]) );
  MUX2_X1 prince_inst_S_39__mux_inv_x2_U1 ( .A(final_x[7]), .B(
        prince_inst_sout_x[39]), .S(prince_inst_n22), .Z(prince_inst_min_x[39]) );
  MUX2_X1 prince_inst_S_39__mux_inv_y2_U1 ( .A(final_y[7]), .B(final_y[7]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[39]) );
  XOR2_X1 prince_inst_S_40__x_U1 ( .A(rc[40]), .B(prince_inst_srin_x[8]), .Z(
        prince_inst_xout_x[40]) );
  XOR2_X1 prince_inst_S_40__srx_U1 ( .A(prince_inst_rc2_inv[40]), .B(
        prince_inst_sout_x[40]), .Z(final_x[56]) );
  MUX2_X1 prince_inst_S_40__mux_inv_x1_U1 ( .A(prince_inst_srin_x[40]), .B(
        prince_inst_xout_x[40]), .S(prince_inst_n29), .Z(prince_inst_sin_x[40]) );
  MUX2_X1 prince_inst_S_40__mux_inv_y1_U1 ( .A(prince_inst_srin_y[40]), .B(
        prince_inst_srin_y[8]), .S(prince_inst_n29), .Z(prince_inst_sin_y[40])
         );
  MUX2_X1 prince_inst_S_40__mux_inv_x2_U1 ( .A(final_x[56]), .B(
        prince_inst_sout_x[40]), .S(prince_inst_n22), .Z(prince_inst_min_x[40]) );
  MUX2_X1 prince_inst_S_40__mux_inv_y2_U1 ( .A(final_y[56]), .B(final_y[56]), 
        .S(prince_inst_n22), .Z(prince_inst_min_y[40]) );
  XOR2_X1 prince_inst_S_41__x_U1 ( .A(rc[41]), .B(prince_inst_srin_x[9]), .Z(
        prince_inst_xout_x[41]) );
  XOR2_X1 prince_inst_S_41__srx_U1 ( .A(prince_inst_rc2_inv[41]), .B(
        prince_inst_sout_x[41]), .Z(final_x[57]) );
  MUX2_X1 prince_inst_S_41__mux_inv_x1_U1 ( .A(prince_inst_srin_x[41]), .B(
        prince_inst_xout_x[41]), .S(prince_inst_n28), .Z(prince_inst_sin_x[41]) );
  MUX2_X1 prince_inst_S_41__mux_inv_y1_U1 ( .A(prince_inst_srin_y[41]), .B(
        prince_inst_srin_y[9]), .S(prince_inst_n28), .Z(prince_inst_sin_y[41])
         );
  MUX2_X1 prince_inst_S_41__mux_inv_x2_U1 ( .A(final_x[57]), .B(
        prince_inst_sout_x[41]), .S(prince_inst_n22), .Z(prince_inst_min_x[41]) );
  MUX2_X1 prince_inst_S_41__mux_inv_y2_U1 ( .A(final_y[57]), .B(final_y[57]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[41]) );
  XOR2_X1 prince_inst_S_42__x_U1 ( .A(rc[42]), .B(prince_inst_srin_x[10]), .Z(
        prince_inst_xout_x[42]) );
  XOR2_X1 prince_inst_S_42__srx_U1 ( .A(prince_inst_rc2_inv[42]), .B(
        prince_inst_sout_x[42]), .Z(final_x[58]) );
  MUX2_X1 prince_inst_S_42__mux_inv_x1_U1 ( .A(prince_inst_srin_x[42]), .B(
        prince_inst_xout_x[42]), .S(prince_inst_n28), .Z(prince_inst_sin_x[42]) );
  MUX2_X1 prince_inst_S_42__mux_inv_y1_U1 ( .A(prince_inst_srin_y[42]), .B(
        prince_inst_srin_y[10]), .S(prince_inst_n28), .Z(prince_inst_sin_y[42]) );
  MUX2_X1 prince_inst_S_42__mux_inv_x2_U1 ( .A(final_x[58]), .B(
        prince_inst_sout_x[42]), .S(prince_inst_n22), .Z(prince_inst_min_x[42]) );
  MUX2_X1 prince_inst_S_42__mux_inv_y2_U1 ( .A(final_y[58]), .B(final_y[58]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[42]) );
  XOR2_X1 prince_inst_S_43__x_U1 ( .A(rc[43]), .B(prince_inst_srin_x[11]), .Z(
        prince_inst_xout_x[43]) );
  XOR2_X1 prince_inst_S_43__srx_U1 ( .A(prince_inst_rc2_inv[43]), .B(
        prince_inst_sout_x[43]), .Z(final_x[59]) );
  MUX2_X1 prince_inst_S_43__mux_inv_x1_U1 ( .A(prince_inst_srin_x[43]), .B(
        prince_inst_xout_x[43]), .S(prince_inst_n28), .Z(prince_inst_sin_x[43]) );
  MUX2_X1 prince_inst_S_43__mux_inv_y1_U1 ( .A(prince_inst_srin_y[43]), .B(
        prince_inst_srin_y[11]), .S(prince_inst_n28), .Z(prince_inst_sin_y[43]) );
  MUX2_X1 prince_inst_S_43__mux_inv_x2_U1 ( .A(final_x[59]), .B(
        prince_inst_sout_x[43]), .S(prince_inst_n22), .Z(prince_inst_min_x[43]) );
  MUX2_X1 prince_inst_S_43__mux_inv_y2_U1 ( .A(final_y[59]), .B(final_y[59]), 
        .S(inv_sig2), .Z(prince_inst_min_y[43]) );
  XOR2_X1 prince_inst_S_44__x_U1 ( .A(rc[44]), .B(prince_inst_srin_x[44]), .Z(
        prince_inst_xout_x[44]) );
  XOR2_X1 prince_inst_S_44__srx_U1 ( .A(prince_inst_rc2_inv[44]), .B(
        prince_inst_sout_x[44]), .Z(final_x[44]) );
  MUX2_X1 prince_inst_S_44__mux_inv_x1_U1 ( .A(prince_inst_srin_x[44]), .B(
        prince_inst_xout_x[44]), .S(prince_inst_n28), .Z(prince_inst_sin_x[44]) );
  MUX2_X1 prince_inst_S_44__mux_inv_y1_U1 ( .A(prince_inst_srin_y[44]), .B(
        prince_inst_srin_y[44]), .S(prince_inst_n28), .Z(prince_inst_sin_y[44]) );
  MUX2_X1 prince_inst_S_44__mux_inv_x2_U1 ( .A(final_x[44]), .B(
        prince_inst_sout_x[44]), .S(prince_inst_n22), .Z(prince_inst_min_x[44]) );
  MUX2_X1 prince_inst_S_44__mux_inv_y2_U1 ( .A(final_y[44]), .B(final_y[44]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[44]) );
  XOR2_X1 prince_inst_S_45__x_U1 ( .A(rc[45]), .B(prince_inst_srin_x[45]), .Z(
        prince_inst_xout_x[45]) );
  XOR2_X1 prince_inst_S_45__srx_U1 ( .A(prince_inst_rc2_inv[45]), .B(
        prince_inst_sout_x[45]), .Z(final_x[45]) );
  MUX2_X1 prince_inst_S_45__mux_inv_x1_U1 ( .A(prince_inst_srin_x[45]), .B(
        prince_inst_xout_x[45]), .S(prince_inst_n28), .Z(prince_inst_sin_x[45]) );
  MUX2_X1 prince_inst_S_45__mux_inv_y1_U1 ( .A(prince_inst_srin_y[45]), .B(
        prince_inst_srin_y[45]), .S(prince_inst_n28), .Z(prince_inst_sin_y[45]) );
  MUX2_X1 prince_inst_S_45__mux_inv_x2_U1 ( .A(final_x[45]), .B(
        prince_inst_sout_x[45]), .S(prince_inst_n22), .Z(prince_inst_min_x[45]) );
  MUX2_X1 prince_inst_S_45__mux_inv_y2_U1 ( .A(final_y[45]), .B(final_y[45]), 
        .S(prince_inst_n19), .Z(prince_inst_min_y[45]) );
  XOR2_X1 prince_inst_S_46__x_U1 ( .A(rc[46]), .B(prince_inst_srin_x[46]), .Z(
        prince_inst_xout_x[46]) );
  XOR2_X1 prince_inst_S_46__srx_U1 ( .A(prince_inst_rc2_inv[46]), .B(
        prince_inst_sout_x[46]), .Z(final_x[46]) );
  MUX2_X1 prince_inst_S_46__mux_inv_x1_U1 ( .A(prince_inst_srin_x[46]), .B(
        prince_inst_xout_x[46]), .S(prince_inst_n28), .Z(prince_inst_sin_x[46]) );
  MUX2_X1 prince_inst_S_46__mux_inv_y1_U1 ( .A(prince_inst_srin_y[46]), .B(
        prince_inst_srin_y[46]), .S(prince_inst_n28), .Z(prince_inst_sin_y[46]) );
  MUX2_X1 prince_inst_S_46__mux_inv_x2_U1 ( .A(final_x[46]), .B(
        prince_inst_sout_x[46]), .S(prince_inst_n22), .Z(prince_inst_min_x[46]) );
  MUX2_X1 prince_inst_S_46__mux_inv_y2_U1 ( .A(final_y[46]), .B(final_y[46]), 
        .S(prince_inst_n20), .Z(prince_inst_min_y[46]) );
  XOR2_X1 prince_inst_S_47__x_U1 ( .A(rc[47]), .B(prince_inst_srin_x[47]), .Z(
        prince_inst_xout_x[47]) );
  XOR2_X1 prince_inst_S_47__srx_U1 ( .A(prince_inst_rc2_inv[47]), .B(
        prince_inst_sout_x[47]), .Z(final_x[47]) );
  MUX2_X1 prince_inst_S_47__mux_inv_x1_U1 ( .A(prince_inst_srin_x[47]), .B(
        prince_inst_xout_x[47]), .S(prince_inst_n27), .Z(prince_inst_sin_x[47]) );
  MUX2_X1 prince_inst_S_47__mux_inv_y1_U1 ( .A(prince_inst_srin_y[47]), .B(
        prince_inst_srin_y[47]), .S(prince_inst_n27), .Z(prince_inst_sin_y[47]) );
  MUX2_X1 prince_inst_S_47__mux_inv_x2_U1 ( .A(final_x[47]), .B(
        prince_inst_sout_x[47]), .S(prince_inst_n22), .Z(prince_inst_min_x[47]) );
  MUX2_X1 prince_inst_S_47__mux_inv_y2_U1 ( .A(final_y[47]), .B(final_y[47]), 
        .S(inv_sig2), .Z(prince_inst_min_y[47]) );
  XOR2_X1 prince_inst_S_48__x_U1 ( .A(rc[48]), .B(prince_inst_srin_x[16]), .Z(
        prince_inst_xout_x[48]) );
  XOR2_X1 prince_inst_S_48__srx_U1 ( .A(prince_inst_rc2_inv[48]), .B(
        prince_inst_sout_x[48]), .Z(final_x[32]) );
  MUX2_X1 prince_inst_S_48__mux_inv_x1_U1 ( .A(prince_inst_srin_x[48]), .B(
        prince_inst_xout_x[48]), .S(prince_inst_n27), .Z(prince_inst_sin_x[48]) );
  MUX2_X1 prince_inst_S_48__mux_inv_y1_U1 ( .A(prince_inst_srin_y[48]), .B(
        prince_inst_srin_y[16]), .S(prince_inst_n27), .Z(prince_inst_sin_y[48]) );
  MUX2_X1 prince_inst_S_48__mux_inv_x2_U1 ( .A(final_x[32]), .B(
        prince_inst_sout_x[48]), .S(prince_inst_n22), .Z(prince_inst_min_x[48]) );
  MUX2_X1 prince_inst_S_48__mux_inv_y2_U1 ( .A(final_y[32]), .B(final_y[32]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[48]) );
  XOR2_X1 prince_inst_S_49__x_U1 ( .A(rc[49]), .B(prince_inst_srin_x[17]), .Z(
        prince_inst_xout_x[49]) );
  XOR2_X1 prince_inst_S_49__srx_U1 ( .A(prince_inst_rc2_inv[49]), .B(
        prince_inst_sout_x[49]), .Z(final_x[33]) );
  MUX2_X1 prince_inst_S_49__mux_inv_x1_U1 ( .A(prince_inst_srin_x[49]), .B(
        prince_inst_xout_x[49]), .S(prince_inst_n27), .Z(prince_inst_sin_x[49]) );
  MUX2_X1 prince_inst_S_49__mux_inv_y1_U1 ( .A(prince_inst_srin_y[49]), .B(
        prince_inst_srin_y[17]), .S(prince_inst_n27), .Z(prince_inst_sin_y[49]) );
  MUX2_X1 prince_inst_S_49__mux_inv_x2_U1 ( .A(final_x[33]), .B(
        prince_inst_sout_x[49]), .S(prince_inst_n22), .Z(prince_inst_min_x[49]) );
  MUX2_X1 prince_inst_S_49__mux_inv_y2_U1 ( .A(final_y[33]), .B(final_y[33]), 
        .S(prince_inst_n19), .Z(prince_inst_min_y[49]) );
  XOR2_X1 prince_inst_S_50__x_U1 ( .A(rc[50]), .B(prince_inst_srin_x[18]), .Z(
        prince_inst_xout_x[50]) );
  XOR2_X1 prince_inst_S_50__srx_U1 ( .A(prince_inst_rc2_inv[50]), .B(
        prince_inst_sout_x[50]), .Z(final_x[34]) );
  MUX2_X1 prince_inst_S_50__mux_inv_x1_U1 ( .A(prince_inst_srin_x[50]), .B(
        prince_inst_xout_x[50]), .S(prince_inst_n27), .Z(prince_inst_sin_x[50]) );
  MUX2_X1 prince_inst_S_50__mux_inv_y1_U1 ( .A(prince_inst_srin_y[50]), .B(
        prince_inst_srin_y[18]), .S(prince_inst_n27), .Z(prince_inst_sin_y[50]) );
  MUX2_X1 prince_inst_S_50__mux_inv_x2_U1 ( .A(final_x[34]), .B(
        prince_inst_sout_x[50]), .S(prince_inst_n23), .Z(prince_inst_min_x[50]) );
  MUX2_X1 prince_inst_S_50__mux_inv_y2_U1 ( .A(final_y[34]), .B(final_y[34]), 
        .S(prince_inst_n22), .Z(prince_inst_min_y[50]) );
  XOR2_X1 prince_inst_S_51__x_U1 ( .A(rc[51]), .B(prince_inst_srin_x[19]), .Z(
        prince_inst_xout_x[51]) );
  XOR2_X1 prince_inst_S_51__srx_U1 ( .A(prince_inst_rc2_inv[51]), .B(
        prince_inst_sout_x[51]), .Z(final_x[35]) );
  MUX2_X1 prince_inst_S_51__mux_inv_x1_U1 ( .A(prince_inst_srin_x[51]), .B(
        prince_inst_xout_x[51]), .S(prince_inst_n27), .Z(prince_inst_sin_x[51]) );
  MUX2_X1 prince_inst_S_51__mux_inv_y1_U1 ( .A(prince_inst_srin_y[51]), .B(
        prince_inst_srin_y[19]), .S(prince_inst_n27), .Z(prince_inst_sin_y[51]) );
  MUX2_X1 prince_inst_S_51__mux_inv_x2_U1 ( .A(final_x[35]), .B(
        prince_inst_sout_x[51]), .S(prince_inst_n23), .Z(prince_inst_min_x[51]) );
  MUX2_X1 prince_inst_S_51__mux_inv_y2_U1 ( .A(final_y[35]), .B(final_y[35]), 
        .S(inv_sig2), .Z(prince_inst_min_y[51]) );
  XOR2_X1 prince_inst_S_52__x_U1 ( .A(rc[52]), .B(prince_inst_srin_x[52]), .Z(
        prince_inst_xout_x[52]) );
  XOR2_X1 prince_inst_S_52__srx_U1 ( .A(prince_inst_rc2_inv[52]), .B(
        prince_inst_sout_x[52]), .Z(final_x[20]) );
  MUX2_X1 prince_inst_S_52__mux_inv_x1_U1 ( .A(prince_inst_srin_x[52]), .B(
        prince_inst_xout_x[52]), .S(prince_inst_n27), .Z(prince_inst_sin_x[52]) );
  MUX2_X1 prince_inst_S_52__mux_inv_y1_U1 ( .A(prince_inst_srin_y[52]), .B(
        prince_inst_srin_y[52]), .S(prince_inst_n27), .Z(prince_inst_sin_y[52]) );
  MUX2_X1 prince_inst_S_52__mux_inv_x2_U1 ( .A(final_x[20]), .B(
        prince_inst_sout_x[52]), .S(prince_inst_n23), .Z(prince_inst_min_x[52]) );
  MUX2_X1 prince_inst_S_52__mux_inv_y2_U1 ( .A(final_y[20]), .B(final_y[20]), 
        .S(inv_sig2), .Z(prince_inst_min_y[52]) );
  XOR2_X1 prince_inst_S_53__x_U1 ( .A(rc[53]), .B(prince_inst_srin_x[53]), .Z(
        prince_inst_xout_x[53]) );
  XOR2_X1 prince_inst_S_53__srx_U1 ( .A(prince_inst_rc2_inv[53]), .B(
        prince_inst_sout_x[53]), .Z(final_x[21]) );
  MUX2_X1 prince_inst_S_53__mux_inv_x1_U1 ( .A(prince_inst_srin_x[53]), .B(
        prince_inst_xout_x[53]), .S(prince_inst_n26), .Z(prince_inst_sin_x[53]) );
  MUX2_X1 prince_inst_S_53__mux_inv_y1_U1 ( .A(prince_inst_srin_y[53]), .B(
        prince_inst_srin_y[53]), .S(prince_inst_n26), .Z(prince_inst_sin_y[53]) );
  MUX2_X1 prince_inst_S_53__mux_inv_x2_U1 ( .A(final_x[21]), .B(
        prince_inst_sout_x[53]), .S(prince_inst_n23), .Z(prince_inst_min_x[53]) );
  MUX2_X1 prince_inst_S_53__mux_inv_y2_U1 ( .A(final_y[21]), .B(final_y[21]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[53]) );
  XOR2_X1 prince_inst_S_54__x_U1 ( .A(rc[54]), .B(prince_inst_srin_x[54]), .Z(
        prince_inst_xout_x[54]) );
  XOR2_X1 prince_inst_S_54__srx_U1 ( .A(prince_inst_rc2_inv[54]), .B(
        prince_inst_sout_x[54]), .Z(final_x[22]) );
  MUX2_X1 prince_inst_S_54__mux_inv_x1_U1 ( .A(prince_inst_srin_x[54]), .B(
        prince_inst_xout_x[54]), .S(prince_inst_n26), .Z(prince_inst_sin_x[54]) );
  MUX2_X1 prince_inst_S_54__mux_inv_y1_U1 ( .A(prince_inst_srin_y[54]), .B(
        prince_inst_srin_y[54]), .S(prince_inst_n26), .Z(prince_inst_sin_y[54]) );
  MUX2_X1 prince_inst_S_54__mux_inv_x2_U1 ( .A(final_x[22]), .B(
        prince_inst_sout_x[54]), .S(prince_inst_n23), .Z(prince_inst_min_x[54]) );
  MUX2_X1 prince_inst_S_54__mux_inv_y2_U1 ( .A(final_y[22]), .B(final_y[22]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[54]) );
  XOR2_X1 prince_inst_S_55__x_U1 ( .A(rc[55]), .B(prince_inst_srin_x[55]), .Z(
        prince_inst_xout_x[55]) );
  XOR2_X1 prince_inst_S_55__srx_U1 ( .A(prince_inst_rc2_inv[55]), .B(
        prince_inst_sout_x[55]), .Z(final_x[23]) );
  MUX2_X1 prince_inst_S_55__mux_inv_x1_U1 ( .A(prince_inst_srin_x[55]), .B(
        prince_inst_xout_x[55]), .S(prince_inst_n26), .Z(prince_inst_sin_x[55]) );
  MUX2_X1 prince_inst_S_55__mux_inv_y1_U1 ( .A(prince_inst_srin_y[55]), .B(
        prince_inst_srin_y[55]), .S(prince_inst_n26), .Z(prince_inst_sin_y[55]) );
  MUX2_X1 prince_inst_S_55__mux_inv_x2_U1 ( .A(final_x[23]), .B(
        prince_inst_sout_x[55]), .S(prince_inst_n23), .Z(prince_inst_min_x[55]) );
  MUX2_X1 prince_inst_S_55__mux_inv_y2_U1 ( .A(final_y[23]), .B(final_y[23]), 
        .S(inv_sig2), .Z(prince_inst_min_y[55]) );
  XOR2_X1 prince_inst_S_56__x_U1 ( .A(rc[56]), .B(prince_inst_srin_x[24]), .Z(
        prince_inst_xout_x[56]) );
  XOR2_X1 prince_inst_S_56__srx_U1 ( .A(prince_inst_rc2_inv[56]), .B(
        prince_inst_sout_x[56]), .Z(final_x[8]) );
  MUX2_X1 prince_inst_S_56__mux_inv_x1_U1 ( .A(prince_inst_srin_x[56]), .B(
        prince_inst_xout_x[56]), .S(prince_inst_n26), .Z(prince_inst_sin_x[56]) );
  MUX2_X1 prince_inst_S_56__mux_inv_y1_U1 ( .A(prince_inst_srin_y[56]), .B(
        prince_inst_srin_y[24]), .S(prince_inst_n26), .Z(prince_inst_sin_y[56]) );
  MUX2_X1 prince_inst_S_56__mux_inv_x2_U1 ( .A(final_x[8]), .B(
        prince_inst_sout_x[56]), .S(prince_inst_n23), .Z(prince_inst_min_x[56]) );
  MUX2_X1 prince_inst_S_56__mux_inv_y2_U1 ( .A(final_y[8]), .B(final_y[8]), 
        .S(prince_inst_n23), .Z(prince_inst_min_y[56]) );
  XOR2_X1 prince_inst_S_57__x_U1 ( .A(rc[57]), .B(prince_inst_srin_x[25]), .Z(
        prince_inst_xout_x[57]) );
  XOR2_X1 prince_inst_S_57__srx_U1 ( .A(prince_inst_rc2_inv[57]), .B(
        prince_inst_sout_x[57]), .Z(final_x[9]) );
  MUX2_X1 prince_inst_S_57__mux_inv_x1_U1 ( .A(prince_inst_srin_x[57]), .B(
        prince_inst_xout_x[57]), .S(prince_inst_n26), .Z(prince_inst_sin_x[57]) );
  MUX2_X1 prince_inst_S_57__mux_inv_y1_U1 ( .A(prince_inst_srin_y[57]), .B(
        prince_inst_srin_y[25]), .S(prince_inst_n26), .Z(prince_inst_sin_y[57]) );
  MUX2_X1 prince_inst_S_57__mux_inv_x2_U1 ( .A(final_x[9]), .B(
        prince_inst_sout_x[57]), .S(prince_inst_n23), .Z(prince_inst_min_x[57]) );
  MUX2_X1 prince_inst_S_57__mux_inv_y2_U1 ( .A(final_y[9]), .B(final_y[9]), 
        .S(inv_sig2), .Z(prince_inst_min_y[57]) );
  XOR2_X1 prince_inst_S_58__x_U1 ( .A(rc[58]), .B(prince_inst_srin_x[26]), .Z(
        prince_inst_xout_x[58]) );
  XOR2_X1 prince_inst_S_58__srx_U1 ( .A(prince_inst_rc2_inv[58]), .B(
        prince_inst_sout_x[58]), .Z(final_x[10]) );
  MUX2_X1 prince_inst_S_58__mux_inv_x1_U1 ( .A(prince_inst_srin_x[58]), .B(
        prince_inst_xout_x[58]), .S(prince_inst_n26), .Z(prince_inst_sin_x[58]) );
  MUX2_X1 prince_inst_S_58__mux_inv_y1_U1 ( .A(prince_inst_srin_y[58]), .B(
        prince_inst_srin_y[26]), .S(prince_inst_n26), .Z(prince_inst_sin_y[58]) );
  MUX2_X1 prince_inst_S_58__mux_inv_x2_U1 ( .A(final_x[10]), .B(
        prince_inst_sout_x[58]), .S(prince_inst_n23), .Z(prince_inst_min_x[58]) );
  MUX2_X1 prince_inst_S_58__mux_inv_y2_U1 ( .A(final_y[10]), .B(final_y[10]), 
        .S(inv_sig2), .Z(prince_inst_min_y[58]) );
  XOR2_X1 prince_inst_S_59__x_U1 ( .A(rc[59]), .B(prince_inst_srin_x[27]), .Z(
        prince_inst_xout_x[59]) );
  XOR2_X1 prince_inst_S_59__srx_U1 ( .A(prince_inst_rc2_inv[59]), .B(
        prince_inst_sout_x[59]), .Z(final_x[11]) );
  MUX2_X1 prince_inst_S_59__mux_inv_x1_U1 ( .A(prince_inst_srin_x[59]), .B(
        prince_inst_xout_x[59]), .S(inv_sig), .Z(prince_inst_sin_x[59]) );
  MUX2_X1 prince_inst_S_59__mux_inv_y1_U1 ( .A(prince_inst_srin_y[59]), .B(
        prince_inst_srin_y[27]), .S(inv_sig), .Z(prince_inst_sin_y[59]) );
  MUX2_X1 prince_inst_S_59__mux_inv_x2_U1 ( .A(final_x[11]), .B(
        prince_inst_sout_x[59]), .S(prince_inst_n23), .Z(prince_inst_min_x[59]) );
  MUX2_X1 prince_inst_S_59__mux_inv_y2_U1 ( .A(final_y[11]), .B(final_y[11]), 
        .S(prince_inst_n20), .Z(prince_inst_min_y[59]) );
  XOR2_X1 prince_inst_S_60__x_U1 ( .A(rc[60]), .B(prince_inst_srin_x[60]), .Z(
        prince_inst_xout_x[60]) );
  XOR2_X1 prince_inst_S_60__srx_U1 ( .A(prince_inst_rc2_inv[60]), .B(
        prince_inst_sout_x[60]), .Z(final_x[60]) );
  MUX2_X1 prince_inst_S_60__mux_inv_x1_U1 ( .A(prince_inst_srin_x[60]), .B(
        prince_inst_xout_x[60]), .S(prince_inst_n28), .Z(prince_inst_sin_x[60]) );
  MUX2_X1 prince_inst_S_60__mux_inv_y1_U1 ( .A(prince_inst_srin_y[60]), .B(
        prince_inst_srin_y[60]), .S(inv_sig), .Z(prince_inst_sin_y[60]) );
  MUX2_X1 prince_inst_S_60__mux_inv_x2_U1 ( .A(final_x[60]), .B(
        prince_inst_sout_x[60]), .S(prince_inst_n23), .Z(prince_inst_min_x[60]) );
  MUX2_X1 prince_inst_S_60__mux_inv_y2_U1 ( .A(final_y[60]), .B(final_y[60]), 
        .S(inv_sig2), .Z(prince_inst_min_y[60]) );
  XOR2_X1 prince_inst_S_61__x_U1 ( .A(rc[61]), .B(prince_inst_srin_x[61]), .Z(
        prince_inst_xout_x[61]) );
  XOR2_X1 prince_inst_S_61__srx_U1 ( .A(prince_inst_rc2_inv[61]), .B(
        prince_inst_sout_x[61]), .Z(final_x[61]) );
  MUX2_X1 prince_inst_S_61__mux_inv_x1_U1 ( .A(prince_inst_srin_x[61]), .B(
        prince_inst_xout_x[61]), .S(prince_inst_n31), .Z(prince_inst_sin_x[61]) );
  MUX2_X1 prince_inst_S_61__mux_inv_y1_U1 ( .A(prince_inst_srin_y[61]), .B(
        prince_inst_srin_y[61]), .S(prince_inst_n26), .Z(prince_inst_sin_y[61]) );
  MUX2_X1 prince_inst_S_61__mux_inv_x2_U1 ( .A(final_x[61]), .B(
        prince_inst_sout_x[61]), .S(prince_inst_n23), .Z(prince_inst_min_x[61]) );
  MUX2_X1 prince_inst_S_61__mux_inv_y2_U1 ( .A(final_y[61]), .B(final_y[61]), 
        .S(prince_inst_n24), .Z(prince_inst_min_y[61]) );
  XOR2_X1 prince_inst_S_62__x_U1 ( .A(rc[62]), .B(prince_inst_srin_x[62]), .Z(
        prince_inst_xout_x[62]) );
  XOR2_X1 prince_inst_S_62__srx_U1 ( .A(prince_inst_rc2_inv[62]), .B(
        prince_inst_sout_x[62]), .Z(final_x[62]) );
  MUX2_X1 prince_inst_S_62__mux_inv_x1_U1 ( .A(prince_inst_srin_x[62]), .B(
        prince_inst_xout_x[62]), .S(prince_inst_n29), .Z(prince_inst_sin_x[62]) );
  MUX2_X1 prince_inst_S_62__mux_inv_y1_U1 ( .A(prince_inst_srin_y[62]), .B(
        prince_inst_srin_y[62]), .S(prince_inst_n26), .Z(prince_inst_sin_y[62]) );
  MUX2_X1 prince_inst_S_62__mux_inv_x2_U1 ( .A(final_x[62]), .B(
        prince_inst_sout_x[62]), .S(prince_inst_n24), .Z(prince_inst_min_x[62]) );
  MUX2_X1 prince_inst_S_62__mux_inv_y2_U1 ( .A(final_y[62]), .B(final_y[62]), 
        .S(inv_sig2), .Z(prince_inst_min_y[62]) );
  XOR2_X1 prince_inst_S_63__x_U1 ( .A(rc[63]), .B(prince_inst_srin_x[63]), .Z(
        prince_inst_xout_x[63]) );
  XOR2_X1 prince_inst_S_63__srx_U1 ( .A(prince_inst_rc2_inv[63]), .B(
        prince_inst_sout_x[63]), .Z(final_x[63]) );
  MUX2_X1 prince_inst_S_63__mux_inv_x1_U1 ( .A(prince_inst_srin_x[63]), .B(
        prince_inst_xout_x[63]), .S(inv_sig), .Z(prince_inst_sin_x[63]) );
  MUX2_X1 prince_inst_S_63__mux_inv_y1_U1 ( .A(prince_inst_srin_y[63]), .B(
        prince_inst_srin_y[63]), .S(inv_sig), .Z(prince_inst_sin_y[63]) );
  MUX2_X1 prince_inst_S_63__mux_inv_x2_U1 ( .A(final_x[63]), .B(
        prince_inst_sout_x[63]), .S(prince_inst_n24), .Z(prince_inst_min_x[63]) );
  MUX2_X1 prince_inst_S_63__mux_inv_y2_U1 ( .A(final_y[63]), .B(final_y[63]), 
        .S(prince_inst_n21), .Z(prince_inst_min_y[63]) );
  INV_X1 prince_inst_sbox_inst0_U7 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst0_n13) );
  INV_X1 prince_inst_sbox_inst0_U6 ( .A(inv_sig), .ZN(
        prince_inst_sbox_inst0_n11) );
  INV_X4 prince_inst_sbox_inst0_U5 ( .A(prince_inst_sbox_inst0_n13), .ZN(
        prince_inst_sbox_inst0_n12) );
  INV_X1 prince_inst_sbox_inst0_U4 ( .A(prince_inst_sbox_inst0_n11), .ZN(
        prince_inst_sbox_inst0_n9) );
  INV_X1 prince_inst_sbox_inst0_U3 ( .A(prince_inst_sbox_inst0_n11), .ZN(
        prince_inst_sbox_inst0_n10) );
  INV_X1 prince_inst_sbox_inst0_U2 ( .A(rst), .ZN(prince_inst_sbox_inst0_n8)
         );
  INV_X2 prince_inst_sbox_inst0_U1 ( .A(prince_inst_sbox_inst0_n8), .ZN(
        prince_inst_sbox_inst0_n7) );
  NAND3_X1 prince_inst_sbox_inst0_xxxy_inst_U28 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n20), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n19), .A3(prince_inst_sin_x[0]), .ZN(
        prince_inst_sbox_inst0_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n18), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n17), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n19) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U26 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sbox_inst0_xxxy_inst_n16), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n20) );
  NAND3_X1 prince_inst_sbox_inst0_xxxy_inst_U25 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n15), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n14), .A3(
        prince_inst_sbox_inst0_xxxy_inst_n13), .ZN(
        prince_inst_sbox_inst0_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst0_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n18), .A2(prince_inst_sin_x[2]), .A3(
        prince_inst_sin_x[0]), .A4(prince_inst_sin_y[3]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n13) );
  NAND3_X1 prince_inst_sbox_inst0_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n12), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n11), .A3(prince_inst_sin_x[2]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n14) );
  NAND4_X1 prince_inst_sbox_inst0_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n10), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n17), .A3(
        prince_inst_sbox_inst0_xxxy_inst_n11), .A4(prince_inst_sin_x[0]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n15) );
  XOR2_X1 prince_inst_sbox_inst0_xxxy_inst_U21 ( .A(
        prince_inst_sbox_inst0_xxxy_inst_n9), .B(prince_inst_sin_y[3]), .Z(
        prince_inst_sbox_inst0_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U20 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n8), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n7), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n9) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U19 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sbox_inst0_xxxy_inst_n11), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n8) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U18 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n6), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n5), .ZN(
        prince_inst_sbox_inst0_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst0_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n16), .A2(prince_inst_sin_x[2]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n5) );
  NAND3_X1 prince_inst_sbox_inst0_xxxy_inst_U16 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sin_y[3]), .A3(prince_inst_sbox_inst0_xxxy_inst_n18), 
        .ZN(prince_inst_sbox_inst0_xxxy_inst_n6) );
  NAND3_X1 prince_inst_sbox_inst0_xxxy_inst_U15 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n10), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n7), .A3(
        prince_inst_sbox_inst0_xxxy_inst_n4), .ZN(
        prince_inst_sbox_inst0_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst0_xxxy_inst_U14 ( .A(prince_inst_sin_x[0]), .B(
        prince_inst_sbox_inst0_xxxy_inst_n11), .S(
        prince_inst_sbox_inst0_xxxy_inst_n17), .Z(
        prince_inst_sbox_inst0_xxxy_inst_n4) );
  INV_X1 prince_inst_sbox_inst0_xxxy_inst_U13 ( .A(prince_inst_sin_y[3]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n17) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U12 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n11), .A2(prince_inst_sin_x[0]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n7) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U11 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n3), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n16), .ZN(
        prince_inst_sbox_inst0_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst0_xxxy_inst_U10 ( .A(
        prince_inst_sbox_inst0_xxxy_inst_n10), .B(
        prince_inst_sbox_inst0_xxxy_inst_n3), .S(
        prince_inst_sbox_inst0_xxxy_inst_n2), .Z(
        prince_inst_sbox_inst0_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U9 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sbox_inst0_xxxy_inst_n16), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n2) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U8 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n11), .A2(prince_inst_sin_y[3]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n16) );
  INV_X1 prince_inst_sbox_inst0_xxxy_inst_U7 ( .A(
        prince_inst_sbox_inst0_xxxy_inst_n18), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n11) );
  INV_X1 prince_inst_sbox_inst0_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst0_t1_sh[0]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n3) );
  INV_X1 prince_inst_sbox_inst0_xxxy_inst_U5 ( .A(prince_inst_sin_x[2]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n10) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U4 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sbox_inst0_xxxy_inst_n1), .ZN(
        prince_inst_sbox_inst0_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst0_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst0_xxxy_inst_n18), .A2(
        prince_inst_sbox_inst0_xxxy_inst_n12), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n1) );
  INV_X1 prince_inst_sbox_inst0_xxxy_inst_U2 ( .A(prince_inst_sin_x[0]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n12) );
  INV_X1 prince_inst_sbox_inst0_xxxy_inst_U1 ( .A(prince_inst_sin_x[1]), .ZN(
        prince_inst_sbox_inst0_xxxy_inst_n18) );
  XOR2_X1 prince_inst_sbox_inst0_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst0_t1_sh[1]), .B(
        prince_inst_sbox_inst0_xxyx_inst_n18), .Z(
        prince_inst_sbox_inst0_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst0_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n17), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n16), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n18) );
  XOR2_X1 prince_inst_sbox_inst0_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst0_xxyx_inst_n15), .B(
        prince_inst_sbox_inst0_xxyx_inst_n14), .Z(
        prince_inst_sbox_inst0_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U23 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_xxyx_inst_n14)
         );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n13), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n12), .ZN(
        prince_inst_sbox_inst0_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst0_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n11), .A2(prince_inst_sin_x[3]), .A3(
        prince_inst_sin_x[0]), .ZN(prince_inst_sbox_inst0_xxyx_inst_n12) );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n10), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n9), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n11) );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n15), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n8), .ZN(
        prince_inst_sbox_inst0_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst0_xxyx_inst_U18 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sbox_inst0_xxyx_inst_n17), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n15) );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n7), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n8), .ZN(
        prince_inst_sbox_inst0_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst0_xxyx_inst_U16 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sin_x[0]), .A3(prince_inst_sbox_inst0_xxyx_inst_n16), 
        .ZN(prince_inst_sbox_inst0_xxyx_inst_n8) );
  NAND3_X1 prince_inst_sbox_inst0_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n9), .A2(prince_inst_sin_x[3]), .A3(
        prince_inst_sin_x[1]), .ZN(prince_inst_sbox_inst0_xxyx_inst_n7) );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n6), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n13), .ZN(
        prince_inst_sbox_inst0_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst0_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst0_xxyx_inst_n17), .B(
        prince_inst_sbox_inst0_xxyx_inst_n16), .Z(
        prince_inst_sbox_inst0_xxyx_inst_n13) );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U12 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sin_y[2]), .ZN(prince_inst_sbox_inst0_xxyx_inst_n17)
         );
  NOR4_X1 prince_inst_sbox_inst0_xxyx_inst_U11 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sbox_inst0_xxyx_inst_n5), .A3(
        prince_inst_sbox_inst0_xxyx_inst_n4), .A4(
        prince_inst_sbox_inst0_xxyx_inst_n3), .ZN(
        prince_inst_sbox_inst0_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst0_xxyx_inst_U10 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_xxyx_inst_n3) );
  NOR2_X1 prince_inst_sbox_inst0_xxyx_inst_U9 ( .A1(prince_inst_sin_x[3]), 
        .A2(prince_inst_sbox_inst0_xxyx_inst_n9), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n4) );
  NOR2_X1 prince_inst_sbox_inst0_xxyx_inst_U8 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sbox_inst0_xxyx_inst_n9), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n5) );
  INV_X1 prince_inst_sbox_inst0_xxyx_inst_U7 ( .A(prince_inst_sin_y[2]), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n9) );
  NAND2_X1 prince_inst_sbox_inst0_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n2), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n1), .ZN(
        prince_inst_sbox_inst0_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst0_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n16), .A2(prince_inst_sin_x[1]), .A3(
        prince_inst_sin_y[2]), .A4(prince_inst_sin_x[0]), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n1) );
  INV_X1 prince_inst_sbox_inst0_xxyx_inst_U4 ( .A(prince_inst_sin_x[3]), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n16) );
  NAND4_X1 prince_inst_sbox_inst0_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst0_xxyx_inst_n10), .A2(
        prince_inst_sbox_inst0_xxyx_inst_n6), .A3(prince_inst_sin_x[3]), .A4(
        prince_inst_sin_y[2]), .ZN(prince_inst_sbox_inst0_xxyx_inst_n2) );
  INV_X1 prince_inst_sbox_inst0_xxyx_inst_U2 ( .A(prince_inst_sin_x[0]), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n6) );
  INV_X1 prince_inst_sbox_inst0_xxyx_inst_U1 ( .A(prince_inst_sin_x[1]), .ZN(
        prince_inst_sbox_inst0_xxyx_inst_n10) );
  XNOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst0_xyxx_inst_n22), .B(
        prince_inst_sbox_inst0_xyxx_inst_n21), .ZN(
        prince_inst_sbox_inst0_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n20), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n19), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n21) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n18), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n17), .ZN(
        prince_inst_sbox_inst0_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst0_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n16), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n15), .A3(
        prince_inst_sbox_inst0_xyxx_inst_n14), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n17) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U26 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sbox_inst0_xyxx_inst_n13), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n14) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U25 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_xyxx_inst_n13)
         );
  MUX2_X1 prince_inst_sbox_inst0_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst0_xyxx_inst_n20), .B(
        prince_inst_sbox_inst0_s0_sh[2]), .S(
        prince_inst_sbox_inst0_xyxx_inst_n12), .Z(
        prince_inst_sbox_inst0_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst0_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n22), .A2(prince_inst_sin_x[3]), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n12) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n20), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n11), .ZN(
        prince_inst_sbox_inst0_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U21 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sbox_inst0_xyxx_inst_n22), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n11) );
  INV_X1 prince_inst_sbox_inst0_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst0_xyxx_inst_n10), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n22) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n19), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n9), .ZN(
        prince_inst_sbox_inst0_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n8), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n16), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n9) );
  INV_X1 prince_inst_sbox_inst0_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst0_xyxx_inst_n7), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n16) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n15), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n10), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n8) );
  NAND2_X1 prince_inst_sbox_inst0_xyxx_inst_U15 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sin_x[0]), .ZN(prince_inst_sbox_inst0_xyxx_inst_n10)
         );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n18), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n7), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n19) );
  NAND2_X1 prince_inst_sbox_inst0_xyxx_inst_U13 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_xyxx_inst_n7) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U12 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sin_x[2]), .ZN(prince_inst_sbox_inst0_xyxx_inst_n18)
         );
  XNOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst0_xyxx_inst_n6), .B(
        prince_inst_sbox_inst0_xyxx_inst_n5), .ZN(
        prince_inst_sbox_inst0_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst0_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n20), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n4), .A3(
        prince_inst_sbox_inst0_xyxx_inst_n3), .ZN(
        prince_inst_sbox_inst0_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst0_xyxx_inst_U9 ( .A(prince_inst_sin_x[3]), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n3) );
  AND2_X1 prince_inst_sbox_inst0_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n2), .A2(prince_inst_sin_x[0]), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n4) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n2), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n15), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n20) );
  OR2_X1 prince_inst_sbox_inst0_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst0_xyxx_inst_n6), .A2(
        prince_inst_sbox_inst0_xyxx_inst_n1), .ZN(
        prince_inst_sbox_inst0_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst0_xyxx_inst_U5 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sbox_inst0_xyxx_inst_n5), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n1) );
  NAND2_X1 prince_inst_sbox_inst0_xyxx_inst_U4 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_xyxx_inst_n5) );
  NOR3_X1 prince_inst_sbox_inst0_xyxx_inst_U3 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sbox_inst0_xyxx_inst_n15), .A3(
        prince_inst_sbox_inst0_xyxx_inst_n2), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n6) );
  INV_X1 prince_inst_sbox_inst0_xyxx_inst_U2 ( .A(prince_inst_sin_y[1]), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n2) );
  INV_X1 prince_inst_sbox_inst0_xyxx_inst_U1 ( .A(prince_inst_sin_x[2]), .ZN(
        prince_inst_sbox_inst0_xyxx_inst_n15) );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n31), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n30), .ZN(
        prince_inst_sbox_inst0_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst0_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst0_xyyy_inst_n29), .B(
        prince_inst_sbox_inst0_xyyy_inst_n28), .Z(
        prince_inst_sbox_inst0_xyyy_inst_n31) );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n27), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n26), .ZN(
        prince_inst_sbox_inst0_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst0_xyyy_inst_U25 ( .A1(prince_inst_sin_y[2]), 
        .A2(prince_inst_sin_y[3]), .A3(prince_inst_sbox_inst0_xyyy_inst_n30), 
        .ZN(prince_inst_sbox_inst0_xyyy_inst_n26) );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U24 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sbox_inst0_xyyy_inst_n25), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n30) );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U23 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sbox_inst0_xyyy_inst_n24), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n27) );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n23), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n22), .ZN(
        prince_inst_sbox_inst0_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n21), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n20), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n22) );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n24), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n25), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n23) );
  NOR3_X1 prince_inst_sbox_inst0_xyyy_inst_U19 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sin_y[2]), .A3(prince_inst_sbox_inst0_xyyy_inst_n20), 
        .ZN(prince_inst_sbox_inst0_xyyy_inst_n24) );
  MUX2_X1 prince_inst_sbox_inst0_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst0_xyyy_inst_n19), .B(
        prince_inst_sbox_inst0_xyyy_inst_n18), .S(
        prince_inst_sbox_inst0_xyyy_inst_n17), .Z(
        prince_inst_sbox_inst0_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst0_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n18), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n21), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n19) );
  NOR2_X1 prince_inst_sbox_inst0_xyyy_inst_U16 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sbox_inst0_xyyy_inst_n16), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n21) );
  INV_X1 prince_inst_sbox_inst0_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst0_xyyy_inst_n15), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n16) );
  NOR3_X1 prince_inst_sbox_inst0_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n14), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n13), .A3(
        prince_inst_sbox_inst0_xyyy_inst_n28), .ZN(
        prince_inst_sbox_inst0_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst0_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n12), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n18), .A3(
        prince_inst_sbox_inst0_xyyy_inst_n20), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n13) );
  INV_X1 prince_inst_sbox_inst0_xyyy_inst_U12 ( .A(prince_inst_sin_y[3]), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n20) );
  NOR2_X1 prince_inst_sbox_inst0_xyyy_inst_U11 ( .A1(prince_inst_sin_y[3]), 
        .A2(prince_inst_sbox_inst0_xyyy_inst_n15), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n14) );
  MUX2_X1 prince_inst_sbox_inst0_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst0_t1_sh[3]), .B(
        prince_inst_sbox_inst0_xyyy_inst_n18), .S(
        prince_inst_sbox_inst0_xyyy_inst_n28), .Z(
        prince_inst_sbox_inst0_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst0_xyyy_inst_U9 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sbox_inst0_xyyy_inst_n17), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n28) );
  AND2_X1 prince_inst_sbox_inst0_xyyy_inst_U8 ( .A1(prince_inst_sin_x[0]), 
        .A2(prince_inst_sin_y[3]), .ZN(prince_inst_sbox_inst0_xyyy_inst_n17)
         );
  AND2_X1 prince_inst_sbox_inst0_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n29), .A2(
        prince_inst_sbox_inst0_t1_sh[3]), .ZN(prince_inst_sbox_inst0_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst0_xyyy_inst_U6 ( .A1(prince_inst_sin_y[3]), 
        .A2(prince_inst_sbox_inst0_xyyy_inst_n15), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n29) );
  NOR2_X1 prince_inst_sbox_inst0_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n25), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n18), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n15) );
  INV_X1 prince_inst_sbox_inst0_xyyy_inst_U4 ( .A(prince_inst_sin_y[1]), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n25) );
  NOR2_X1 prince_inst_sbox_inst0_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst0_xyyy_inst_n18), .A2(
        prince_inst_sbox_inst0_xyyy_inst_n12), .ZN(
        prince_inst_sbox_inst0_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst0_xyyy_inst_U2 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sin_x[0]), .ZN(prince_inst_sbox_inst0_xyyy_inst_n12)
         );
  INV_X1 prince_inst_sbox_inst0_xyyy_inst_U1 ( .A(prince_inst_sin_y[2]), .ZN(
        prince_inst_sbox_inst0_xyyy_inst_n18) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n21), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n20), .ZN(
        prince_inst_sbox_inst0_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U27 ( .A1(prince_inst_sin_y[0]), 
        .A2(prince_inst_sbox_inst0_yxxx_inst_n19), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n20) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n18), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n17), .ZN(
        prince_inst_sbox_inst0_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n16), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n15), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n17) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U24 ( .A1(prince_inst_sin_y[0]), 
        .A2(prince_inst_sbox_inst0_yxxx_inst_n14), .ZN(
        prince_inst_sbox_inst0_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n19), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n13), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n14) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n12), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n11), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n13) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U21 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_yxxx_inst_n11)
         );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n10), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n15), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n19) );
  INV_X1 prince_inst_sbox_inst0_yxxx_inst_U19 ( .A(prince_inst_sin_x[3]), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n15) );
  MUX2_X1 prince_inst_sbox_inst0_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst0_yxxx_inst_n9), .B(
        prince_inst_sbox_inst0_yxxx_inst_n8), .S(
        prince_inst_sbox_inst0_yxxx_inst_n7), .Z(
        prince_inst_sbox_inst0_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n10), .A2(prince_inst_sin_x[3]), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n9) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n18), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n6), .ZN(
        prince_inst_sbox_inst0_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n5), .A2(prince_inst_sin_y[0]), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n6) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n4), .A2(prince_inst_sin_x[3]), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n5) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U13 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sbox_inst0_yxxx_inst_n12), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n4) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n3), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n7), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n18) );
  XNOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst0_yxxx_inst_n16), .B(
        prince_inst_sbox_inst0_yxxx_inst_n2), .ZN(
        prince_inst_sbox_inst0_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst0_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n3), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n16), .ZN(
        prince_inst_sbox_inst0_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst0_yxxx_inst_U9 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sbox_inst0_yxxx_inst_n7), .A3(
        prince_inst_sbox_inst0_yxxx_inst_n12), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n16) );
  INV_X1 prince_inst_sbox_inst0_yxxx_inst_U8 ( .A(prince_inst_sin_x[2]), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n12) );
  NOR2_X1 prince_inst_sbox_inst0_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n10), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n2), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n3) );
  OR2_X1 prince_inst_sbox_inst0_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst0_yxxx_inst_n8), .A2(
        prince_inst_sbox_inst0_yxxx_inst_n21), .ZN(
        prince_inst_sbox_inst0_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst0_yxxx_inst_U5 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sbox_inst0_yxxx_inst_n10), .A3(
        prince_inst_sbox_inst0_yxxx_inst_n7), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n21) );
  INV_X1 prince_inst_sbox_inst0_yxxx_inst_U4 ( .A(prince_inst_sin_y[0]), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n7) );
  INV_X1 prince_inst_sbox_inst0_yxxx_inst_U3 ( .A(prince_inst_sin_x[1]), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n10) );
  INV_X1 prince_inst_sbox_inst0_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst0_yxxx_inst_n2), .ZN(
        prince_inst_sbox_inst0_yxxx_inst_n8) );
  NAND2_X1 prince_inst_sbox_inst0_yxxx_inst_U1 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_yxxx_inst_n2) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n19), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n18), .ZN(
        prince_inst_sbox_inst0_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst0_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n17), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n18), .A3(
        prince_inst_sbox_inst0_yxyy_inst_n19), .ZN(
        prince_inst_sbox_inst0_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst0_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n16), .A2(prince_inst_sin_x[1]), .A3(
        prince_inst_sin_y[3]), .ZN(prince_inst_sbox_inst0_yxyy_inst_n18) );
  NAND3_X1 prince_inst_sbox_inst0_yxyy_inst_U24 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n15), .A2(prince_inst_sin_y[2]), .A3(
        prince_inst_sin_y[3]), .ZN(prince_inst_sbox_inst0_yxyy_inst_n17) );
  MUX2_X1 prince_inst_sbox_inst0_yxyy_inst_U23 ( .A(
        prince_inst_sbox_inst0_yxyy_inst_n14), .B(
        prince_inst_sbox_inst0_yxyy_inst_n13), .S(prince_inst_sin_y[0]), .Z(
        prince_inst_sbox_inst0_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst0_yxyy_inst_U22 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n16), .A2(prince_inst_sin_x[1]), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n13) );
  MUX2_X1 prince_inst_sbox_inst0_yxyy_inst_U21 ( .A(prince_inst_sin_x[1]), .B(
        prince_inst_sbox_inst0_yxyy_inst_n12), .S(
        prince_inst_sbox_inst0_yxyy_inst_n16), .Z(
        prince_inst_sbox_inst0_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n11), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n10), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n12) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n15), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n9), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n11) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U18 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n8), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n7), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n9) );
  MUX2_X1 prince_inst_sbox_inst0_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst0_yxyy_inst_n14), .B(
        prince_inst_sbox_inst0_yxyy_inst_n6), .S(
        prince_inst_sbox_inst0_yxyy_inst_n7), .Z(
        prince_inst_sbox_inst0_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst0_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst0_yxyy_inst_n5), .B(
        prince_inst_sbox_inst0_yxyy_inst_n6), .Z(
        prince_inst_sbox_inst0_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst0_yxyy_inst_U15 ( .A(
        prince_inst_sbox_inst0_yxyy_inst_n19), .B(
        prince_inst_sbox_inst0_yxyy_inst_n10), .Z(
        prince_inst_sbox_inst0_yxyy_inst_n5) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U14 ( .A1(prince_inst_sin_y[3]), 
        .A2(prince_inst_sin_y[0]), .ZN(prince_inst_sbox_inst0_yxyy_inst_n10)
         );
  NOR4_X1 prince_inst_sbox_inst0_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n4), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n6), .A3(
        prince_inst_sbox_inst0_yxyy_inst_n14), .A4(
        prince_inst_sbox_inst0_yxyy_inst_n7), .ZN(
        prince_inst_sbox_inst0_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst0_yxyy_inst_U12 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n15), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n8), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n14) );
  INV_X1 prince_inst_sbox_inst0_yxyy_inst_U11 ( .A(
        prince_inst_sbox_inst0_yxyy_inst_n19), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n4) );
  NAND3_X1 prince_inst_sbox_inst0_yxyy_inst_U10 ( .A1(prince_inst_sin_x[1]), 
        .A2(prince_inst_sin_y[2]), .A3(prince_inst_sin_y[0]), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n19) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U9 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n3), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n2), .ZN(
        prince_inst_sbox_inst0_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U8 ( .A1(prince_inst_sin_y[3]), 
        .A2(prince_inst_sbox_inst0_yxyy_inst_n1), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n2) );
  NAND2_X1 prince_inst_sbox_inst0_yxyy_inst_U7 ( .A1(prince_inst_sin_y[2]), 
        .A2(prince_inst_sin_x[1]), .ZN(prince_inst_sbox_inst0_yxyy_inst_n1) );
  OR3_X1 prince_inst_sbox_inst0_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n6), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n15), .A3(
        prince_inst_sbox_inst0_yxyy_inst_n7), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n3) );
  INV_X1 prince_inst_sbox_inst0_yxyy_inst_U5 ( .A(prince_inst_sin_y[0]), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n7) );
  INV_X1 prince_inst_sbox_inst0_yxyy_inst_U4 ( .A(prince_inst_sin_x[1]), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n15) );
  NOR2_X1 prince_inst_sbox_inst0_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst0_yxyy_inst_n16), .A2(
        prince_inst_sbox_inst0_yxyy_inst_n8), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n6) );
  INV_X1 prince_inst_sbox_inst0_yxyy_inst_U2 ( .A(prince_inst_sin_y[3]), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n8) );
  INV_X1 prince_inst_sbox_inst0_yxyy_inst_U1 ( .A(prince_inst_sin_y[2]), .ZN(
        prince_inst_sbox_inst0_yxyy_inst_n16) );
  NOR2_X1 prince_inst_sbox_inst0_yyxy_inst_U24 ( .A1(prince_inst_sin_y[0]), 
        .A2(prince_inst_sbox_inst0_yyxy_inst_n16), .ZN(
        prince_inst_sbox_inst0_s3_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst0_yyxy_inst_U23 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n15), .A2(
        prince_inst_sbox_inst0_yyxy_inst_n14), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n16) );
  NAND2_X1 prince_inst_sbox_inst0_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n13), .A2(
        prince_inst_sbox_inst0_yyxy_inst_n12), .ZN(
        prince_inst_sbox_inst0_t2_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst0_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n11), .A2(prince_inst_sin_y[1]), .A3(
        prince_inst_sin_y[3]), .ZN(prince_inst_sbox_inst0_yyxy_inst_n12) );
  NAND3_X1 prince_inst_sbox_inst0_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n10), .A2(prince_inst_sin_y[0]), .A3(
        prince_inst_sin_x[2]), .ZN(prince_inst_sbox_inst0_yyxy_inst_n13) );
  MUX2_X1 prince_inst_sbox_inst0_yyxy_inst_U19 ( .A(
        prince_inst_sbox_inst0_yyxy_inst_n15), .B(
        prince_inst_sbox_inst0_yyxy_inst_n9), .S(
        prince_inst_sbox_inst0_yyxy_inst_n11), .Z(
        prince_inst_sbox_inst0_t3_sh[6]) );
  INV_X1 prince_inst_sbox_inst0_yyxy_inst_U18 ( .A(prince_inst_sin_y[0]), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n11) );
  AND3_X1 prince_inst_sbox_inst0_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n8), .A2(
        prince_inst_sbox_inst0_yyxy_inst_n10), .A3(prince_inst_sin_y[3]), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n9) );
  NOR3_X1 prince_inst_sbox_inst0_yyxy_inst_U16 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sin_y[3]), .A3(prince_inst_sbox_inst0_yyxy_inst_n10), 
        .ZN(prince_inst_sbox_inst0_yyxy_inst_n15) );
  NAND2_X1 prince_inst_sbox_inst0_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n7), .A2(
        prince_inst_sbox_inst0_yyxy_inst_n6), .ZN(
        prince_inst_sbox_inst0_s0_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst0_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n8), .A2(prince_inst_sin_y[1]), .A3(
        prince_inst_sin_y[0]), .ZN(prince_inst_sbox_inst0_yyxy_inst_n7) );
  NAND2_X1 prince_inst_sbox_inst0_yyxy_inst_U13 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n5), .A2(
        prince_inst_sbox_inst0_yyxy_inst_n4), .ZN(
        prince_inst_sbox_inst0_s2_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst0_yyxy_inst_U12 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n10), .A2(prince_inst_sin_y[3]), .A3(
        prince_inst_sin_y[0]), .ZN(prince_inst_sbox_inst0_yyxy_inst_n5) );
  MUX2_X1 prince_inst_sbox_inst0_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst0_yyxy_inst_n3), .B(
        prince_inst_sbox_inst0_yyxy_inst_n2), .S(prince_inst_sin_y[0]), .Z(
        prince_inst_sbox_inst0_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst0_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n10), .A2(prince_inst_sin_y[3]), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n2) );
  INV_X1 prince_inst_sbox_inst0_yyxy_inst_U9 ( .A(prince_inst_sin_y[1]), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n10) );
  INV_X1 prince_inst_sbox_inst0_yyxy_inst_U8 ( .A(
        prince_inst_sbox_inst0_yyxy_inst_n6), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n3) );
  OR2_X1 prince_inst_sbox_inst0_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n14), .A2(
        prince_inst_sbox_inst0_s1_sh[6]), .ZN(prince_inst_sbox_inst0_t1_sh[6])
         );
  NOR2_X1 prince_inst_sbox_inst0_yyxy_inst_U6 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sbox_inst0_yyxy_inst_n6), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n14) );
  NAND2_X1 prince_inst_sbox_inst0_yyxy_inst_U5 ( .A1(prince_inst_sin_x[2]), 
        .A2(prince_inst_sin_y[3]), .ZN(prince_inst_sbox_inst0_yyxy_inst_n6) );
  NAND2_X1 prince_inst_sbox_inst0_yyxy_inst_U4 ( .A1(
        prince_inst_sbox_inst0_yyxy_inst_n1), .A2(
        prince_inst_sbox_inst0_yyxy_inst_n4), .ZN(
        prince_inst_sbox_inst0_s1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst0_yyxy_inst_U3 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sin_y[3]), .A3(prince_inst_sbox_inst0_yyxy_inst_n8), 
        .ZN(prince_inst_sbox_inst0_yyxy_inst_n4) );
  INV_X1 prince_inst_sbox_inst0_yyxy_inst_U2 ( .A(prince_inst_sin_x[2]), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n8) );
  NAND3_X1 prince_inst_sbox_inst0_yyxy_inst_U1 ( .A1(prince_inst_sin_y[0]), 
        .A2(prince_inst_sin_y[1]), .A3(prince_inst_sin_x[2]), .ZN(
        prince_inst_sbox_inst0_yyxy_inst_n1) );
  XNOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst0_yyyx_inst_n38), .B(
        prince_inst_sbox_inst0_yyyx_inst_n37), .ZN(
        prince_inst_sbox_inst0_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst0_yyyx_inst_n36), .B(
        prince_inst_sbox_inst0_yyyx_inst_n35), .Z(
        prince_inst_sbox_inst0_yyyx_inst_n37) );
  XNOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst0_yyyx_inst_n34), .B(
        prince_inst_sbox_inst0_yyyx_inst_n38), .ZN(
        prince_inst_sbox_inst0_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst0_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n33), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n32), .ZN(
        prince_inst_sbox_inst0_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst0_yyyx_inst_U21 ( .A1(prince_inst_sin_x[3]), 
        .A2(prince_inst_sbox_inst0_yyyx_inst_n34), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n32) );
  NAND3_X1 prince_inst_sbox_inst0_yyyx_inst_U20 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sin_y[2]), .A3(prince_inst_sbox_inst0_yyyx_inst_n31), 
        .ZN(prince_inst_sbox_inst0_yyyx_inst_n33) );
  XNOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst0_yyyx_inst_n30), .B(
        prince_inst_sbox_inst0_yyyx_inst_n29), .ZN(
        prince_inst_sbox_inst0_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst0_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n36), .A2(prince_inst_sin_y[2]), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n30) );
  NAND3_X1 prince_inst_sbox_inst0_yyyx_inst_U17 ( .A1(prince_inst_sin_y[1]), 
        .A2(prince_inst_sin_y[0]), .A3(prince_inst_sin_y[2]), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n36) );
  NOR3_X1 prince_inst_sbox_inst0_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n28), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n27), .A3(
        prince_inst_sbox_inst0_yyyx_inst_n26), .ZN(
        prince_inst_sbox_inst0_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst0_yyyx_inst_U15 ( .A1(prince_inst_sin_x[3]), 
        .A2(prince_inst_sin_y[2]), .A3(prince_inst_sbox_inst0_yyyx_inst_n25), 
        .ZN(prince_inst_sbox_inst0_yyyx_inst_n26) );
  INV_X1 prince_inst_sbox_inst0_yyyx_inst_U14 ( .A(prince_inst_sin_y[0]), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n27) );
  NOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n38), .A2(prince_inst_sin_y[1]), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n28) );
  OR2_X1 prince_inst_sbox_inst0_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n24), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n23), .ZN(
        prince_inst_sbox_inst0_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U11 ( .A1(prince_inst_sin_y[0]), 
        .A2(prince_inst_sbox_inst0_yyyx_inst_n38), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n23) );
  NOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n25), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n35), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n24) );
  NAND2_X1 prince_inst_sbox_inst0_yyyx_inst_U9 ( .A1(prince_inst_sin_y[0]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_yyyx_inst_n35)
         );
  OR2_X1 prince_inst_sbox_inst0_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n34), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n22), .ZN(
        prince_inst_sbox_inst0_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n25), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n38), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n22) );
  AND3_X1 prince_inst_sbox_inst0_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n25), .A2(prince_inst_sin_y[0]), .A3(
        prince_inst_sin_y[2]), .ZN(prince_inst_sbox_inst0_yyyx_inst_n34) );
  AND2_X1 prince_inst_sbox_inst0_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n29), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n38), .ZN(
        prince_inst_sbox_inst0_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst0_yyyx_inst_U4 ( .A1(prince_inst_sin_x[3]), 
        .A2(prince_inst_sin_y[2]), .ZN(prince_inst_sbox_inst0_yyyx_inst_n38)
         );
  NOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst0_yyyx_inst_n31), .A2(
        prince_inst_sbox_inst0_yyyx_inst_n25), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n29) );
  INV_X1 prince_inst_sbox_inst0_yyyx_inst_U2 ( .A(prince_inst_sin_y[1]), .ZN(
        prince_inst_sbox_inst0_yyyx_inst_n25) );
  NOR2_X1 prince_inst_sbox_inst0_yyyx_inst_U1 ( .A1(prince_inst_sin_y[0]), 
        .A2(prince_inst_sin_x[3]), .ZN(prince_inst_sbox_inst0_yyyx_inst_n31)
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s00_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[0]), .B(prince_inst_sbox_inst0_s0_sh[0]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s01_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[1]), .B(prince_inst_sbox_inst0_s0_sh[1]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s02_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[2]), .B(prince_inst_sbox_inst0_s0_sh[2]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s03_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[3]), .B(prince_inst_sbox_inst0_s0_sh[3]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s04_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[4]), .B(prince_inst_sbox_inst0_s0_sh[4]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s05_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[5]), .B(prince_inst_sbox_inst0_s0_sh[5]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s06_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[6]), .B(prince_inst_sbox_inst0_s0_sh[6]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s07_U1 ( .A(
        prince_inst_sbox_inst0_t0_sh[7]), .B(prince_inst_sbox_inst0_s0_sh[7]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s10_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[0]), .B(prince_inst_sbox_inst0_s1_sh[0]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s11_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[1]), .B(prince_inst_sbox_inst0_s1_sh[1]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s12_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[2]), .B(prince_inst_sbox_inst0_s1_sh[2]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s13_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[3]), .B(prince_inst_sbox_inst0_s1_sh[3]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s14_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[4]), .B(prince_inst_sbox_inst0_s1_sh[4]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s15_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[5]), .B(prince_inst_sbox_inst0_s1_sh[5]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s16_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[6]), .B(prince_inst_sbox_inst0_s1_sh[6]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s17_U1 ( .A(
        prince_inst_sbox_inst0_t1_sh[7]), .B(prince_inst_sbox_inst0_s1_sh[7]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s20_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[0]), .B(prince_inst_sbox_inst0_s2_sh[0]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s21_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[1]), .B(prince_inst_sbox_inst0_s2_sh[1]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s22_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[2]), .B(prince_inst_sbox_inst0_s2_sh[2]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s23_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[3]), .B(prince_inst_sbox_inst0_s2_sh[3]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s24_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[4]), .B(prince_inst_sbox_inst0_s2_sh[4]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s25_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[5]), .B(prince_inst_sbox_inst0_s2_sh[5]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s26_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[6]), .B(prince_inst_sbox_inst0_s2_sh[6]), 
        .S(prince_inst_sbox_inst0_n9), .Z(prince_inst_sbox_inst0_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s27_U1 ( .A(
        prince_inst_sbox_inst0_t2_sh[7]), .B(prince_inst_sbox_inst0_s2_sh[7]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s30_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[0]), .B(prince_inst_sbox_inst0_s3_sh[0]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s31_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[1]), .B(prince_inst_sbox_inst0_s3_sh[1]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s32_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[2]), .B(prince_inst_sbox_inst0_s3_sh[2]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s33_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[3]), .B(prince_inst_sbox_inst0_s3_sh[3]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s34_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[4]), .B(prince_inst_sbox_inst0_s3_sh[4]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s35_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[5]), .B(prince_inst_sbox_inst0_s3_sh[5]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s36_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[6]), .B(prince_inst_sbox_inst0_s3_sh[6]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst0_mux_s37_U1 ( .A(
        prince_inst_sbox_inst0_t3_sh[7]), .B(prince_inst_sbox_inst0_s3_sh[7]), 
        .S(prince_inst_sbox_inst0_n10), .Z(prince_inst_sbox_inst0_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk0_U1 ( .A(r[0]), .B(
        prince_inst_sbox_inst0_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n4), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n3), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n5) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n3) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n2), .A2(
        prince_inst_sbox_inst0_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n4) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n2) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk0_reg_xr_n5), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk1_U1 ( .A(r[1]), .B(
        prince_inst_sbox_inst0_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk2_U1 ( .A(r[2]), .B(
        prince_inst_sbox_inst0_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk3_U1 ( .A(r[3]), .B(
        prince_inst_sbox_inst0_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk4_U1 ( .A(r[0]), .B(
        prince_inst_sbox_inst0_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk5_U1 ( .A(r[1]), .B(
        prince_inst_sbox_inst0_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk6_U1 ( .A(r[2]), .B(
        prince_inst_sbox_inst0_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_msk7_U1 ( .A(r[3]), .B(
        prince_inst_sbox_inst0_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst0_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst0_c_inst0_ax_n2), .B(
        prince_inst_sbox_inst0_c_inst0_ax_n1), .ZN(prince_inst_sout_x[0]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst0_c_inst0_y[1]), .B(
        prince_inst_sbox_inst0_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst0_c_inst0_ax_n1) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst0_c_inst0_y[2]), .B(
        prince_inst_sbox_inst0_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst0_c_inst0_ax_n2) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst0_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst0_c_inst0_ay_n5), .ZN(final_y[48]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst0_c_inst0_y[5]), .B(
        prince_inst_sbox_inst0_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst0_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst0_c_inst0_y[6]), .B(
        prince_inst_sbox_inst0_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst0_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk0_U1 ( .A(r[4]), .B(
        prince_inst_sbox_inst0_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk1_U1 ( .A(r[5]), .B(
        prince_inst_sbox_inst0_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk2_U1 ( .A(r[6]), .B(
        prince_inst_sbox_inst0_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk3_U1 ( .A(r[7]), .B(
        prince_inst_sbox_inst0_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk4_U1 ( .A(r[4]), .B(
        prince_inst_sbox_inst0_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk5_U1 ( .A(r[5]), .B(
        prince_inst_sbox_inst0_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk6_U1 ( .A(r[6]), .B(
        prince_inst_sbox_inst0_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_msk7_U1 ( .A(r[7]), .B(
        prince_inst_sbox_inst0_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst0_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst0_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst0_c_inst1_ax_n5), .ZN(prince_inst_sout_x[1]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst0_c_inst1_y[1]), .B(
        prince_inst_sbox_inst0_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst0_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst0_c_inst1_y[2]), .B(
        prince_inst_sbox_inst0_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst0_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst0_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst0_c_inst1_ay_n5), .ZN(final_y[49]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst0_c_inst1_y[5]), .B(
        prince_inst_sbox_inst0_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst0_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst0_c_inst1_y[6]), .B(
        prince_inst_sbox_inst0_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst0_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk0_U1 ( .A(r[8]), .B(
        prince_inst_sbox_inst0_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk1_U1 ( .A(r[9]), .B(
        prince_inst_sbox_inst0_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk2_U1 ( .A(r[10]), .B(
        prince_inst_sbox_inst0_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk3_U1 ( .A(r[11]), .B(
        prince_inst_sbox_inst0_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk4_U1 ( .A(r[8]), .B(
        prince_inst_sbox_inst0_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk5_U1 ( .A(r[9]), .B(
        prince_inst_sbox_inst0_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk6_U1 ( .A(r[10]), .B(
        prince_inst_sbox_inst0_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_msk7_U1 ( .A(r[11]), .B(
        prince_inst_sbox_inst0_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst0_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst0_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst0_c_inst2_ax_n5), .ZN(prince_inst_sout_x[2]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst0_c_inst2_y[1]), .B(
        prince_inst_sbox_inst0_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst0_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst0_c_inst2_y[2]), .B(
        prince_inst_sbox_inst0_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst0_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst0_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst0_c_inst2_ay_n5), .ZN(final_y[50]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst0_c_inst2_y[5]), .B(
        prince_inst_sbox_inst0_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst0_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst0_c_inst2_y[6]), .B(
        prince_inst_sbox_inst0_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst0_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk0_U1 ( .A(r[12]), .B(
        prince_inst_sbox_inst0_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk1_U1 ( .A(r[13]), .B(
        prince_inst_sbox_inst0_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk2_U1 ( .A(r[14]), .B(
        prince_inst_sbox_inst0_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk3_U1 ( .A(r[15]), .B(
        prince_inst_sbox_inst0_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk4_U1 ( .A(r[12]), .B(
        prince_inst_sbox_inst0_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk5_U1 ( .A(r[13]), .B(
        prince_inst_sbox_inst0_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk6_U1 ( .A(r[14]), .B(
        prince_inst_sbox_inst0_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_msk7_U1 ( .A(r[15]), .B(
        prince_inst_sbox_inst0_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst0_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst0_n7), .A3(
        prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst0_n12), .A2(prince_inst_sbox_inst0_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst0_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst0_n12), .ZN(
        prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst0_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst0_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst0_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst0_c_inst3_ax_n5), .ZN(prince_inst_sout_x[3]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst0_c_inst3_y[1]), .B(
        prince_inst_sbox_inst0_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst0_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst0_c_inst3_y[2]), .B(
        prince_inst_sbox_inst0_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst0_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst0_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst0_c_inst3_ay_n5), .ZN(final_y[51]) );
  XNOR2_X1 prince_inst_sbox_inst0_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst0_c_inst3_y[5]), .B(
        prince_inst_sbox_inst0_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst0_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst0_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst0_c_inst3_y[6]), .B(
        prince_inst_sbox_inst0_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst0_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst1_U7 ( .A(prince_inst_sbox_inst1_n13), .ZN(
        prince_inst_sbox_inst1_n12) );
  INV_X1 prince_inst_sbox_inst1_U6 ( .A(prince_inst_n29), .ZN(
        prince_inst_sbox_inst1_n11) );
  INV_X1 prince_inst_sbox_inst1_U5 ( .A(prince_inst_sbox_inst1_n11), .ZN(
        prince_inst_sbox_inst1_n10) );
  INV_X1 prince_inst_sbox_inst1_U4 ( .A(prince_inst_sbox_inst1_n11), .ZN(
        prince_inst_sbox_inst1_n9) );
  INV_X1 prince_inst_sbox_inst1_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst1_n13) );
  INV_X1 prince_inst_sbox_inst1_U2 ( .A(rst), .ZN(prince_inst_sbox_inst1_n8)
         );
  INV_X2 prince_inst_sbox_inst1_U1 ( .A(prince_inst_sbox_inst1_n8), .ZN(
        prince_inst_sbox_inst1_n7) );
  NAND3_X1 prince_inst_sbox_inst1_xxxy_inst_U28 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n70), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n69), .A3(prince_inst_sin_x[4]), .ZN(
        prince_inst_sbox_inst1_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n67), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n69) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U26 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n70) );
  NAND3_X1 prince_inst_sbox_inst1_xxxy_inst_U25 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n65), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n64), .A3(
        prince_inst_sbox_inst1_xxxy_inst_n63), .ZN(
        prince_inst_sbox_inst1_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst1_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n68), .A2(prince_inst_sin_x[6]), .A3(
        prince_inst_sin_x[4]), .A4(prince_inst_sin_y[7]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n63) );
  NAND3_X1 prince_inst_sbox_inst1_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n62), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n61), .A3(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n64) );
  NAND4_X1 prince_inst_sbox_inst1_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n67), .A3(
        prince_inst_sbox_inst1_xxxy_inst_n61), .A4(prince_inst_sin_x[4]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n65) );
  XOR2_X1 prince_inst_sbox_inst1_xxxy_inst_U21 ( .A(
        prince_inst_sbox_inst1_xxxy_inst_n59), .B(prince_inst_sin_y[7]), .Z(
        prince_inst_sbox_inst1_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U20 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U19 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n58) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U18 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst1_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst1_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n66), .A2(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst1_xxxy_inst_U16 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sin_y[7]), .A3(prince_inst_sbox_inst1_xxxy_inst_n68), 
        .ZN(prince_inst_sbox_inst1_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst1_xxxy_inst_U15 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst1_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst1_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst1_xxxy_inst_U14 ( .A(prince_inst_sin_x[4]), .B(
        prince_inst_sbox_inst1_xxxy_inst_n61), .S(
        prince_inst_sbox_inst1_xxxy_inst_n67), .Z(
        prince_inst_sbox_inst1_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst1_xxxy_inst_U13 ( .A(prince_inst_sin_y[7]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U12 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n61), .A2(prince_inst_sin_x[4]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U11 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst1_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst1_xxxy_inst_U10 ( .A(
        prince_inst_sbox_inst1_xxxy_inst_n60), .B(
        prince_inst_sbox_inst1_xxxy_inst_n53), .S(
        prince_inst_sbox_inst1_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst1_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U9 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sbox_inst1_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U8 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n61), .A2(prince_inst_sin_y[7]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n66) );
  INV_X1 prince_inst_sbox_inst1_xxxy_inst_U7 ( .A(
        prince_inst_sbox_inst1_xxxy_inst_n68), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst1_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst1_t1_sh[0]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst1_xxxy_inst_U5 ( .A(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U4 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst1_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst1_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst1_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst1_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst1_xxxy_inst_U2 ( .A(prince_inst_sin_x[4]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n62) );
  INV_X1 prince_inst_sbox_inst1_xxxy_inst_U1 ( .A(prince_inst_sin_x[5]), .ZN(
        prince_inst_sbox_inst1_xxxy_inst_n68) );
  XOR2_X1 prince_inst_sbox_inst1_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst1_t1_sh[1]), .B(
        prince_inst_sbox_inst1_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst1_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst1_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst1_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst1_xxyx_inst_n52), .B(
        prince_inst_sbox_inst1_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst1_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U23 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst1_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst1_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n48), .A2(prince_inst_sin_x[7]), .A3(
        prince_inst_sin_x[4]), .ZN(prince_inst_sbox_inst1_xxyx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst1_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst1_xxyx_inst_U18 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sbox_inst1_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst1_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst1_xxyx_inst_U16 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sin_x[4]), .A3(prince_inst_sbox_inst1_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst1_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst1_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n46), .A2(prince_inst_sin_x[7]), .A3(
        prince_inst_sin_x[5]), .ZN(prince_inst_sbox_inst1_xxyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst1_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst1_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst1_xxyx_inst_n54), .B(
        prince_inst_sbox_inst1_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst1_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U12 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sin_y[6]), .ZN(prince_inst_sbox_inst1_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst1_xxyx_inst_U11 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sbox_inst1_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst1_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst1_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst1_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst1_xxyx_inst_U10 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst1_xxyx_inst_U9 ( .A1(prince_inst_sin_x[7]), 
        .A2(prince_inst_sbox_inst1_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst1_xxyx_inst_U8 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sbox_inst1_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst1_xxyx_inst_U7 ( .A(prince_inst_sin_y[6]), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst1_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst1_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst1_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n53), .A2(prince_inst_sin_x[5]), .A3(
        prince_inst_sin_y[6]), .A4(prince_inst_sin_x[4]), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst1_xxyx_inst_U4 ( .A(prince_inst_sin_x[7]), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst1_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst1_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst1_xxyx_inst_n43), .A3(prince_inst_sin_x[7]), .A4(
        prince_inst_sin_y[6]), .ZN(prince_inst_sbox_inst1_xxyx_inst_n39) );
  INV_X1 prince_inst_sbox_inst1_xxyx_inst_U2 ( .A(prince_inst_sin_x[4]), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst1_xxyx_inst_U1 ( .A(prince_inst_sin_x[5]), .ZN(
        prince_inst_sbox_inst1_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst1_xyxx_inst_n74), .B(
        prince_inst_sbox_inst1_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst1_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst1_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst1_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst1_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U26 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sbox_inst1_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U25 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst1_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst1_xyxx_inst_n72), .B(
        prince_inst_sbox_inst1_s0_sh[2]), .S(
        prince_inst_sbox_inst1_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst1_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst1_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n74), .A2(prince_inst_sin_x[7]), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst1_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U21 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst1_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst1_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n74) );
  XNOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U19 ( .A(
        prince_inst_sbox_inst1_xyxx_inst_n61), .B(
        prince_inst_sbox_inst1_xyxx_inst_n60), .ZN(
        prince_inst_sbox_inst1_t1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst1_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U17 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst1_xyxx_inst_U16 ( .A(
        prince_inst_sbox_inst1_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U15 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n58) );
  NAND2_X1 prince_inst_sbox_inst1_xyxx_inst_U14 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_x[4]), .ZN(prince_inst_sbox_inst1_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U13 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst1_xyxx_inst_U12 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_xyxx_inst_n57)
         );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U11 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_x[6]), .ZN(prince_inst_sbox_inst1_xyxx_inst_n70)
         );
  NOR3_X1 prince_inst_sbox_inst1_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst1_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst1_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst1_xyxx_inst_U9 ( .A(prince_inst_sin_x[7]), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst1_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n54), .A2(prince_inst_sin_x[4]), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst1_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst1_xyxx_inst_n61), .A2(
        prince_inst_sbox_inst1_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst1_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst1_xyxx_inst_U5 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_xyxx_inst_n60), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst1_xyxx_inst_U4 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_xyxx_inst_n60)
         );
  NOR3_X1 prince_inst_sbox_inst1_xyxx_inst_U3 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sbox_inst1_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst1_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst1_xyxx_inst_U2 ( .A(prince_inst_sin_y[5]), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst1_xyxx_inst_U1 ( .A(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst1_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst1_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst1_xyyy_inst_n59), .B(
        prince_inst_sbox_inst1_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst1_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst1_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst1_xyyy_inst_U25 ( .A1(prince_inst_sin_y[6]), 
        .A2(prince_inst_sin_y[7]), .A3(prince_inst_sbox_inst1_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst1_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U24 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sbox_inst1_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U23 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sbox_inst1_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst1_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst1_xyyy_inst_U19 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sin_y[6]), .A3(prince_inst_sbox_inst1_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst1_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst1_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst1_xyyy_inst_n49), .B(
        prince_inst_sbox_inst1_xyyy_inst_n48), .S(
        prince_inst_sbox_inst1_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst1_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst1_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst1_xyyy_inst_U16 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sbox_inst1_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst1_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst1_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst1_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst1_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst1_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst1_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst1_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst1_xyyy_inst_U12 ( .A(prince_inst_sin_y[7]), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst1_xyyy_inst_U11 ( .A1(prince_inst_sin_y[7]), 
        .A2(prince_inst_sbox_inst1_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst1_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst1_t1_sh[3]), .B(
        prince_inst_sbox_inst1_xyyy_inst_n48), .S(
        prince_inst_sbox_inst1_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst1_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst1_xyyy_inst_U9 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sbox_inst1_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst1_xyyy_inst_U8 ( .A1(prince_inst_sin_x[4]), 
        .A2(prince_inst_sin_y[7]), .ZN(prince_inst_sbox_inst1_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst1_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst1_t1_sh[3]), .ZN(prince_inst_sbox_inst1_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst1_xyyy_inst_U6 ( .A1(prince_inst_sin_y[7]), 
        .A2(prince_inst_sbox_inst1_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst1_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst1_xyyy_inst_U4 ( .A(prince_inst_sin_y[5]), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst1_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst1_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst1_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst1_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst1_xyyy_inst_U2 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_x[4]), .ZN(prince_inst_sbox_inst1_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst1_xyyy_inst_U1 ( .A(prince_inst_sin_y[6]), .ZN(
        prince_inst_sbox_inst1_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst1_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U27 ( .A1(prince_inst_sin_y[4]), 
        .A2(prince_inst_sbox_inst1_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst1_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U24 ( .A1(prince_inst_sin_y[4]), 
        .A2(prince_inst_sbox_inst1_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst1_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U21 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst1_yxxx_inst_U19 ( .A(prince_inst_sin_x[7]), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst1_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst1_yxxx_inst_n52), .B(
        prince_inst_sbox_inst1_yxxx_inst_n51), .S(
        prince_inst_sbox_inst1_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst1_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n53), .A2(prince_inst_sin_x[7]), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst1_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n48), .A2(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n47), .A2(prince_inst_sin_x[7]), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U13 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sbox_inst1_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst1_yxxx_inst_n59), .B(
        prince_inst_sbox_inst1_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst1_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst1_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst1_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst1_yxxx_inst_U9 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sbox_inst1_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst1_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst1_yxxx_inst_U8 ( .A(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst1_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst1_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst1_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst1_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst1_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst1_yxxx_inst_U5 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst1_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst1_yxxx_inst_U4 ( .A(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst1_yxxx_inst_U3 ( .A(prince_inst_sin_x[5]), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst1_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst1_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst1_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst1_yxxx_inst_U1 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n67), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n66), .ZN(
        prince_inst_sbox_inst1_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst1_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n66), .A3(
        prince_inst_sbox_inst1_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst1_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst1_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n64), .A2(prince_inst_sin_x[5]), .A3(
        prince_inst_sin_y[7]), .ZN(prince_inst_sbox_inst1_yxyy_inst_n66) );
  NAND3_X1 prince_inst_sbox_inst1_yxyy_inst_U24 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n63), .A2(prince_inst_sin_y[6]), .A3(
        prince_inst_sin_y[7]), .ZN(prince_inst_sbox_inst1_yxyy_inst_n65) );
  MUX2_X1 prince_inst_sbox_inst1_yxyy_inst_U23 ( .A(
        prince_inst_sbox_inst1_yxyy_inst_n62), .B(
        prince_inst_sbox_inst1_yxyy_inst_n61), .S(prince_inst_sin_y[4]), .Z(
        prince_inst_sbox_inst1_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst1_yxyy_inst_U22 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n64), .A2(prince_inst_sin_x[5]), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst1_yxyy_inst_U21 ( .A(prince_inst_sin_x[5]), .B(
        prince_inst_sbox_inst1_yxyy_inst_n60), .S(
        prince_inst_sbox_inst1_yxyy_inst_n64), .Z(
        prince_inst_sbox_inst1_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U18 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst1_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst1_yxyy_inst_n62), .B(
        prince_inst_sbox_inst1_yxyy_inst_n54), .S(
        prince_inst_sbox_inst1_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst1_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst1_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst1_yxyy_inst_n53), .B(
        prince_inst_sbox_inst1_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst1_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst1_yxyy_inst_U15 ( .A(
        prince_inst_sbox_inst1_yxyy_inst_n67), .B(
        prince_inst_sbox_inst1_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst1_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U14 ( .A1(prince_inst_sin_y[7]), 
        .A2(prince_inst_sin_y[4]), .ZN(prince_inst_sbox_inst1_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst1_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst1_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst1_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst1_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst1_yxyy_inst_U12 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst1_yxyy_inst_U11 ( .A(
        prince_inst_sbox_inst1_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst1_yxyy_inst_U10 ( .A1(prince_inst_sin_x[5]), 
        .A2(prince_inst_sin_y[6]), .A3(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U9 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst1_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U8 ( .A1(prince_inst_sin_y[7]), 
        .A2(prince_inst_sbox_inst1_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst1_yxyy_inst_U7 ( .A1(prince_inst_sin_y[6]), 
        .A2(prince_inst_sin_x[5]), .ZN(prince_inst_sbox_inst1_yxyy_inst_n49)
         );
  OR3_X1 prince_inst_sbox_inst1_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst1_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst1_yxyy_inst_U5 ( .A(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst1_yxyy_inst_U4 ( .A(prince_inst_sin_x[5]), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst1_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst1_yxyy_inst_n64), .A2(
        prince_inst_sbox_inst1_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst1_yxyy_inst_U2 ( .A(prince_inst_sin_y[7]), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst1_yxyy_inst_U1 ( .A(prince_inst_sin_y[6]), .ZN(
        prince_inst_sbox_inst1_yxyy_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst1_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U29 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst1_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst1_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst1_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n75), .A2(prince_inst_sin_y[7]), .A3(
        prince_inst_sbox_inst1_yyxy_inst_n70), .A4(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst1_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n69), .A3(prince_inst_sin_y[5]), .A4(
        prince_inst_sbox_inst1_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst1_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst1_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst1_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst1_yyxy_inst_U23 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_x[6]), .A3(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst1_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n69), .A2(prince_inst_sin_y[5]), .A3(
        prince_inst_sin_y[7]), .ZN(prince_inst_sbox_inst1_yyxy_inst_n65) );
  NAND3_X1 prince_inst_sbox_inst1_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n75), .A2(prince_inst_sin_x[6]), .A3(
        prince_inst_sin_y[7]), .ZN(prince_inst_sbox_inst1_yyxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst1_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst1_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst1_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n61), .A2(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst1_yyxy_inst_U18 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_y[7]), .A3(prince_inst_sbox_inst1_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst1_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst1_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst1_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst1_yyxy_inst_U16 ( .A1(prince_inst_sin_y[7]), 
        .A2(prince_inst_sbox_inst1_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst1_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst1_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst1_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n58), .A3(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst1_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst1_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst1_yyxy_inst_U13 ( .A1(prince_inst_sin_y[4]), 
        .A2(prince_inst_sbox_inst1_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst1_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst1_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst1_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst1_yyxy_inst_n54), .B(
        prince_inst_sbox_inst1_yyxy_inst_n55), .S(
        prince_inst_sbox_inst1_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst1_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst1_yyxy_inst_U9 ( .A(prince_inst_sin_x[6]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n75), .A2(prince_inst_sin_y[7]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst1_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst1_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst1_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U5 ( .A1(prince_inst_sin_x[6]), 
        .A2(prince_inst_sbox_inst1_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst1_yyxy_inst_U4 ( .A(prince_inst_sin_y[5]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst1_yyxy_inst_U3 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sbox_inst1_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst1_yyxy_inst_U2 ( .A(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst1_yyxy_inst_U1 ( .A(prince_inst_sin_y[7]), .ZN(
        prince_inst_sbox_inst1_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst1_yyyx_inst_n58), .B(
        prince_inst_sbox_inst1_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst1_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst1_yyyx_inst_n56), .B(
        prince_inst_sbox_inst1_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst1_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst1_yyyx_inst_n54), .B(
        prince_inst_sbox_inst1_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst1_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst1_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst1_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst1_yyyx_inst_U21 ( .A1(prince_inst_sin_x[7]), 
        .A2(prince_inst_sbox_inst1_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst1_yyyx_inst_U20 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_y[6]), .A3(prince_inst_sbox_inst1_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst1_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst1_yyyx_inst_n50), .B(
        prince_inst_sbox_inst1_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst1_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst1_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n56), .A2(prince_inst_sin_y[6]), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst1_yyyx_inst_U17 ( .A1(prince_inst_sin_y[5]), 
        .A2(prince_inst_sin_y[4]), .A3(prince_inst_sin_y[6]), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst1_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst1_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst1_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst1_yyyx_inst_U15 ( .A1(prince_inst_sin_x[7]), 
        .A2(prince_inst_sin_y[6]), .A3(prince_inst_sbox_inst1_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst1_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst1_yyyx_inst_U14 ( .A(prince_inst_sin_y[4]), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n58), .A2(prince_inst_sin_y[5]), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst1_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst1_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U11 ( .A1(prince_inst_sin_y[4]), 
        .A2(prince_inst_sbox_inst1_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst1_yyyx_inst_U9 ( .A1(prince_inst_sin_y[4]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst1_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst1_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst1_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n45), .A2(prince_inst_sin_y[4]), .A3(
        prince_inst_sin_y[6]), .ZN(prince_inst_sbox_inst1_yyyx_inst_n54) );
  AND2_X1 prince_inst_sbox_inst1_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst1_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst1_yyyx_inst_U4 ( .A1(prince_inst_sin_x[7]), 
        .A2(prince_inst_sin_y[6]), .ZN(prince_inst_sbox_inst1_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst1_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst1_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst1_yyyx_inst_U2 ( .A(prince_inst_sin_y[5]), .ZN(
        prince_inst_sbox_inst1_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst1_yyyx_inst_U1 ( .A1(prince_inst_sin_y[4]), 
        .A2(prince_inst_sin_x[7]), .ZN(prince_inst_sbox_inst1_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s00_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[0]), .B(prince_inst_sbox_inst1_s0_sh[0]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s01_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[1]), .B(prince_inst_sbox_inst1_s0_sh[1]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s02_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[2]), .B(prince_inst_sbox_inst1_s0_sh[2]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s03_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[3]), .B(prince_inst_sbox_inst1_s0_sh[3]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s04_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[4]), .B(prince_inst_sbox_inst1_s0_sh[4]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s05_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[5]), .B(prince_inst_sbox_inst1_s0_sh[5]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s06_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[6]), .B(prince_inst_sbox_inst1_s0_sh[6]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s07_U1 ( .A(
        prince_inst_sbox_inst1_t0_sh[7]), .B(prince_inst_sbox_inst1_s0_sh[7]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s10_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[0]), .B(prince_inst_sbox_inst1_s1_sh[0]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s11_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[1]), .B(prince_inst_sbox_inst1_s1_sh[1]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s12_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[2]), .B(prince_inst_sbox_inst1_s1_sh[2]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s13_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[3]), .B(prince_inst_sbox_inst1_s1_sh[3]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s14_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[4]), .B(prince_inst_sbox_inst1_s1_sh[4]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s15_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[5]), .B(prince_inst_sbox_inst1_s1_sh[5]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s16_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[6]), .B(prince_inst_sbox_inst1_s1_sh[6]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s17_U1 ( .A(
        prince_inst_sbox_inst1_t1_sh[7]), .B(prince_inst_sbox_inst1_s1_sh[7]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s20_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[0]), .B(prince_inst_sbox_inst1_s2_sh[0]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s21_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[1]), .B(prince_inst_sbox_inst1_s2_sh[1]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s22_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[2]), .B(prince_inst_sbox_inst1_s2_sh[2]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s23_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[3]), .B(prince_inst_sbox_inst1_s2_sh[3]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s24_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[4]), .B(prince_inst_sbox_inst1_s2_sh[4]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s25_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[5]), .B(prince_inst_sbox_inst1_s2_sh[5]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s26_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[6]), .B(prince_inst_sbox_inst1_s2_sh[6]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s27_U1 ( .A(
        prince_inst_sbox_inst1_t2_sh[7]), .B(prince_inst_sbox_inst1_s2_sh[7]), 
        .S(prince_inst_sbox_inst1_n9), .Z(prince_inst_sbox_inst1_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s30_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[0]), .B(prince_inst_sbox_inst1_s3_sh[0]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s31_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[1]), .B(prince_inst_sbox_inst1_s3_sh[1]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s32_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[2]), .B(prince_inst_sbox_inst1_s3_sh[2]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s33_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[3]), .B(prince_inst_sbox_inst1_s3_sh[3]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s34_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[4]), .B(prince_inst_sbox_inst1_s3_sh[4]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s35_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[5]), .B(prince_inst_sbox_inst1_s3_sh[5]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s36_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[6]), .B(prince_inst_sbox_inst1_s3_sh[6]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst1_mux_s37_U1 ( .A(
        prince_inst_sbox_inst1_t3_sh[7]), .B(prince_inst_sbox_inst1_s3_sh[7]), 
        .S(prince_inst_sbox_inst1_n10), .Z(prince_inst_sbox_inst1_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk0_U1 ( .A(r[16]), .B(
        prince_inst_sbox_inst1_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk1_U1 ( .A(r[17]), .B(
        prince_inst_sbox_inst1_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk2_U1 ( .A(r[18]), .B(
        prince_inst_sbox_inst1_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk3_U1 ( .A(r[19]), .B(
        prince_inst_sbox_inst1_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk4_U1 ( .A(r[16]), .B(
        prince_inst_sbox_inst1_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk5_U1 ( .A(r[17]), .B(
        prince_inst_sbox_inst1_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk6_U1 ( .A(r[18]), .B(
        prince_inst_sbox_inst1_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_msk7_U1 ( .A(r[19]), .B(
        prince_inst_sbox_inst1_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst1_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst1_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst1_c_inst0_ax_n5), .ZN(prince_inst_sout_x[4]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst1_c_inst0_y[1]), .B(
        prince_inst_sbox_inst1_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst1_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst1_c_inst0_y[2]), .B(
        prince_inst_sbox_inst1_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst1_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst1_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst1_c_inst0_ay_n5), .ZN(final_y[36]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst1_c_inst0_y[5]), .B(
        prince_inst_sbox_inst1_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst1_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst1_c_inst0_y[6]), .B(
        prince_inst_sbox_inst1_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst1_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk0_U1 ( .A(r[20]), .B(
        prince_inst_sbox_inst1_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk1_U1 ( .A(r[21]), .B(
        prince_inst_sbox_inst1_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk2_U1 ( .A(r[22]), .B(
        prince_inst_sbox_inst1_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk3_U1 ( .A(r[23]), .B(
        prince_inst_sbox_inst1_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk4_U1 ( .A(r[20]), .B(
        prince_inst_sbox_inst1_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk5_U1 ( .A(r[21]), .B(
        prince_inst_sbox_inst1_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk6_U1 ( .A(r[22]), .B(
        prince_inst_sbox_inst1_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_msk7_U1 ( .A(r[23]), .B(
        prince_inst_sbox_inst1_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst1_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst1_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst1_c_inst1_ax_n5), .ZN(prince_inst_sout_x[5]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst1_c_inst1_y[1]), .B(
        prince_inst_sbox_inst1_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst1_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst1_c_inst1_y[2]), .B(
        prince_inst_sbox_inst1_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst1_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst1_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst1_c_inst1_ay_n5), .ZN(final_y[37]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst1_c_inst1_y[5]), .B(
        prince_inst_sbox_inst1_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst1_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst1_c_inst1_y[6]), .B(
        prince_inst_sbox_inst1_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst1_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk0_U1 ( .A(r[24]), .B(
        prince_inst_sbox_inst1_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk1_U1 ( .A(r[25]), .B(
        prince_inst_sbox_inst1_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk2_U1 ( .A(r[26]), .B(
        prince_inst_sbox_inst1_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk3_U1 ( .A(r[27]), .B(
        prince_inst_sbox_inst1_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk4_U1 ( .A(r[24]), .B(
        prince_inst_sbox_inst1_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk5_U1 ( .A(r[25]), .B(
        prince_inst_sbox_inst1_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk6_U1 ( .A(r[26]), .B(
        prince_inst_sbox_inst1_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_msk7_U1 ( .A(r[27]), .B(
        prince_inst_sbox_inst1_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst1_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst1_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst1_c_inst2_ax_n5), .ZN(prince_inst_sout_x[6]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst1_c_inst2_y[1]), .B(
        prince_inst_sbox_inst1_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst1_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst1_c_inst2_y[2]), .B(
        prince_inst_sbox_inst1_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst1_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst1_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst1_c_inst2_ay_n5), .ZN(final_y[38]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst1_c_inst2_y[5]), .B(
        prince_inst_sbox_inst1_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst1_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst1_c_inst2_y[6]), .B(
        prince_inst_sbox_inst1_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst1_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk0_U1 ( .A(r[28]), .B(
        prince_inst_sbox_inst1_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk1_U1 ( .A(r[29]), .B(
        prince_inst_sbox_inst1_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk2_U1 ( .A(r[30]), .B(
        prince_inst_sbox_inst1_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk3_U1 ( .A(r[31]), .B(
        prince_inst_sbox_inst1_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk4_U1 ( .A(r[28]), .B(
        prince_inst_sbox_inst1_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk5_U1 ( .A(r[29]), .B(
        prince_inst_sbox_inst1_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk6_U1 ( .A(r[30]), .B(
        prince_inst_sbox_inst1_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_msk7_U1 ( .A(r[31]), .B(
        prince_inst_sbox_inst1_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst1_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst1_n7), .A3(
        prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst1_n12), .A2(prince_inst_sbox_inst1_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst1_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst1_n12), .ZN(
        prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst1_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst1_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst1_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst1_c_inst3_ax_n5), .ZN(prince_inst_sout_x[7]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst1_c_inst3_y[1]), .B(
        prince_inst_sbox_inst1_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst1_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst1_c_inst3_y[2]), .B(
        prince_inst_sbox_inst1_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst1_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst1_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst1_c_inst3_ay_n5), .ZN(final_y[39]) );
  XNOR2_X1 prince_inst_sbox_inst1_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst1_c_inst3_y[5]), .B(
        prince_inst_sbox_inst1_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst1_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst1_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst1_c_inst3_y[6]), .B(
        prince_inst_sbox_inst1_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst1_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst2_U7 ( .A(prince_inst_sbox_inst2_n12), .ZN(
        prince_inst_sbox_inst2_n11) );
  INV_X1 prince_inst_sbox_inst2_U6 ( .A(prince_inst_n26), .ZN(
        prince_inst_sbox_inst2_n10) );
  INV_X1 prince_inst_sbox_inst2_U5 ( .A(prince_inst_sbox_inst2_n10), .ZN(
        prince_inst_sbox_inst2_n8) );
  INV_X1 prince_inst_sbox_inst2_U4 ( .A(prince_inst_sbox_inst2_n10), .ZN(
        prince_inst_sbox_inst2_n9) );
  INV_X1 prince_inst_sbox_inst2_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst2_n12) );
  INV_X1 prince_inst_sbox_inst2_U2 ( .A(rst), .ZN(prince_inst_sbox_inst2_n7)
         );
  INV_X2 prince_inst_sbox_inst2_U1 ( .A(prince_inst_sbox_inst2_n7), .ZN(
        prince_inst_sbox_inst2_n6) );
  NAND3_X1 prince_inst_sbox_inst2_xxxy_inst_U28 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n70), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n69), .A3(prince_inst_sin_x[8]), .ZN(
        prince_inst_sbox_inst2_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n67), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n69) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U26 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n70) );
  NAND3_X1 prince_inst_sbox_inst2_xxxy_inst_U25 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n65), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n64), .A3(
        prince_inst_sbox_inst2_xxxy_inst_n63), .ZN(
        prince_inst_sbox_inst2_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst2_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n68), .A2(prince_inst_sin_x[10]), 
        .A3(prince_inst_sin_x[8]), .A4(prince_inst_sin_y[11]), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n63) );
  NAND3_X1 prince_inst_sbox_inst2_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n62), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n61), .A3(prince_inst_sin_x[10]), 
        .ZN(prince_inst_sbox_inst2_xxxy_inst_n64) );
  NAND4_X1 prince_inst_sbox_inst2_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n67), .A3(
        prince_inst_sbox_inst2_xxxy_inst_n61), .A4(prince_inst_sin_x[8]), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n65) );
  XOR2_X1 prince_inst_sbox_inst2_xxxy_inst_U21 ( .A(
        prince_inst_sbox_inst2_xxxy_inst_n59), .B(prince_inst_sin_y[11]), .Z(
        prince_inst_sbox_inst2_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U20 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U19 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n58) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U18 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst2_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst2_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n66), .A2(prince_inst_sin_x[10]), 
        .ZN(prince_inst_sbox_inst2_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst2_xxxy_inst_U16 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sin_y[11]), .A3(prince_inst_sbox_inst2_xxxy_inst_n68), 
        .ZN(prince_inst_sbox_inst2_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst2_xxxy_inst_U15 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst2_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst2_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst2_xxxy_inst_U14 ( .A(prince_inst_sin_x[8]), .B(
        prince_inst_sbox_inst2_xxxy_inst_n61), .S(
        prince_inst_sbox_inst2_xxxy_inst_n67), .Z(
        prince_inst_sbox_inst2_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst2_xxxy_inst_U13 ( .A(prince_inst_sin_y[11]), 
        .ZN(prince_inst_sbox_inst2_xxxy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U12 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n61), .A2(prince_inst_sin_x[8]), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U11 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst2_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst2_xxxy_inst_U10 ( .A(
        prince_inst_sbox_inst2_xxxy_inst_n60), .B(
        prince_inst_sbox_inst2_xxxy_inst_n53), .S(
        prince_inst_sbox_inst2_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst2_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U9 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sbox_inst2_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U8 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n61), .A2(prince_inst_sin_y[11]), 
        .ZN(prince_inst_sbox_inst2_xxxy_inst_n66) );
  INV_X1 prince_inst_sbox_inst2_xxxy_inst_U7 ( .A(
        prince_inst_sbox_inst2_xxxy_inst_n68), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst2_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst2_t1_sh[0]), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst2_xxxy_inst_U5 ( .A(prince_inst_sin_x[10]), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U4 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst2_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst2_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst2_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst2_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst2_xxxy_inst_U2 ( .A(prince_inst_sin_x[8]), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n62) );
  INV_X1 prince_inst_sbox_inst2_xxxy_inst_U1 ( .A(prince_inst_sin_x[9]), .ZN(
        prince_inst_sbox_inst2_xxxy_inst_n68) );
  XOR2_X1 prince_inst_sbox_inst2_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst2_t1_sh[1]), .B(
        prince_inst_sbox_inst2_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst2_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst2_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst2_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst2_xxyx_inst_n52), .B(
        prince_inst_sbox_inst2_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst2_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U23 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst2_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst2_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n48), .A2(prince_inst_sin_x[11]), 
        .A3(prince_inst_sin_x[8]), .ZN(prince_inst_sbox_inst2_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n45), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst2_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst2_xxyx_inst_U18 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n46), .A2(prince_inst_sin_x[11]), 
        .A3(prince_inst_sin_x[9]), .ZN(prince_inst_sbox_inst2_xxyx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst2_t2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst2_xxyx_inst_U16 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sin_x[8]), .A3(prince_inst_sbox_inst2_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst2_xxyx_inst_n44) );
  OR2_X1 prince_inst_sbox_inst2_xxyx_inst_U15 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sbox_inst2_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst2_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst2_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst2_xxyx_inst_n54), .B(
        prince_inst_sbox_inst2_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst2_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U12 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sin_y[10]), .ZN(prince_inst_sbox_inst2_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst2_xxyx_inst_U11 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sbox_inst2_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst2_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst2_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst2_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst2_xxyx_inst_U10 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst2_xxyx_inst_U9 ( .A1(prince_inst_sin_x[11]), 
        .A2(prince_inst_sbox_inst2_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst2_xxyx_inst_U8 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sbox_inst2_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst2_xxyx_inst_U7 ( .A(prince_inst_sin_y[10]), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst2_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst2_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst2_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n53), .A2(prince_inst_sin_x[9]), .A3(
        prince_inst_sin_y[10]), .A4(prince_inst_sin_x[8]), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst2_xxyx_inst_U4 ( .A(prince_inst_sin_x[11]), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst2_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst2_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst2_xxyx_inst_n43), .A3(prince_inst_sin_x[11]), 
        .A4(prince_inst_sin_y[10]), .ZN(prince_inst_sbox_inst2_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst2_xxyx_inst_U2 ( .A(prince_inst_sin_x[8]), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst2_xxyx_inst_U1 ( .A(prince_inst_sin_x[9]), .ZN(
        prince_inst_sbox_inst2_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst2_xyxx_inst_n74), .B(
        prince_inst_sbox_inst2_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst2_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst2_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst2_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst2_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U26 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sbox_inst2_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U25 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst2_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst2_xyxx_inst_n72), .B(
        prince_inst_sbox_inst2_s0_sh[2]), .S(
        prince_inst_sbox_inst2_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst2_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst2_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n74), .A2(prince_inst_sin_x[11]), 
        .ZN(prince_inst_sbox_inst2_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst2_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U21 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst2_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst2_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst2_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst2_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst2_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst2_xyxx_inst_U15 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_x[8]), .ZN(prince_inst_sbox_inst2_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst2_xyxx_inst_U13 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U12 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_x[10]), .ZN(prince_inst_sbox_inst2_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst2_xyxx_inst_n58), .B(
        prince_inst_sbox_inst2_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst2_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst2_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst2_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst2_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst2_xyxx_inst_U9 ( .A(prince_inst_sin_x[11]), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst2_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n54), .A2(prince_inst_sin_x[8]), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst2_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst2_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst2_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst2_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst2_xyxx_inst_U5 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst2_xyxx_inst_U4 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst2_xyxx_inst_U3 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sbox_inst2_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst2_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst2_xyxx_inst_U2 ( .A(prince_inst_sin_y[9]), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst2_xyxx_inst_U1 ( .A(prince_inst_sin_x[10]), .ZN(
        prince_inst_sbox_inst2_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst2_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst2_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst2_xyyy_inst_n59), .B(
        prince_inst_sbox_inst2_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst2_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst2_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst2_xyyy_inst_U25 ( .A1(prince_inst_sin_y[10]), 
        .A2(prince_inst_sin_y[11]), .A3(prince_inst_sbox_inst2_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst2_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U24 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sbox_inst2_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U23 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sbox_inst2_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst2_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst2_xyyy_inst_U19 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sin_y[10]), .A3(prince_inst_sbox_inst2_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst2_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst2_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst2_xyyy_inst_n49), .B(
        prince_inst_sbox_inst2_xyyy_inst_n48), .S(
        prince_inst_sbox_inst2_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst2_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst2_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst2_xyyy_inst_U16 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sbox_inst2_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst2_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst2_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst2_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst2_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst2_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst2_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst2_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst2_xyyy_inst_U12 ( .A(prince_inst_sin_y[11]), 
        .ZN(prince_inst_sbox_inst2_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst2_xyyy_inst_U11 ( .A1(prince_inst_sin_y[11]), 
        .A2(prince_inst_sbox_inst2_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst2_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst2_t1_sh[3]), .B(
        prince_inst_sbox_inst2_xyyy_inst_n48), .S(
        prince_inst_sbox_inst2_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst2_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst2_xyyy_inst_U9 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sbox_inst2_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst2_xyyy_inst_U8 ( .A1(prince_inst_sin_x[8]), 
        .A2(prince_inst_sin_y[11]), .ZN(prince_inst_sbox_inst2_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst2_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst2_t1_sh[3]), .ZN(prince_inst_sbox_inst2_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst2_xyyy_inst_U6 ( .A1(prince_inst_sin_y[11]), 
        .A2(prince_inst_sbox_inst2_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst2_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst2_xyyy_inst_U4 ( .A(prince_inst_sin_y[9]), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst2_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst2_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst2_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst2_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst2_xyyy_inst_U2 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_x[8]), .ZN(prince_inst_sbox_inst2_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst2_xyyy_inst_U1 ( .A(prince_inst_sin_y[10]), .ZN(
        prince_inst_sbox_inst2_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst2_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U27 ( .A1(prince_inst_sin_y[8]), 
        .A2(prince_inst_sbox_inst2_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst2_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U24 ( .A1(prince_inst_sin_y[8]), 
        .A2(prince_inst_sbox_inst2_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst2_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U21 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst2_yxxx_inst_U19 ( .A(prince_inst_sin_x[11]), 
        .ZN(prince_inst_sbox_inst2_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst2_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst2_yxxx_inst_n52), .B(
        prince_inst_sbox_inst2_yxxx_inst_n51), .S(
        prince_inst_sbox_inst2_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst2_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n53), .A2(prince_inst_sin_x[11]), 
        .ZN(prince_inst_sbox_inst2_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst2_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n48), .A2(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n47), .A2(prince_inst_sin_x[11]), 
        .ZN(prince_inst_sbox_inst2_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U13 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sbox_inst2_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst2_yxxx_inst_n59), .B(
        prince_inst_sbox_inst2_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst2_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst2_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst2_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst2_yxxx_inst_U9 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sbox_inst2_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst2_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst2_yxxx_inst_U8 ( .A(prince_inst_sin_x[10]), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst2_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst2_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst2_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst2_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst2_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst2_yxxx_inst_U5 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst2_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst2_yxxx_inst_U4 ( .A(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst2_yxxx_inst_U3 ( .A(prince_inst_sin_x[9]), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst2_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst2_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst2_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst2_yxxx_inst_U1 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n67), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n66), .ZN(
        prince_inst_sbox_inst2_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst2_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n66), .A3(
        prince_inst_sbox_inst2_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst2_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst2_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n64), .A2(prince_inst_sin_x[9]), .A3(
        prince_inst_sin_y[11]), .ZN(prince_inst_sbox_inst2_yxyy_inst_n66) );
  NAND3_X1 prince_inst_sbox_inst2_yxyy_inst_U24 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n63), .A2(prince_inst_sin_y[10]), 
        .A3(prince_inst_sin_y[11]), .ZN(prince_inst_sbox_inst2_yxyy_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst2_yxyy_inst_U23 ( .A(
        prince_inst_sbox_inst2_yxyy_inst_n62), .B(
        prince_inst_sbox_inst2_yxyy_inst_n61), .S(prince_inst_sin_y[8]), .Z(
        prince_inst_sbox_inst2_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst2_yxyy_inst_U22 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n64), .A2(prince_inst_sin_x[9]), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst2_yxyy_inst_U21 ( .A(prince_inst_sin_x[9]), .B(
        prince_inst_sbox_inst2_yxyy_inst_n60), .S(
        prince_inst_sbox_inst2_yxyy_inst_n64), .Z(
        prince_inst_sbox_inst2_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U18 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst2_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst2_yxyy_inst_n62), .B(
        prince_inst_sbox_inst2_yxyy_inst_n54), .S(
        prince_inst_sbox_inst2_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst2_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst2_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst2_yxyy_inst_n53), .B(
        prince_inst_sbox_inst2_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst2_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst2_yxyy_inst_U15 ( .A(
        prince_inst_sbox_inst2_yxyy_inst_n67), .B(
        prince_inst_sbox_inst2_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst2_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U14 ( .A1(prince_inst_sin_y[11]), 
        .A2(prince_inst_sin_y[8]), .ZN(prince_inst_sbox_inst2_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst2_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst2_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst2_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst2_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst2_yxyy_inst_U12 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst2_yxyy_inst_U11 ( .A(
        prince_inst_sbox_inst2_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst2_yxyy_inst_U10 ( .A1(prince_inst_sin_x[9]), 
        .A2(prince_inst_sin_y[10]), .A3(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U9 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst2_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U8 ( .A1(prince_inst_sin_y[11]), 
        .A2(prince_inst_sbox_inst2_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst2_yxyy_inst_U7 ( .A1(prince_inst_sin_y[10]), 
        .A2(prince_inst_sin_x[9]), .ZN(prince_inst_sbox_inst2_yxyy_inst_n49)
         );
  OR3_X1 prince_inst_sbox_inst2_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst2_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst2_yxyy_inst_U5 ( .A(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst2_yxyy_inst_U4 ( .A(prince_inst_sin_x[9]), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst2_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst2_yxyy_inst_n64), .A2(
        prince_inst_sbox_inst2_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst2_yxyy_inst_U2 ( .A(prince_inst_sin_y[11]), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst2_yxyy_inst_U1 ( .A(prince_inst_sin_y[10]), .ZN(
        prince_inst_sbox_inst2_yxyy_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst2_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U29 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst2_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst2_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst2_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n75), .A2(prince_inst_sin_y[11]), 
        .A3(prince_inst_sbox_inst2_yyxy_inst_n70), .A4(prince_inst_sin_x[10]), 
        .ZN(prince_inst_sbox_inst2_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst2_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n69), .A3(prince_inst_sin_y[9]), .A4(
        prince_inst_sbox_inst2_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst2_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst2_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst2_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst2_yyxy_inst_U23 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_x[10]), .A3(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst2_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n69), .A2(prince_inst_sin_y[9]), .A3(
        prince_inst_sin_y[11]), .ZN(prince_inst_sbox_inst2_yyxy_inst_n65) );
  NAND3_X1 prince_inst_sbox_inst2_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n75), .A2(prince_inst_sin_x[10]), 
        .A3(prince_inst_sin_y[11]), .ZN(prince_inst_sbox_inst2_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst2_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst2_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst2_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n61), .A2(prince_inst_sin_x[10]), 
        .ZN(prince_inst_sbox_inst2_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst2_yyxy_inst_U18 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_y[11]), .A3(prince_inst_sbox_inst2_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst2_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst2_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst2_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst2_yyxy_inst_U16 ( .A1(prince_inst_sin_y[11]), 
        .A2(prince_inst_sbox_inst2_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst2_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst2_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst2_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n58), .A3(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst2_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst2_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst2_yyxy_inst_U13 ( .A1(prince_inst_sin_y[8]), 
        .A2(prince_inst_sbox_inst2_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst2_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst2_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst2_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst2_yyxy_inst_n54), .B(
        prince_inst_sbox_inst2_yyxy_inst_n55), .S(
        prince_inst_sbox_inst2_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst2_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst2_yyxy_inst_U9 ( .A(prince_inst_sin_x[10]), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n75), .A2(prince_inst_sin_y[11]), 
        .ZN(prince_inst_sbox_inst2_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst2_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst2_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst2_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U5 ( .A1(prince_inst_sin_x[10]), 
        .A2(prince_inst_sbox_inst2_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst2_yyxy_inst_U4 ( .A(prince_inst_sin_y[9]), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst2_yyxy_inst_U3 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sbox_inst2_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst2_yyxy_inst_U2 ( .A(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst2_yyxy_inst_U1 ( .A(prince_inst_sin_y[11]), .ZN(
        prince_inst_sbox_inst2_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst2_yyyx_inst_n58), .B(
        prince_inst_sbox_inst2_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst2_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst2_yyyx_inst_n56), .B(
        prince_inst_sbox_inst2_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst2_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst2_yyyx_inst_n54), .B(
        prince_inst_sbox_inst2_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst2_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst2_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst2_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst2_yyyx_inst_U21 ( .A1(prince_inst_sin_x[11]), 
        .A2(prince_inst_sbox_inst2_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst2_yyyx_inst_U20 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_y[10]), .A3(prince_inst_sbox_inst2_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst2_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst2_yyyx_inst_n50), .B(
        prince_inst_sbox_inst2_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst2_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst2_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n56), .A2(prince_inst_sin_y[10]), 
        .ZN(prince_inst_sbox_inst2_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst2_yyyx_inst_U17 ( .A1(prince_inst_sin_y[9]), 
        .A2(prince_inst_sin_y[8]), .A3(prince_inst_sin_y[10]), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst2_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst2_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst2_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst2_yyyx_inst_U15 ( .A1(prince_inst_sin_x[11]), 
        .A2(prince_inst_sin_y[10]), .A3(prince_inst_sbox_inst2_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst2_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst2_yyyx_inst_U14 ( .A(prince_inst_sin_y[8]), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n58), .A2(prince_inst_sin_y[9]), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst2_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst2_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U11 ( .A1(prince_inst_sin_y[8]), 
        .A2(prince_inst_sbox_inst2_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst2_yyyx_inst_U9 ( .A1(prince_inst_sin_y[8]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst2_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst2_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst2_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n45), .A2(prince_inst_sin_y[8]), .A3(
        prince_inst_sin_y[10]), .ZN(prince_inst_sbox_inst2_yyyx_inst_n54) );
  AND2_X1 prince_inst_sbox_inst2_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst2_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst2_yyyx_inst_U4 ( .A1(prince_inst_sin_x[11]), 
        .A2(prince_inst_sin_y[10]), .ZN(prince_inst_sbox_inst2_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst2_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst2_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst2_yyyx_inst_U2 ( .A(prince_inst_sin_y[9]), .ZN(
        prince_inst_sbox_inst2_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst2_yyyx_inst_U1 ( .A1(prince_inst_sin_y[8]), 
        .A2(prince_inst_sin_x[11]), .ZN(prince_inst_sbox_inst2_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s00_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[0]), .B(prince_inst_sbox_inst2_s0_sh[0]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s01_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[1]), .B(prince_inst_sbox_inst2_s0_sh[1]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s02_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[2]), .B(prince_inst_sbox_inst2_s0_sh[2]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s03_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[3]), .B(prince_inst_sbox_inst2_s0_sh[3]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s04_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[4]), .B(prince_inst_sbox_inst2_s0_sh[4]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s05_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[5]), .B(prince_inst_sbox_inst2_s0_sh[5]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s06_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[6]), .B(prince_inst_sbox_inst2_s0_sh[6]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s07_U1 ( .A(
        prince_inst_sbox_inst2_t0_sh[7]), .B(prince_inst_sbox_inst2_s0_sh[7]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s10_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[0]), .B(prince_inst_sbox_inst2_s1_sh[0]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s11_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[1]), .B(prince_inst_sbox_inst2_s1_sh[1]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s12_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[2]), .B(prince_inst_sbox_inst2_s1_sh[2]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s13_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[3]), .B(prince_inst_sbox_inst2_s1_sh[3]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s14_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[4]), .B(prince_inst_sbox_inst2_s1_sh[4]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s15_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[5]), .B(prince_inst_sbox_inst2_s1_sh[5]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s16_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[6]), .B(prince_inst_sbox_inst2_s1_sh[6]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s17_U1 ( .A(
        prince_inst_sbox_inst2_t1_sh[7]), .B(prince_inst_sbox_inst2_s1_sh[7]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s20_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[0]), .B(prince_inst_sbox_inst2_s2_sh[0]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s21_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[1]), .B(prince_inst_sbox_inst2_s2_sh[1]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s22_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[2]), .B(prince_inst_sbox_inst2_s2_sh[2]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s23_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[3]), .B(prince_inst_sbox_inst2_s2_sh[3]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s24_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[4]), .B(prince_inst_sbox_inst2_s2_sh[4]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s25_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[5]), .B(prince_inst_sbox_inst2_s2_sh[5]), 
        .S(prince_inst_sbox_inst2_n8), .Z(prince_inst_sbox_inst2_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s26_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[6]), .B(prince_inst_sbox_inst2_s2_sh[6]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s27_U1 ( .A(
        prince_inst_sbox_inst2_t2_sh[7]), .B(prince_inst_sbox_inst2_s2_sh[7]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s30_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[0]), .B(prince_inst_sbox_inst2_s3_sh[0]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s31_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[1]), .B(prince_inst_sbox_inst2_s3_sh[1]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s32_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[2]), .B(prince_inst_sbox_inst2_s3_sh[2]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s33_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[3]), .B(prince_inst_sbox_inst2_s3_sh[3]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s34_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[4]), .B(prince_inst_sbox_inst2_s3_sh[4]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s35_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[5]), .B(prince_inst_sbox_inst2_s3_sh[5]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s36_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[6]), .B(prince_inst_sbox_inst2_s3_sh[6]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst2_mux_s37_U1 ( .A(
        prince_inst_sbox_inst2_t3_sh[7]), .B(prince_inst_sbox_inst2_s3_sh[7]), 
        .S(prince_inst_sbox_inst2_n9), .Z(prince_inst_sbox_inst2_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk0_U1 ( .A(r[32]), .B(
        prince_inst_sbox_inst2_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk1_U1 ( .A(r[33]), .B(
        prince_inst_sbox_inst2_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk2_U1 ( .A(r[34]), .B(
        prince_inst_sbox_inst2_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk3_U1 ( .A(r[35]), .B(
        prince_inst_sbox_inst2_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk4_U1 ( .A(r[32]), .B(
        prince_inst_sbox_inst2_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk5_U1 ( .A(r[33]), .B(
        prince_inst_sbox_inst2_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk6_U1 ( .A(r[34]), .B(
        prince_inst_sbox_inst2_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_msk7_U1 ( .A(r[35]), .B(
        prince_inst_sbox_inst2_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst2_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst2_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst2_c_inst0_ax_n5), .ZN(prince_inst_sout_x[8]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst2_c_inst0_y[1]), .B(
        prince_inst_sbox_inst2_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst2_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst2_c_inst0_y[2]), .B(
        prince_inst_sbox_inst2_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst2_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst2_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst2_c_inst0_ay_n5), .ZN(final_y[24]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst2_c_inst0_y[5]), .B(
        prince_inst_sbox_inst2_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst2_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst2_c_inst0_y[6]), .B(
        prince_inst_sbox_inst2_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst2_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk0_U1 ( .A(r[36]), .B(
        prince_inst_sbox_inst2_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk1_U1 ( .A(r[37]), .B(
        prince_inst_sbox_inst2_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk2_U1 ( .A(r[38]), .B(
        prince_inst_sbox_inst2_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk3_U1 ( .A(r[39]), .B(
        prince_inst_sbox_inst2_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk4_U1 ( .A(r[36]), .B(
        prince_inst_sbox_inst2_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk5_U1 ( .A(r[37]), .B(
        prince_inst_sbox_inst2_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk6_U1 ( .A(r[38]), .B(
        prince_inst_sbox_inst2_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_msk7_U1 ( .A(r[39]), .B(
        prince_inst_sbox_inst2_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst2_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst2_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst2_c_inst1_ax_n5), .ZN(prince_inst_sout_x[9]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst2_c_inst1_y[1]), .B(
        prince_inst_sbox_inst2_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst2_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst2_c_inst1_y[2]), .B(
        prince_inst_sbox_inst2_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst2_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst2_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst2_c_inst1_ay_n5), .ZN(final_y[25]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst2_c_inst1_y[5]), .B(
        prince_inst_sbox_inst2_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst2_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst2_c_inst1_y[6]), .B(
        prince_inst_sbox_inst2_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst2_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk0_U1 ( .A(r[40]), .B(
        prince_inst_sbox_inst2_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk1_U1 ( .A(r[41]), .B(
        prince_inst_sbox_inst2_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk2_U1 ( .A(r[42]), .B(
        prince_inst_sbox_inst2_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk3_U1 ( .A(r[43]), .B(
        prince_inst_sbox_inst2_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk4_U1 ( .A(r[40]), .B(
        prince_inst_sbox_inst2_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk5_U1 ( .A(r[41]), .B(
        prince_inst_sbox_inst2_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk6_U1 ( .A(r[42]), .B(
        prince_inst_sbox_inst2_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_msk7_U1 ( .A(r[43]), .B(
        prince_inst_sbox_inst2_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst2_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst2_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst2_c_inst2_ax_n5), .ZN(prince_inst_sout_x[10]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst2_c_inst2_y[1]), .B(
        prince_inst_sbox_inst2_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst2_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst2_c_inst2_y[2]), .B(
        prince_inst_sbox_inst2_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst2_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst2_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst2_c_inst2_ay_n5), .ZN(final_y[26]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst2_c_inst2_y[5]), .B(
        prince_inst_sbox_inst2_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst2_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst2_c_inst2_y[6]), .B(
        prince_inst_sbox_inst2_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst2_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk0_U1 ( .A(r[44]), .B(
        prince_inst_sbox_inst2_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk1_U1 ( .A(r[45]), .B(
        prince_inst_sbox_inst2_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk2_U1 ( .A(r[46]), .B(
        prince_inst_sbox_inst2_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk3_U1 ( .A(r[47]), .B(
        prince_inst_sbox_inst2_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk4_U1 ( .A(r[44]), .B(
        prince_inst_sbox_inst2_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk5_U1 ( .A(r[45]), .B(
        prince_inst_sbox_inst2_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk6_U1 ( .A(r[46]), .B(
        prince_inst_sbox_inst2_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_msk7_U1 ( .A(r[47]), .B(
        prince_inst_sbox_inst2_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst2_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst2_n6), .A3(
        prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst2_n11), .A2(prince_inst_sbox_inst2_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst2_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst2_n11), .ZN(
        prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst2_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst2_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst2_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst2_c_inst3_ax_n5), .ZN(prince_inst_sout_x[11]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst2_c_inst3_y[1]), .B(
        prince_inst_sbox_inst2_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst2_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst2_c_inst3_y[2]), .B(
        prince_inst_sbox_inst2_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst2_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst2_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst2_c_inst3_ay_n5), .ZN(final_y[27]) );
  XNOR2_X1 prince_inst_sbox_inst2_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst2_c_inst3_y[5]), .B(
        prince_inst_sbox_inst2_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst2_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst2_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst2_c_inst3_y[6]), .B(
        prince_inst_sbox_inst2_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst2_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst3_U7 ( .A(prince_inst_sbox_inst3_n12), .ZN(
        prince_inst_sbox_inst3_n11) );
  INV_X1 prince_inst_sbox_inst3_U6 ( .A(prince_inst_n27), .ZN(
        prince_inst_sbox_inst3_n10) );
  INV_X1 prince_inst_sbox_inst3_U5 ( .A(prince_inst_sbox_inst3_n10), .ZN(
        prince_inst_sbox_inst3_n8) );
  INV_X1 prince_inst_sbox_inst3_U4 ( .A(prince_inst_sbox_inst3_n10), .ZN(
        prince_inst_sbox_inst3_n9) );
  INV_X1 prince_inst_sbox_inst3_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst3_n12) );
  INV_X1 prince_inst_sbox_inst3_U2 ( .A(rst), .ZN(prince_inst_sbox_inst3_n7)
         );
  INV_X2 prince_inst_sbox_inst3_U1 ( .A(prince_inst_sbox_inst3_n7), .ZN(
        prince_inst_sbox_inst3_n6) );
  NAND3_X1 prince_inst_sbox_inst3_xxxy_inst_U28 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n70), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n69), .A3(prince_inst_sin_x[12]), 
        .ZN(prince_inst_sbox_inst3_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n67), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n69) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U26 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n70) );
  NAND3_X1 prince_inst_sbox_inst3_xxxy_inst_U25 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n65), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n64), .A3(
        prince_inst_sbox_inst3_xxxy_inst_n63), .ZN(
        prince_inst_sbox_inst3_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst3_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n68), .A2(prince_inst_sin_x[14]), 
        .A3(prince_inst_sin_x[12]), .A4(prince_inst_sin_y[15]), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n63) );
  NAND3_X1 prince_inst_sbox_inst3_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n62), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n61), .A3(prince_inst_sin_x[14]), 
        .ZN(prince_inst_sbox_inst3_xxxy_inst_n64) );
  NAND4_X1 prince_inst_sbox_inst3_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n67), .A3(
        prince_inst_sbox_inst3_xxxy_inst_n61), .A4(prince_inst_sin_x[12]), 
        .ZN(prince_inst_sbox_inst3_xxxy_inst_n65) );
  XOR2_X1 prince_inst_sbox_inst3_xxxy_inst_U21 ( .A(
        prince_inst_sbox_inst3_xxxy_inst_n59), .B(prince_inst_sin_y[15]), .Z(
        prince_inst_sbox_inst3_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U20 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U19 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n58) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U18 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst3_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst3_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n66), .A2(prince_inst_sin_x[14]), 
        .ZN(prince_inst_sbox_inst3_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst3_xxxy_inst_U16 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sin_y[15]), .A3(prince_inst_sbox_inst3_xxxy_inst_n68), 
        .ZN(prince_inst_sbox_inst3_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst3_xxxy_inst_U15 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst3_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst3_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst3_xxxy_inst_U14 ( .A(prince_inst_sin_x[12]), 
        .B(prince_inst_sbox_inst3_xxxy_inst_n61), .S(
        prince_inst_sbox_inst3_xxxy_inst_n67), .Z(
        prince_inst_sbox_inst3_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst3_xxxy_inst_U13 ( .A(prince_inst_sin_y[15]), 
        .ZN(prince_inst_sbox_inst3_xxxy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U12 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n61), .A2(prince_inst_sin_x[12]), 
        .ZN(prince_inst_sbox_inst3_xxxy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U11 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst3_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst3_xxxy_inst_U10 ( .A(
        prince_inst_sbox_inst3_xxxy_inst_n60), .B(
        prince_inst_sbox_inst3_xxxy_inst_n53), .S(
        prince_inst_sbox_inst3_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst3_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U9 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sbox_inst3_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U8 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n61), .A2(prince_inst_sin_y[15]), 
        .ZN(prince_inst_sbox_inst3_xxxy_inst_n66) );
  INV_X1 prince_inst_sbox_inst3_xxxy_inst_U7 ( .A(
        prince_inst_sbox_inst3_xxxy_inst_n68), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst3_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst3_t1_sh[0]), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst3_xxxy_inst_U5 ( .A(prince_inst_sin_x[14]), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U4 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst3_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst3_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst3_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst3_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst3_xxxy_inst_U2 ( .A(prince_inst_sin_x[12]), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n62) );
  INV_X1 prince_inst_sbox_inst3_xxxy_inst_U1 ( .A(prince_inst_sin_x[13]), .ZN(
        prince_inst_sbox_inst3_xxxy_inst_n68) );
  XOR2_X1 prince_inst_sbox_inst3_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst3_t1_sh[1]), .B(
        prince_inst_sbox_inst3_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst3_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst3_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst3_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst3_xxyx_inst_n52), .B(
        prince_inst_sbox_inst3_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst3_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U23 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst3_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst3_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n48), .A2(prince_inst_sin_x[15]), 
        .A3(prince_inst_sin_x[12]), .ZN(prince_inst_sbox_inst3_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n45), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst3_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst3_xxyx_inst_U18 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n46), .A2(prince_inst_sin_x[15]), 
        .A3(prince_inst_sin_x[13]), .ZN(prince_inst_sbox_inst3_xxyx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst3_t2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst3_xxyx_inst_U16 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sin_x[12]), .A3(prince_inst_sbox_inst3_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst3_xxyx_inst_n44) );
  OR2_X1 prince_inst_sbox_inst3_xxyx_inst_U15 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sbox_inst3_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst3_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst3_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst3_xxyx_inst_n54), .B(
        prince_inst_sbox_inst3_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst3_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U12 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sin_y[14]), .ZN(prince_inst_sbox_inst3_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst3_xxyx_inst_U11 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sbox_inst3_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst3_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst3_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst3_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst3_xxyx_inst_U10 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst3_xxyx_inst_U9 ( .A1(prince_inst_sin_x[15]), 
        .A2(prince_inst_sbox_inst3_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst3_xxyx_inst_U8 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sbox_inst3_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst3_xxyx_inst_U7 ( .A(prince_inst_sin_y[14]), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst3_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst3_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst3_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n53), .A2(prince_inst_sin_x[13]), 
        .A3(prince_inst_sin_y[14]), .A4(prince_inst_sin_x[12]), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst3_xxyx_inst_U4 ( .A(prince_inst_sin_x[15]), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst3_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst3_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst3_xxyx_inst_n43), .A3(prince_inst_sin_x[15]), 
        .A4(prince_inst_sin_y[14]), .ZN(prince_inst_sbox_inst3_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst3_xxyx_inst_U2 ( .A(prince_inst_sin_x[12]), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst3_xxyx_inst_U1 ( .A(prince_inst_sin_x[13]), .ZN(
        prince_inst_sbox_inst3_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst3_xyxx_inst_n74), .B(
        prince_inst_sbox_inst3_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst3_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst3_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst3_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst3_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U26 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sbox_inst3_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U25 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst3_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst3_xyxx_inst_n72), .B(
        prince_inst_sbox_inst3_s0_sh[2]), .S(
        prince_inst_sbox_inst3_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst3_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst3_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n74), .A2(prince_inst_sin_x[15]), 
        .ZN(prince_inst_sbox_inst3_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst3_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U21 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst3_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst3_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst3_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst3_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst3_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst3_xyxx_inst_U15 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_x[12]), .ZN(prince_inst_sbox_inst3_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst3_xyxx_inst_U13 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U12 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_x[14]), .ZN(prince_inst_sbox_inst3_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst3_xyxx_inst_n58), .B(
        prince_inst_sbox_inst3_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst3_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst3_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst3_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst3_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst3_xyxx_inst_U9 ( .A(prince_inst_sin_x[15]), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst3_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n54), .A2(prince_inst_sin_x[12]), 
        .ZN(prince_inst_sbox_inst3_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst3_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst3_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst3_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst3_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst3_xyxx_inst_U5 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst3_xyxx_inst_U4 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst3_xyxx_inst_U3 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sbox_inst3_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst3_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst3_xyxx_inst_U2 ( .A(prince_inst_sin_y[13]), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst3_xyxx_inst_U1 ( .A(prince_inst_sin_x[14]), .ZN(
        prince_inst_sbox_inst3_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst3_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst3_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst3_xyyy_inst_n59), .B(
        prince_inst_sbox_inst3_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst3_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst3_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst3_xyyy_inst_U25 ( .A1(prince_inst_sin_y[14]), 
        .A2(prince_inst_sin_y[15]), .A3(prince_inst_sbox_inst3_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst3_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U24 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sbox_inst3_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U23 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sbox_inst3_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst3_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst3_xyyy_inst_U19 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sin_y[14]), .A3(prince_inst_sbox_inst3_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst3_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst3_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst3_xyyy_inst_n49), .B(
        prince_inst_sbox_inst3_xyyy_inst_n48), .S(
        prince_inst_sbox_inst3_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst3_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst3_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst3_xyyy_inst_U16 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sbox_inst3_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst3_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst3_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst3_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst3_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst3_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst3_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst3_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst3_xyyy_inst_U12 ( .A(prince_inst_sin_y[15]), 
        .ZN(prince_inst_sbox_inst3_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst3_xyyy_inst_U11 ( .A1(prince_inst_sin_y[15]), 
        .A2(prince_inst_sbox_inst3_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst3_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst3_t1_sh[3]), .B(
        prince_inst_sbox_inst3_xyyy_inst_n48), .S(
        prince_inst_sbox_inst3_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst3_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst3_xyyy_inst_U9 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sbox_inst3_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst3_xyyy_inst_U8 ( .A1(prince_inst_sin_x[12]), 
        .A2(prince_inst_sin_y[15]), .ZN(prince_inst_sbox_inst3_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst3_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst3_t1_sh[3]), .ZN(prince_inst_sbox_inst3_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst3_xyyy_inst_U6 ( .A1(prince_inst_sin_y[15]), 
        .A2(prince_inst_sbox_inst3_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst3_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst3_xyyy_inst_U4 ( .A(prince_inst_sin_y[13]), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst3_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst3_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst3_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst3_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst3_xyyy_inst_U2 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_x[12]), .ZN(prince_inst_sbox_inst3_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst3_xyyy_inst_U1 ( .A(prince_inst_sin_y[14]), .ZN(
        prince_inst_sbox_inst3_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst3_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U27 ( .A1(prince_inst_sin_y[12]), 
        .A2(prince_inst_sbox_inst3_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst3_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U24 ( .A1(prince_inst_sin_y[12]), 
        .A2(prince_inst_sbox_inst3_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst3_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U21 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst3_yxxx_inst_U19 ( .A(prince_inst_sin_x[15]), 
        .ZN(prince_inst_sbox_inst3_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst3_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst3_yxxx_inst_n52), .B(
        prince_inst_sbox_inst3_yxxx_inst_n51), .S(
        prince_inst_sbox_inst3_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst3_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n53), .A2(prince_inst_sin_x[15]), 
        .ZN(prince_inst_sbox_inst3_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst3_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n48), .A2(prince_inst_sin_y[12]), 
        .ZN(prince_inst_sbox_inst3_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n47), .A2(prince_inst_sin_x[15]), 
        .ZN(prince_inst_sbox_inst3_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U13 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sbox_inst3_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst3_yxxx_inst_n59), .B(
        prince_inst_sbox_inst3_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst3_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst3_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst3_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst3_yxxx_inst_U9 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sbox_inst3_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst3_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst3_yxxx_inst_U8 ( .A(prince_inst_sin_x[14]), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst3_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst3_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst3_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst3_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst3_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst3_yxxx_inst_U5 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst3_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst3_yxxx_inst_U4 ( .A(prince_inst_sin_y[12]), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst3_yxxx_inst_U3 ( .A(prince_inst_sin_x[13]), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst3_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst3_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst3_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst3_yxxx_inst_U1 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n67), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n66), .ZN(
        prince_inst_sbox_inst3_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst3_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n66), .A3(
        prince_inst_sbox_inst3_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst3_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst3_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n64), .A2(prince_inst_sin_x[13]), 
        .A3(prince_inst_sin_y[15]), .ZN(prince_inst_sbox_inst3_yxyy_inst_n66)
         );
  NAND3_X1 prince_inst_sbox_inst3_yxyy_inst_U24 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n63), .A2(prince_inst_sin_y[14]), 
        .A3(prince_inst_sin_y[15]), .ZN(prince_inst_sbox_inst3_yxyy_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst3_yxyy_inst_U23 ( .A(
        prince_inst_sbox_inst3_yxyy_inst_n62), .B(
        prince_inst_sbox_inst3_yxyy_inst_n61), .S(prince_inst_sin_y[12]), .Z(
        prince_inst_sbox_inst3_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst3_yxyy_inst_U22 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n64), .A2(prince_inst_sin_x[13]), 
        .ZN(prince_inst_sbox_inst3_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst3_yxyy_inst_U21 ( .A(prince_inst_sin_x[13]), 
        .B(prince_inst_sbox_inst3_yxyy_inst_n60), .S(
        prince_inst_sbox_inst3_yxyy_inst_n64), .Z(
        prince_inst_sbox_inst3_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U18 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst3_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst3_yxyy_inst_n62), .B(
        prince_inst_sbox_inst3_yxyy_inst_n54), .S(
        prince_inst_sbox_inst3_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst3_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst3_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst3_yxyy_inst_n53), .B(
        prince_inst_sbox_inst3_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst3_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst3_yxyy_inst_U15 ( .A(
        prince_inst_sbox_inst3_yxyy_inst_n67), .B(
        prince_inst_sbox_inst3_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst3_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U14 ( .A1(prince_inst_sin_y[15]), 
        .A2(prince_inst_sin_y[12]), .ZN(prince_inst_sbox_inst3_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst3_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst3_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst3_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst3_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst3_yxyy_inst_U12 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst3_yxyy_inst_U11 ( .A(
        prince_inst_sbox_inst3_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst3_yxyy_inst_U10 ( .A1(prince_inst_sin_x[13]), 
        .A2(prince_inst_sin_y[14]), .A3(prince_inst_sin_y[12]), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U9 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst3_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U8 ( .A1(prince_inst_sin_y[15]), 
        .A2(prince_inst_sbox_inst3_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst3_yxyy_inst_U7 ( .A1(prince_inst_sin_y[14]), 
        .A2(prince_inst_sin_x[13]), .ZN(prince_inst_sbox_inst3_yxyy_inst_n49)
         );
  OR3_X1 prince_inst_sbox_inst3_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst3_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst3_yxyy_inst_U5 ( .A(prince_inst_sin_y[12]), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst3_yxyy_inst_U4 ( .A(prince_inst_sin_x[13]), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst3_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst3_yxyy_inst_n64), .A2(
        prince_inst_sbox_inst3_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst3_yxyy_inst_U2 ( .A(prince_inst_sin_y[15]), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst3_yxyy_inst_U1 ( .A(prince_inst_sin_y[14]), .ZN(
        prince_inst_sbox_inst3_yxyy_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst3_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U29 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst3_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst3_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst3_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n75), .A2(prince_inst_sin_y[15]), 
        .A3(prince_inst_sbox_inst3_yyxy_inst_n70), .A4(prince_inst_sin_x[14]), 
        .ZN(prince_inst_sbox_inst3_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst3_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n69), .A3(prince_inst_sin_y[13]), 
        .A4(prince_inst_sbox_inst3_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst3_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst3_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst3_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst3_yyxy_inst_U23 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_x[14]), .A3(prince_inst_sin_y[12]), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst3_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n69), .A2(prince_inst_sin_y[13]), 
        .A3(prince_inst_sin_y[15]), .ZN(prince_inst_sbox_inst3_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst3_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n75), .A2(prince_inst_sin_x[14]), 
        .A3(prince_inst_sin_y[15]), .ZN(prince_inst_sbox_inst3_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst3_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst3_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst3_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n61), .A2(prince_inst_sin_x[14]), 
        .ZN(prince_inst_sbox_inst3_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst3_yyxy_inst_U18 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_y[15]), .A3(prince_inst_sbox_inst3_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst3_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst3_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst3_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst3_yyxy_inst_U16 ( .A1(prince_inst_sin_y[15]), 
        .A2(prince_inst_sbox_inst3_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst3_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst3_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst3_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n58), .A3(prince_inst_sin_y[12]), 
        .ZN(prince_inst_sbox_inst3_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst3_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst3_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst3_yyxy_inst_U13 ( .A1(prince_inst_sin_y[12]), 
        .A2(prince_inst_sbox_inst3_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst3_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst3_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst3_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst3_yyxy_inst_n54), .B(
        prince_inst_sbox_inst3_yyxy_inst_n55), .S(
        prince_inst_sbox_inst3_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst3_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst3_yyxy_inst_U9 ( .A(prince_inst_sin_x[14]), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n75), .A2(prince_inst_sin_y[15]), 
        .ZN(prince_inst_sbox_inst3_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst3_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst3_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst3_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U5 ( .A1(prince_inst_sin_x[14]), 
        .A2(prince_inst_sbox_inst3_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst3_yyxy_inst_U4 ( .A(prince_inst_sin_y[13]), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst3_yyxy_inst_U3 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sbox_inst3_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst3_yyxy_inst_U2 ( .A(prince_inst_sin_y[12]), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst3_yyxy_inst_U1 ( .A(prince_inst_sin_y[15]), .ZN(
        prince_inst_sbox_inst3_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst3_yyyx_inst_n58), .B(
        prince_inst_sbox_inst3_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst3_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst3_yyyx_inst_n56), .B(
        prince_inst_sbox_inst3_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst3_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst3_yyyx_inst_n54), .B(
        prince_inst_sbox_inst3_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst3_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst3_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst3_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst3_yyyx_inst_U21 ( .A1(prince_inst_sin_x[15]), 
        .A2(prince_inst_sbox_inst3_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst3_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst3_yyyx_inst_U20 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_y[14]), .A3(prince_inst_sbox_inst3_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst3_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst3_yyyx_inst_n50), .B(
        prince_inst_sbox_inst3_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst3_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst3_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n56), .A2(prince_inst_sin_y[14]), 
        .ZN(prince_inst_sbox_inst3_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst3_yyyx_inst_U17 ( .A1(prince_inst_sin_y[13]), 
        .A2(prince_inst_sin_y[12]), .A3(prince_inst_sin_y[14]), .ZN(
        prince_inst_sbox_inst3_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst3_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst3_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst3_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst3_yyyx_inst_U15 ( .A1(prince_inst_sin_x[15]), 
        .A2(prince_inst_sin_y[14]), .A3(prince_inst_sbox_inst3_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst3_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst3_yyyx_inst_U14 ( .A(prince_inst_sin_y[12]), 
        .ZN(prince_inst_sbox_inst3_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n58), .A2(prince_inst_sin_y[13]), 
        .ZN(prince_inst_sbox_inst3_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst3_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst3_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U11 ( .A1(prince_inst_sin_y[12]), 
        .A2(prince_inst_sbox_inst3_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst3_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst3_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst3_yyyx_inst_U9 ( .A1(prince_inst_sin_y[12]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst3_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst3_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst3_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst3_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n45), .A2(prince_inst_sin_y[12]), 
        .A3(prince_inst_sin_y[14]), .ZN(prince_inst_sbox_inst3_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst3_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst3_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst3_yyyx_inst_U4 ( .A1(prince_inst_sin_x[15]), 
        .A2(prince_inst_sin_y[14]), .ZN(prince_inst_sbox_inst3_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst3_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst3_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst3_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst3_yyyx_inst_U2 ( .A(prince_inst_sin_y[13]), .ZN(
        prince_inst_sbox_inst3_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst3_yyyx_inst_U1 ( .A1(prince_inst_sin_y[12]), 
        .A2(prince_inst_sin_x[15]), .ZN(prince_inst_sbox_inst3_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s00_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[0]), .B(prince_inst_sbox_inst3_s0_sh[0]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s01_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[1]), .B(prince_inst_sbox_inst3_s0_sh[1]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s02_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[2]), .B(prince_inst_sbox_inst3_s0_sh[2]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s03_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[3]), .B(prince_inst_sbox_inst3_s0_sh[3]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s04_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[4]), .B(prince_inst_sbox_inst3_s0_sh[4]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s05_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[5]), .B(prince_inst_sbox_inst3_s0_sh[5]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s06_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[6]), .B(prince_inst_sbox_inst3_s0_sh[6]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s07_U1 ( .A(
        prince_inst_sbox_inst3_t0_sh[7]), .B(prince_inst_sbox_inst3_s0_sh[7]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s10_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[0]), .B(prince_inst_sbox_inst3_s1_sh[0]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s11_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[1]), .B(prince_inst_sbox_inst3_s1_sh[1]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s12_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[2]), .B(prince_inst_sbox_inst3_s1_sh[2]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s13_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[3]), .B(prince_inst_sbox_inst3_s1_sh[3]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s14_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[4]), .B(prince_inst_sbox_inst3_s1_sh[4]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s15_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[5]), .B(prince_inst_sbox_inst3_s1_sh[5]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s16_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[6]), .B(prince_inst_sbox_inst3_s1_sh[6]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s17_U1 ( .A(
        prince_inst_sbox_inst3_t1_sh[7]), .B(prince_inst_sbox_inst3_s1_sh[7]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s20_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[0]), .B(prince_inst_sbox_inst3_s2_sh[0]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s21_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[1]), .B(prince_inst_sbox_inst3_s2_sh[1]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s22_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[2]), .B(prince_inst_sbox_inst3_s2_sh[2]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s23_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[3]), .B(prince_inst_sbox_inst3_s2_sh[3]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s24_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[4]), .B(prince_inst_sbox_inst3_s2_sh[4]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s25_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[5]), .B(prince_inst_sbox_inst3_s2_sh[5]), 
        .S(prince_inst_sbox_inst3_n8), .Z(prince_inst_sbox_inst3_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s26_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[6]), .B(prince_inst_sbox_inst3_s2_sh[6]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s27_U1 ( .A(
        prince_inst_sbox_inst3_t2_sh[7]), .B(prince_inst_sbox_inst3_s2_sh[7]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s30_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[0]), .B(prince_inst_sbox_inst3_s3_sh[0]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s31_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[1]), .B(prince_inst_sbox_inst3_s3_sh[1]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s32_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[2]), .B(prince_inst_sbox_inst3_s3_sh[2]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s33_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[3]), .B(prince_inst_sbox_inst3_s3_sh[3]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s34_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[4]), .B(prince_inst_sbox_inst3_s3_sh[4]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s35_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[5]), .B(prince_inst_sbox_inst3_s3_sh[5]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s36_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[6]), .B(prince_inst_sbox_inst3_s3_sh[6]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst3_mux_s37_U1 ( .A(
        prince_inst_sbox_inst3_t3_sh[7]), .B(prince_inst_sbox_inst3_s3_sh[7]), 
        .S(prince_inst_sbox_inst3_n9), .Z(prince_inst_sbox_inst3_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk0_U1 ( .A(r[48]), .B(
        prince_inst_sbox_inst3_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk1_U1 ( .A(r[49]), .B(
        prince_inst_sbox_inst3_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk2_U1 ( .A(r[50]), .B(
        prince_inst_sbox_inst3_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk3_U1 ( .A(r[51]), .B(
        prince_inst_sbox_inst3_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk4_U1 ( .A(r[48]), .B(
        prince_inst_sbox_inst3_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk5_U1 ( .A(r[49]), .B(
        prince_inst_sbox_inst3_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk6_U1 ( .A(r[50]), .B(
        prince_inst_sbox_inst3_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_msk7_U1 ( .A(r[51]), .B(
        prince_inst_sbox_inst3_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst3_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst3_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst3_c_inst0_ax_n5), .ZN(prince_inst_sout_x[12]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst3_c_inst0_y[1]), .B(
        prince_inst_sbox_inst3_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst3_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst3_c_inst0_y[2]), .B(
        prince_inst_sbox_inst3_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst3_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst3_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst3_c_inst0_ay_n5), .ZN(final_y[12]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst3_c_inst0_y[5]), .B(
        prince_inst_sbox_inst3_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst3_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst3_c_inst0_y[6]), .B(
        prince_inst_sbox_inst3_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst3_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk0_U1 ( .A(r[52]), .B(
        prince_inst_sbox_inst3_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk1_U1 ( .A(r[53]), .B(
        prince_inst_sbox_inst3_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk2_U1 ( .A(r[54]), .B(
        prince_inst_sbox_inst3_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk3_U1 ( .A(r[55]), .B(
        prince_inst_sbox_inst3_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk4_U1 ( .A(r[52]), .B(
        prince_inst_sbox_inst3_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk5_U1 ( .A(r[53]), .B(
        prince_inst_sbox_inst3_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk6_U1 ( .A(r[54]), .B(
        prince_inst_sbox_inst3_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_msk7_U1 ( .A(r[55]), .B(
        prince_inst_sbox_inst3_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst3_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst3_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst3_c_inst1_ax_n5), .ZN(prince_inst_sout_x[13]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst3_c_inst1_y[1]), .B(
        prince_inst_sbox_inst3_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst3_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst3_c_inst1_y[2]), .B(
        prince_inst_sbox_inst3_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst3_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst3_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst3_c_inst1_ay_n5), .ZN(final_y[13]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst3_c_inst1_y[5]), .B(
        prince_inst_sbox_inst3_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst3_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst3_c_inst1_y[6]), .B(
        prince_inst_sbox_inst3_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst3_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk0_U1 ( .A(r[56]), .B(
        prince_inst_sbox_inst3_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk1_U1 ( .A(r[57]), .B(
        prince_inst_sbox_inst3_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk2_U1 ( .A(r[58]), .B(
        prince_inst_sbox_inst3_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk3_U1 ( .A(r[59]), .B(
        prince_inst_sbox_inst3_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk4_U1 ( .A(r[56]), .B(
        prince_inst_sbox_inst3_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk5_U1 ( .A(r[57]), .B(
        prince_inst_sbox_inst3_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk6_U1 ( .A(r[58]), .B(
        prince_inst_sbox_inst3_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_msk7_U1 ( .A(r[59]), .B(
        prince_inst_sbox_inst3_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst3_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst3_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst3_c_inst2_ax_n5), .ZN(prince_inst_sout_x[14]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst3_c_inst2_y[1]), .B(
        prince_inst_sbox_inst3_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst3_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst3_c_inst2_y[2]), .B(
        prince_inst_sbox_inst3_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst3_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst3_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst3_c_inst2_ay_n5), .ZN(final_y[14]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst3_c_inst2_y[5]), .B(
        prince_inst_sbox_inst3_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst3_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst3_c_inst2_y[6]), .B(
        prince_inst_sbox_inst3_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst3_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk0_U1 ( .A(r[60]), .B(
        prince_inst_sbox_inst3_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk1_U1 ( .A(r[61]), .B(
        prince_inst_sbox_inst3_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk2_U1 ( .A(r[62]), .B(
        prince_inst_sbox_inst3_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk3_U1 ( .A(r[63]), .B(
        prince_inst_sbox_inst3_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk4_U1 ( .A(r[60]), .B(
        prince_inst_sbox_inst3_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk5_U1 ( .A(r[61]), .B(
        prince_inst_sbox_inst3_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk6_U1 ( .A(r[62]), .B(
        prince_inst_sbox_inst3_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_msk7_U1 ( .A(r[63]), .B(
        prince_inst_sbox_inst3_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst3_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst3_n6), .A3(
        prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst3_n11), .A2(prince_inst_sbox_inst3_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst3_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst3_n11), .ZN(
        prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst3_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst3_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst3_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst3_c_inst3_ax_n5), .ZN(prince_inst_sout_x[15]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst3_c_inst3_y[1]), .B(
        prince_inst_sbox_inst3_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst3_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst3_c_inst3_y[2]), .B(
        prince_inst_sbox_inst3_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst3_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst3_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst3_c_inst3_ay_n5), .ZN(final_y[15]) );
  XNOR2_X1 prince_inst_sbox_inst3_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst3_c_inst3_y[5]), .B(
        prince_inst_sbox_inst3_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst3_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst3_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst3_c_inst3_y[6]), .B(
        prince_inst_sbox_inst3_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst3_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst4_U7 ( .A(prince_inst_sbox_inst4_n12), .ZN(
        prince_inst_sbox_inst4_n11) );
  INV_X1 prince_inst_sbox_inst4_U6 ( .A(prince_inst_n28), .ZN(
        prince_inst_sbox_inst4_n10) );
  INV_X1 prince_inst_sbox_inst4_U5 ( .A(prince_inst_sbox_inst4_n10), .ZN(
        prince_inst_sbox_inst4_n8) );
  INV_X1 prince_inst_sbox_inst4_U4 ( .A(prince_inst_sbox_inst4_n10), .ZN(
        prince_inst_sbox_inst4_n9) );
  INV_X1 prince_inst_sbox_inst4_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst4_n12) );
  INV_X1 prince_inst_sbox_inst4_U2 ( .A(rst), .ZN(prince_inst_sbox_inst4_n7)
         );
  INV_X2 prince_inst_sbox_inst4_U1 ( .A(prince_inst_sbox_inst4_n7), .ZN(
        prince_inst_sbox_inst4_n6) );
  NAND3_X1 prince_inst_sbox_inst4_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n68), .A3(prince_inst_sin_x[16]), 
        .ZN(prince_inst_sbox_inst4_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U25 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sbox_inst4_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst4_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst4_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst4_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst4_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n67), .A2(prince_inst_sin_x[18]), 
        .A3(prince_inst_sin_x[16]), .A4(prince_inst_sin_y[19]), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst4_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n61), .A2(prince_inst_sin_x[17]), 
        .A3(prince_inst_sin_x[18]), .ZN(prince_inst_sbox_inst4_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst4_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n66), .A3(prince_inst_sin_x[17]), 
        .A4(prince_inst_sin_x[16]), .ZN(prince_inst_sbox_inst4_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst4_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst4_xxxy_inst_n59), .B(prince_inst_sin_y[19]), .Z(
        prince_inst_sbox_inst4_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U18 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sin_x[17]), .ZN(prince_inst_sbox_inst4_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst4_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst4_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n65), .A2(prince_inst_sin_x[18]), 
        .ZN(prince_inst_sbox_inst4_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst4_xxxy_inst_U15 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sin_y[19]), .A3(prince_inst_sbox_inst4_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst4_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst4_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst4_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst4_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst4_xxxy_inst_U13 ( .A(prince_inst_sin_x[16]), 
        .B(prince_inst_sin_x[17]), .S(prince_inst_sbox_inst4_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst4_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst4_xxxy_inst_U12 ( .A(prince_inst_sin_y[19]), 
        .ZN(prince_inst_sbox_inst4_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U11 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sin_x[16]), .ZN(prince_inst_sbox_inst4_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst4_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst4_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst4_xxxy_inst_n60), .B(
        prince_inst_sbox_inst4_xxxy_inst_n53), .S(
        prince_inst_sbox_inst4_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst4_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U8 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sbox_inst4_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U7 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sin_y[19]), .ZN(prince_inst_sbox_inst4_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst4_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst4_t1_sh[0]), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst4_xxxy_inst_U5 ( .A(prince_inst_sin_x[18]), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U4 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sbox_inst4_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst4_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst4_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst4_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst4_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst4_xxxy_inst_U2 ( .A(prince_inst_sin_x[16]), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst4_xxxy_inst_U1 ( .A(prince_inst_sin_x[17]), .ZN(
        prince_inst_sbox_inst4_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst4_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst4_t1_sh[1]), .B(
        prince_inst_sbox_inst4_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst4_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst4_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst4_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst4_xxyx_inst_n52), .B(
        prince_inst_sbox_inst4_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst4_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U23 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst4_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst4_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n48), .A2(prince_inst_sin_x[19]), 
        .A3(prince_inst_sin_x[16]), .ZN(prince_inst_sbox_inst4_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst4_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst4_xxyx_inst_U18 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sbox_inst4_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst4_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst4_xxyx_inst_U16 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sin_x[16]), .A3(prince_inst_sbox_inst4_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst4_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst4_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n46), .A2(prince_inst_sin_x[19]), 
        .A3(prince_inst_sin_x[17]), .ZN(prince_inst_sbox_inst4_xxyx_inst_n44)
         );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst4_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst4_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst4_xxyx_inst_n54), .B(
        prince_inst_sbox_inst4_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst4_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U12 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sin_y[18]), .ZN(prince_inst_sbox_inst4_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst4_xxyx_inst_U11 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sbox_inst4_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst4_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst4_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst4_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst4_xxyx_inst_U10 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst4_xxyx_inst_U9 ( .A1(prince_inst_sin_x[19]), 
        .A2(prince_inst_sbox_inst4_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst4_xxyx_inst_U8 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sbox_inst4_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst4_xxyx_inst_U7 ( .A(prince_inst_sin_y[18]), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst4_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst4_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst4_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n53), .A2(prince_inst_sin_x[17]), 
        .A3(prince_inst_sin_y[18]), .A4(prince_inst_sin_x[16]), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst4_xxyx_inst_U4 ( .A(prince_inst_sin_x[19]), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst4_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst4_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst4_xxyx_inst_n43), .A3(prince_inst_sin_x[19]), 
        .A4(prince_inst_sin_y[18]), .ZN(prince_inst_sbox_inst4_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst4_xxyx_inst_U2 ( .A(prince_inst_sin_x[16]), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst4_xxyx_inst_U1 ( .A(prince_inst_sin_x[17]), .ZN(
        prince_inst_sbox_inst4_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst4_xyxx_inst_n74), .B(
        prince_inst_sbox_inst4_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst4_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst4_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst4_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst4_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U26 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sbox_inst4_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U25 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst4_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst4_xyxx_inst_n72), .B(
        prince_inst_sbox_inst4_s0_sh[2]), .S(
        prince_inst_sbox_inst4_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst4_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst4_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n74), .A2(prince_inst_sin_x[19]), 
        .ZN(prince_inst_sbox_inst4_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst4_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U21 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sbox_inst4_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst4_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst4_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst4_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst4_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst4_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst4_xyxx_inst_U15 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_x[16]), .ZN(prince_inst_sbox_inst4_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst4_xyxx_inst_U13 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U12 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_x[18]), .ZN(prince_inst_sbox_inst4_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst4_xyxx_inst_n58), .B(
        prince_inst_sbox_inst4_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst4_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst4_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst4_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst4_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst4_xyxx_inst_U9 ( .A(prince_inst_sin_x[19]), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst4_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n54), .A2(prince_inst_sin_x[16]), 
        .ZN(prince_inst_sbox_inst4_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst4_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst4_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst4_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst4_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst4_xyxx_inst_U5 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sbox_inst4_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst4_xyxx_inst_U4 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst4_xyxx_inst_U3 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sbox_inst4_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst4_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst4_xyxx_inst_U2 ( .A(prince_inst_sin_y[17]), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst4_xyxx_inst_U1 ( .A(prince_inst_sin_x[18]), .ZN(
        prince_inst_sbox_inst4_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst4_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst4_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst4_xyyy_inst_n59), .B(
        prince_inst_sbox_inst4_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst4_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst4_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst4_xyyy_inst_U25 ( .A1(prince_inst_sin_y[18]), 
        .A2(prince_inst_sin_y[19]), .A3(prince_inst_sbox_inst4_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst4_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U24 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sbox_inst4_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U23 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sbox_inst4_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst4_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst4_xyyy_inst_U19 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sin_y[18]), .A3(prince_inst_sbox_inst4_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst4_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst4_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst4_xyyy_inst_n49), .B(
        prince_inst_sbox_inst4_xyyy_inst_n48), .S(
        prince_inst_sbox_inst4_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst4_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst4_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst4_xyyy_inst_U16 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sbox_inst4_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst4_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst4_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst4_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst4_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst4_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst4_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst4_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst4_xyyy_inst_U12 ( .A(prince_inst_sin_y[19]), 
        .ZN(prince_inst_sbox_inst4_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst4_xyyy_inst_U11 ( .A1(prince_inst_sin_y[19]), 
        .A2(prince_inst_sbox_inst4_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst4_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst4_t1_sh[3]), .B(
        prince_inst_sbox_inst4_xyyy_inst_n48), .S(
        prince_inst_sbox_inst4_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst4_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst4_xyyy_inst_U9 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sbox_inst4_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst4_xyyy_inst_U8 ( .A1(prince_inst_sin_x[16]), 
        .A2(prince_inst_sin_y[19]), .ZN(prince_inst_sbox_inst4_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst4_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst4_t1_sh[3]), .ZN(prince_inst_sbox_inst4_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst4_xyyy_inst_U6 ( .A1(prince_inst_sin_y[19]), 
        .A2(prince_inst_sbox_inst4_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst4_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst4_xyyy_inst_U4 ( .A(prince_inst_sin_y[17]), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst4_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst4_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst4_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst4_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst4_xyyy_inst_U2 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_x[16]), .ZN(prince_inst_sbox_inst4_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst4_xyyy_inst_U1 ( .A(prince_inst_sin_y[18]), .ZN(
        prince_inst_sbox_inst4_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst4_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U27 ( .A1(prince_inst_sin_y[16]), 
        .A2(prince_inst_sbox_inst4_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst4_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U24 ( .A1(prince_inst_sin_y[16]), 
        .A2(prince_inst_sbox_inst4_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst4_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U21 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst4_yxxx_inst_U19 ( .A(prince_inst_sin_x[19]), 
        .ZN(prince_inst_sbox_inst4_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst4_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst4_yxxx_inst_n52), .B(
        prince_inst_sbox_inst4_yxxx_inst_n51), .S(
        prince_inst_sbox_inst4_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst4_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n53), .A2(prince_inst_sin_x[19]), 
        .ZN(prince_inst_sbox_inst4_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst4_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n48), .A2(prince_inst_sin_y[16]), 
        .ZN(prince_inst_sbox_inst4_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n47), .A2(prince_inst_sin_x[19]), 
        .ZN(prince_inst_sbox_inst4_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U13 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sbox_inst4_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst4_yxxx_inst_n59), .B(
        prince_inst_sbox_inst4_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst4_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst4_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst4_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst4_yxxx_inst_U9 ( .A1(prince_inst_sin_x[17]), 
        .A2(prince_inst_sbox_inst4_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst4_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst4_yxxx_inst_U8 ( .A(prince_inst_sin_x[18]), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst4_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst4_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst4_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst4_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst4_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst4_yxxx_inst_U5 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sbox_inst4_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst4_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst4_yxxx_inst_U4 ( .A(prince_inst_sin_y[16]), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst4_yxxx_inst_U3 ( .A(prince_inst_sin_x[17]), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst4_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst4_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst4_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst4_yxxx_inst_U1 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst4_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst4_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst4_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst4_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst4_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n64), .A3(prince_inst_sin_y[19]), 
        .ZN(prince_inst_sbox_inst4_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst4_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n63), .A2(prince_inst_sin_y[18]), 
        .A3(prince_inst_sin_y[19]), .ZN(prince_inst_sbox_inst4_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst4_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst4_yxyy_inst_n62), .B(
        prince_inst_sbox_inst4_yxyy_inst_n61), .S(prince_inst_sin_y[16]), .Z(
        prince_inst_sbox_inst4_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst4_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst4_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst4_yxyy_inst_n64), .B(
        prince_inst_sbox_inst4_yxyy_inst_n60), .S(
        prince_inst_sbox_inst4_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst4_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst4_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst4_yxyy_inst_n62), .B(
        prince_inst_sbox_inst4_yxyy_inst_n54), .S(
        prince_inst_sbox_inst4_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst4_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst4_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst4_yxyy_inst_n53), .B(
        prince_inst_sbox_inst4_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst4_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst4_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst4_yxyy_inst_n68), .B(
        prince_inst_sbox_inst4_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst4_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U15 ( .A1(prince_inst_sin_y[19]), 
        .A2(prince_inst_sin_y[16]), .ZN(prince_inst_sbox_inst4_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst4_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst4_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst4_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst4_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst4_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst4_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst4_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst4_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n64), .A2(prince_inst_sin_y[18]), 
        .A3(prince_inst_sin_y[16]), .ZN(prince_inst_sbox_inst4_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst4_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U9 ( .A1(prince_inst_sin_y[19]), 
        .A2(prince_inst_sbox_inst4_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst4_yxyy_inst_U8 ( .A1(prince_inst_sin_y[18]), 
        .A2(prince_inst_sbox_inst4_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst4_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst4_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst4_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst4_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst4_yxyy_inst_U5 ( .A(prince_inst_sin_y[16]), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst4_yxyy_inst_U4 ( .A(prince_inst_sin_x[17]), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst4_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst4_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst4_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst4_yxyy_inst_U2 ( .A(prince_inst_sin_y[19]), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst4_yxyy_inst_U1 ( .A(prince_inst_sin_y[18]), .ZN(
        prince_inst_sbox_inst4_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst4_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U29 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sbox_inst4_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst4_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst4_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst4_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n75), .A2(prince_inst_sin_y[19]), 
        .A3(prince_inst_sbox_inst4_yyxy_inst_n70), .A4(prince_inst_sin_x[18]), 
        .ZN(prince_inst_sbox_inst4_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst4_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n69), .A3(prince_inst_sin_y[17]), 
        .A4(prince_inst_sbox_inst4_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst4_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst4_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst4_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst4_yyxy_inst_U23 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_x[18]), .A3(prince_inst_sin_y[16]), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst4_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n69), .A2(prince_inst_sin_y[17]), 
        .A3(prince_inst_sin_y[19]), .ZN(prince_inst_sbox_inst4_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst4_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n75), .A2(prince_inst_sin_x[18]), 
        .A3(prince_inst_sin_y[19]), .ZN(prince_inst_sbox_inst4_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst4_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst4_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst4_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n61), .A2(prince_inst_sin_x[18]), 
        .ZN(prince_inst_sbox_inst4_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst4_yyxy_inst_U18 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_y[19]), .A3(prince_inst_sbox_inst4_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst4_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst4_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst4_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst4_yyxy_inst_U16 ( .A1(prince_inst_sin_y[19]), 
        .A2(prince_inst_sbox_inst4_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst4_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst4_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst4_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n58), .A3(prince_inst_sin_y[16]), 
        .ZN(prince_inst_sbox_inst4_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst4_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst4_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst4_yyxy_inst_U13 ( .A1(prince_inst_sin_y[16]), 
        .A2(prince_inst_sbox_inst4_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst4_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst4_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst4_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst4_yyxy_inst_n54), .B(
        prince_inst_sbox_inst4_yyxy_inst_n55), .S(
        prince_inst_sbox_inst4_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst4_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst4_yyxy_inst_U9 ( .A(prince_inst_sin_x[18]), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n75), .A2(prince_inst_sin_y[19]), 
        .ZN(prince_inst_sbox_inst4_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst4_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst4_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst4_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U5 ( .A1(prince_inst_sin_x[18]), 
        .A2(prince_inst_sbox_inst4_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst4_yyxy_inst_U4 ( .A(prince_inst_sin_y[17]), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst4_yyxy_inst_U3 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sbox_inst4_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst4_yyxy_inst_U2 ( .A(prince_inst_sin_y[16]), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst4_yyxy_inst_U1 ( .A(prince_inst_sin_y[19]), .ZN(
        prince_inst_sbox_inst4_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst4_yyyx_inst_n58), .B(
        prince_inst_sbox_inst4_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst4_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst4_yyyx_inst_n56), .B(
        prince_inst_sbox_inst4_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst4_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst4_yyyx_inst_n54), .B(
        prince_inst_sbox_inst4_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst4_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst4_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst4_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst4_yyyx_inst_U21 ( .A1(prince_inst_sin_x[19]), 
        .A2(prince_inst_sbox_inst4_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst4_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst4_yyyx_inst_U20 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_y[18]), .A3(prince_inst_sbox_inst4_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst4_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst4_yyyx_inst_n50), .B(
        prince_inst_sbox_inst4_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst4_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst4_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n56), .A2(prince_inst_sin_y[18]), 
        .ZN(prince_inst_sbox_inst4_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst4_yyyx_inst_U17 ( .A1(prince_inst_sin_y[17]), 
        .A2(prince_inst_sin_y[16]), .A3(prince_inst_sin_y[18]), .ZN(
        prince_inst_sbox_inst4_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst4_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst4_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst4_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst4_yyyx_inst_U15 ( .A1(prince_inst_sin_x[19]), 
        .A2(prince_inst_sin_y[18]), .A3(prince_inst_sbox_inst4_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst4_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst4_yyyx_inst_U14 ( .A(prince_inst_sin_y[16]), 
        .ZN(prince_inst_sbox_inst4_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n58), .A2(prince_inst_sin_y[17]), 
        .ZN(prince_inst_sbox_inst4_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst4_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst4_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U11 ( .A1(prince_inst_sin_y[16]), 
        .A2(prince_inst_sbox_inst4_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst4_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst4_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst4_yyyx_inst_U9 ( .A1(prince_inst_sin_y[16]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst4_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst4_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst4_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst4_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n45), .A2(prince_inst_sin_y[16]), 
        .A3(prince_inst_sin_y[18]), .ZN(prince_inst_sbox_inst4_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst4_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst4_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst4_yyyx_inst_U4 ( .A1(prince_inst_sin_x[19]), 
        .A2(prince_inst_sin_y[18]), .ZN(prince_inst_sbox_inst4_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst4_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst4_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst4_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst4_yyyx_inst_U2 ( .A(prince_inst_sin_y[17]), .ZN(
        prince_inst_sbox_inst4_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst4_yyyx_inst_U1 ( .A1(prince_inst_sin_y[16]), 
        .A2(prince_inst_sin_x[19]), .ZN(prince_inst_sbox_inst4_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s00_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[0]), .B(prince_inst_sbox_inst4_s0_sh[0]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s01_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[1]), .B(prince_inst_sbox_inst4_s0_sh[1]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s02_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[2]), .B(prince_inst_sbox_inst4_s0_sh[2]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s03_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[3]), .B(prince_inst_sbox_inst4_s0_sh[3]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s04_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[4]), .B(prince_inst_sbox_inst4_s0_sh[4]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s05_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[5]), .B(prince_inst_sbox_inst4_s0_sh[5]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s06_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[6]), .B(prince_inst_sbox_inst4_s0_sh[6]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s07_U1 ( .A(
        prince_inst_sbox_inst4_t0_sh[7]), .B(prince_inst_sbox_inst4_s0_sh[7]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s10_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[0]), .B(prince_inst_sbox_inst4_s1_sh[0]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s11_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[1]), .B(prince_inst_sbox_inst4_s1_sh[1]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s12_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[2]), .B(prince_inst_sbox_inst4_s1_sh[2]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s13_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[3]), .B(prince_inst_sbox_inst4_s1_sh[3]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s14_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[4]), .B(prince_inst_sbox_inst4_s1_sh[4]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s15_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[5]), .B(prince_inst_sbox_inst4_s1_sh[5]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s16_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[6]), .B(prince_inst_sbox_inst4_s1_sh[6]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s17_U1 ( .A(
        prince_inst_sbox_inst4_t1_sh[7]), .B(prince_inst_sbox_inst4_s1_sh[7]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s20_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[0]), .B(prince_inst_sbox_inst4_s2_sh[0]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s21_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[1]), .B(prince_inst_sbox_inst4_s2_sh[1]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s22_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[2]), .B(prince_inst_sbox_inst4_s2_sh[2]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s23_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[3]), .B(prince_inst_sbox_inst4_s2_sh[3]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s24_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[4]), .B(prince_inst_sbox_inst4_s2_sh[4]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s25_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[5]), .B(prince_inst_sbox_inst4_s2_sh[5]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s26_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[6]), .B(prince_inst_sbox_inst4_s2_sh[6]), 
        .S(prince_inst_sbox_inst4_n8), .Z(prince_inst_sbox_inst4_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s27_U1 ( .A(
        prince_inst_sbox_inst4_t2_sh[7]), .B(prince_inst_sbox_inst4_s2_sh[7]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s30_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[0]), .B(prince_inst_sbox_inst4_s3_sh[0]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s31_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[1]), .B(prince_inst_sbox_inst4_s3_sh[1]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s32_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[2]), .B(prince_inst_sbox_inst4_s3_sh[2]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s33_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[3]), .B(prince_inst_sbox_inst4_s3_sh[3]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s34_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[4]), .B(prince_inst_sbox_inst4_s3_sh[4]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s35_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[5]), .B(prince_inst_sbox_inst4_s3_sh[5]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s36_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[6]), .B(prince_inst_sbox_inst4_s3_sh[6]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst4_mux_s37_U1 ( .A(
        prince_inst_sbox_inst4_t3_sh[7]), .B(prince_inst_sbox_inst4_s3_sh[7]), 
        .S(prince_inst_sbox_inst4_n9), .Z(prince_inst_sbox_inst4_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk0_U1 ( .A(r[0]), .B(
        prince_inst_sbox_inst4_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk1_U1 ( .A(r[1]), .B(
        prince_inst_sbox_inst4_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk2_U1 ( .A(r[2]), .B(
        prince_inst_sbox_inst4_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk3_U1 ( .A(r[3]), .B(
        prince_inst_sbox_inst4_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk4_U1 ( .A(r[0]), .B(
        prince_inst_sbox_inst4_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk5_U1 ( .A(r[1]), .B(
        prince_inst_sbox_inst4_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk6_U1 ( .A(r[2]), .B(
        prince_inst_sbox_inst4_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_msk7_U1 ( .A(r[3]), .B(
        prince_inst_sbox_inst4_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst4_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst4_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst4_c_inst0_ax_n5), .ZN(prince_inst_sout_x[16]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst4_c_inst0_y[1]), .B(
        prince_inst_sbox_inst4_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst4_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst4_c_inst0_y[2]), .B(
        prince_inst_sbox_inst4_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst4_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst4_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst4_c_inst0_ay_n5), .ZN(final_y[0]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst4_c_inst0_y[5]), .B(
        prince_inst_sbox_inst4_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst4_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst4_c_inst0_y[6]), .B(
        prince_inst_sbox_inst4_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst4_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk0_U1 ( .A(r[4]), .B(
        prince_inst_sbox_inst4_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk1_U1 ( .A(r[5]), .B(
        prince_inst_sbox_inst4_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk2_U1 ( .A(r[6]), .B(
        prince_inst_sbox_inst4_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk3_U1 ( .A(r[7]), .B(
        prince_inst_sbox_inst4_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk4_U1 ( .A(r[4]), .B(
        prince_inst_sbox_inst4_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk5_U1 ( .A(r[5]), .B(
        prince_inst_sbox_inst4_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk6_U1 ( .A(r[6]), .B(
        prince_inst_sbox_inst4_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_msk7_U1 ( .A(r[7]), .B(
        prince_inst_sbox_inst4_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst4_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst4_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst4_c_inst1_ax_n5), .ZN(prince_inst_sout_x[17]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst4_c_inst1_y[1]), .B(
        prince_inst_sbox_inst4_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst4_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst4_c_inst1_y[2]), .B(
        prince_inst_sbox_inst4_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst4_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst4_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst4_c_inst1_ay_n5), .ZN(final_y[1]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst4_c_inst1_y[5]), .B(
        prince_inst_sbox_inst4_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst4_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst4_c_inst1_y[6]), .B(
        prince_inst_sbox_inst4_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst4_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk0_U1 ( .A(r[8]), .B(
        prince_inst_sbox_inst4_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk1_U1 ( .A(r[9]), .B(
        prince_inst_sbox_inst4_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk2_U1 ( .A(r[10]), .B(
        prince_inst_sbox_inst4_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk3_U1 ( .A(r[11]), .B(
        prince_inst_sbox_inst4_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk4_U1 ( .A(r[8]), .B(
        prince_inst_sbox_inst4_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk5_U1 ( .A(r[9]), .B(
        prince_inst_sbox_inst4_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk6_U1 ( .A(r[10]), .B(
        prince_inst_sbox_inst4_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_msk7_U1 ( .A(r[11]), .B(
        prince_inst_sbox_inst4_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst4_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst4_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst4_c_inst2_ax_n5), .ZN(prince_inst_sout_x[18]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst4_c_inst2_y[1]), .B(
        prince_inst_sbox_inst4_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst4_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst4_c_inst2_y[2]), .B(
        prince_inst_sbox_inst4_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst4_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst4_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst4_c_inst2_ay_n5), .ZN(final_y[2]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst4_c_inst2_y[5]), .B(
        prince_inst_sbox_inst4_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst4_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst4_c_inst2_y[6]), .B(
        prince_inst_sbox_inst4_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst4_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk0_U1 ( .A(r[12]), .B(
        prince_inst_sbox_inst4_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk1_U1 ( .A(r[13]), .B(
        prince_inst_sbox_inst4_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk2_U1 ( .A(r[14]), .B(
        prince_inst_sbox_inst4_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk3_U1 ( .A(r[15]), .B(
        prince_inst_sbox_inst4_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk4_U1 ( .A(r[12]), .B(
        prince_inst_sbox_inst4_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk5_U1 ( .A(r[13]), .B(
        prince_inst_sbox_inst4_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk6_U1 ( .A(r[14]), .B(
        prince_inst_sbox_inst4_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_msk7_U1 ( .A(r[15]), .B(
        prince_inst_sbox_inst4_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst4_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst4_n6), .A3(
        prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst4_n11), .A2(prince_inst_sbox_inst4_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst4_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst4_n11), .ZN(
        prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst4_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst4_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst4_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst4_c_inst3_ax_n5), .ZN(prince_inst_sout_x[19]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst4_c_inst3_y[1]), .B(
        prince_inst_sbox_inst4_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst4_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst4_c_inst3_y[2]), .B(
        prince_inst_sbox_inst4_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst4_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst4_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst4_c_inst3_ay_n5), .ZN(final_y[3]) );
  XNOR2_X1 prince_inst_sbox_inst4_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst4_c_inst3_y[5]), .B(
        prince_inst_sbox_inst4_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst4_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst4_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst4_c_inst3_y[6]), .B(
        prince_inst_sbox_inst4_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst4_c_inst3_ay_n6) );
  INV_X1 prince_inst_sbox_inst5_U7 ( .A(inv_sig), .ZN(
        prince_inst_sbox_inst5_n10) );
  INV_X4 prince_inst_sbox_inst5_U6 ( .A(prince_inst_sbox_inst5_n12), .ZN(
        prince_inst_sbox_inst5_n11) );
  INV_X1 prince_inst_sbox_inst5_U5 ( .A(prince_inst_sbox_inst5_n10), .ZN(
        prince_inst_sbox_inst5_n8) );
  INV_X1 prince_inst_sbox_inst5_U4 ( .A(prince_inst_sbox_inst5_n10), .ZN(
        prince_inst_sbox_inst5_n9) );
  INV_X1 prince_inst_sbox_inst5_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst5_n12) );
  INV_X1 prince_inst_sbox_inst5_U2 ( .A(rst), .ZN(prince_inst_sbox_inst5_n7)
         );
  INV_X2 prince_inst_sbox_inst5_U1 ( .A(prince_inst_sbox_inst5_n7), .ZN(
        prince_inst_sbox_inst5_n6) );
  NAND3_X1 prince_inst_sbox_inst5_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n68), .A3(prince_inst_sin_x[20]), 
        .ZN(prince_inst_sbox_inst5_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U25 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sbox_inst5_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst5_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst5_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst5_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst5_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n67), .A2(prince_inst_sin_x[22]), 
        .A3(prince_inst_sin_x[20]), .A4(prince_inst_sin_y[23]), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst5_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n61), .A2(prince_inst_sin_x[21]), 
        .A3(prince_inst_sin_x[22]), .ZN(prince_inst_sbox_inst5_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst5_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n66), .A3(prince_inst_sin_x[21]), 
        .A4(prince_inst_sin_x[20]), .ZN(prince_inst_sbox_inst5_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst5_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst5_xxxy_inst_n59), .B(prince_inst_sin_y[23]), .Z(
        prince_inst_sbox_inst5_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U18 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sin_x[21]), .ZN(prince_inst_sbox_inst5_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst5_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst5_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n65), .A2(prince_inst_sin_x[22]), 
        .ZN(prince_inst_sbox_inst5_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst5_xxxy_inst_U15 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sin_y[23]), .A3(prince_inst_sbox_inst5_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst5_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst5_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst5_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst5_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst5_xxxy_inst_U13 ( .A(prince_inst_sin_x[20]), 
        .B(prince_inst_sin_x[21]), .S(prince_inst_sbox_inst5_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst5_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst5_xxxy_inst_U12 ( .A(prince_inst_sin_y[23]), 
        .ZN(prince_inst_sbox_inst5_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U11 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sin_x[20]), .ZN(prince_inst_sbox_inst5_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst5_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst5_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst5_xxxy_inst_n60), .B(
        prince_inst_sbox_inst5_xxxy_inst_n53), .S(
        prince_inst_sbox_inst5_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst5_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U8 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sbox_inst5_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U7 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sin_y[23]), .ZN(prince_inst_sbox_inst5_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst5_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst5_t1_sh[0]), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst5_xxxy_inst_U5 ( .A(prince_inst_sin_x[22]), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U4 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sbox_inst5_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst5_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst5_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst5_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst5_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst5_xxxy_inst_U2 ( .A(prince_inst_sin_x[20]), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst5_xxxy_inst_U1 ( .A(prince_inst_sin_x[21]), .ZN(
        prince_inst_sbox_inst5_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst5_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst5_t1_sh[1]), .B(
        prince_inst_sbox_inst5_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst5_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst5_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst5_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst5_xxyx_inst_n52), .B(
        prince_inst_sbox_inst5_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst5_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U23 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst5_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst5_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n48), .A2(prince_inst_sin_x[23]), 
        .A3(prince_inst_sin_x[20]), .ZN(prince_inst_sbox_inst5_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n45), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst5_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst5_xxyx_inst_U18 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n46), .A2(prince_inst_sin_x[23]), 
        .A3(prince_inst_sin_x[21]), .ZN(prince_inst_sbox_inst5_xxyx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst5_t2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst5_xxyx_inst_U16 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sin_x[20]), .A3(prince_inst_sbox_inst5_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst5_xxyx_inst_n44) );
  OR2_X1 prince_inst_sbox_inst5_xxyx_inst_U15 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sbox_inst5_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst5_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst5_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst5_xxyx_inst_n54), .B(
        prince_inst_sbox_inst5_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst5_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U12 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sin_y[22]), .ZN(prince_inst_sbox_inst5_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst5_xxyx_inst_U11 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sbox_inst5_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst5_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst5_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst5_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst5_xxyx_inst_U10 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst5_xxyx_inst_U9 ( .A1(prince_inst_sin_x[23]), 
        .A2(prince_inst_sbox_inst5_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst5_xxyx_inst_U8 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sbox_inst5_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst5_xxyx_inst_U7 ( .A(prince_inst_sin_y[22]), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst5_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst5_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst5_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n53), .A2(prince_inst_sin_x[21]), 
        .A3(prince_inst_sin_y[22]), .A4(prince_inst_sin_x[20]), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst5_xxyx_inst_U4 ( .A(prince_inst_sin_x[23]), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst5_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst5_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst5_xxyx_inst_n43), .A3(prince_inst_sin_x[23]), 
        .A4(prince_inst_sin_y[22]), .ZN(prince_inst_sbox_inst5_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst5_xxyx_inst_U2 ( .A(prince_inst_sin_x[20]), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst5_xxyx_inst_U1 ( .A(prince_inst_sin_x[21]), .ZN(
        prince_inst_sbox_inst5_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst5_xyxx_inst_n74), .B(
        prince_inst_sbox_inst5_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst5_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst5_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst5_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst5_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U26 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sbox_inst5_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U25 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst5_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst5_xyxx_inst_n72), .B(
        prince_inst_sbox_inst5_s0_sh[2]), .S(
        prince_inst_sbox_inst5_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst5_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst5_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n74), .A2(prince_inst_sin_x[23]), 
        .ZN(prince_inst_sbox_inst5_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst5_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U21 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sbox_inst5_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst5_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst5_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst5_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst5_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst5_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst5_xyxx_inst_U15 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_x[20]), .ZN(prince_inst_sbox_inst5_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst5_xyxx_inst_U13 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U12 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_x[22]), .ZN(prince_inst_sbox_inst5_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst5_xyxx_inst_n58), .B(
        prince_inst_sbox_inst5_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst5_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst5_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst5_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst5_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst5_xyxx_inst_U9 ( .A(prince_inst_sin_x[23]), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst5_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n54), .A2(prince_inst_sin_x[20]), 
        .ZN(prince_inst_sbox_inst5_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst5_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst5_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst5_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst5_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst5_xyxx_inst_U5 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sbox_inst5_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst5_xyxx_inst_U4 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst5_xyxx_inst_U3 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sbox_inst5_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst5_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst5_xyxx_inst_U2 ( .A(prince_inst_sin_y[21]), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst5_xyxx_inst_U1 ( .A(prince_inst_sin_x[22]), .ZN(
        prince_inst_sbox_inst5_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst5_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst5_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst5_xyyy_inst_n59), .B(
        prince_inst_sbox_inst5_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst5_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst5_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst5_xyyy_inst_U25 ( .A1(prince_inst_sin_y[22]), 
        .A2(prince_inst_sin_y[23]), .A3(prince_inst_sbox_inst5_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst5_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U24 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sbox_inst5_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U23 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sbox_inst5_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst5_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst5_xyyy_inst_U19 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sin_y[22]), .A3(prince_inst_sbox_inst5_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst5_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst5_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst5_xyyy_inst_n49), .B(
        prince_inst_sbox_inst5_xyyy_inst_n48), .S(
        prince_inst_sbox_inst5_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst5_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst5_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst5_xyyy_inst_U16 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sbox_inst5_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst5_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst5_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst5_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst5_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst5_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst5_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst5_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst5_xyyy_inst_U12 ( .A(prince_inst_sin_y[23]), 
        .ZN(prince_inst_sbox_inst5_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst5_xyyy_inst_U11 ( .A1(prince_inst_sin_y[23]), 
        .A2(prince_inst_sbox_inst5_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst5_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst5_t1_sh[3]), .B(
        prince_inst_sbox_inst5_xyyy_inst_n48), .S(
        prince_inst_sbox_inst5_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst5_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst5_xyyy_inst_U9 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sbox_inst5_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst5_xyyy_inst_U8 ( .A1(prince_inst_sin_x[20]), 
        .A2(prince_inst_sin_y[23]), .ZN(prince_inst_sbox_inst5_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst5_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst5_t1_sh[3]), .ZN(prince_inst_sbox_inst5_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst5_xyyy_inst_U6 ( .A1(prince_inst_sin_y[23]), 
        .A2(prince_inst_sbox_inst5_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst5_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst5_xyyy_inst_U4 ( .A(prince_inst_sin_y[21]), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst5_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst5_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst5_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst5_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst5_xyyy_inst_U2 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_x[20]), .ZN(prince_inst_sbox_inst5_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst5_xyyy_inst_U1 ( .A(prince_inst_sin_y[22]), .ZN(
        prince_inst_sbox_inst5_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst5_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U27 ( .A1(prince_inst_sin_y[20]), 
        .A2(prince_inst_sbox_inst5_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst5_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U24 ( .A1(prince_inst_sin_y[20]), 
        .A2(prince_inst_sbox_inst5_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst5_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U21 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst5_yxxx_inst_U19 ( .A(prince_inst_sin_x[23]), 
        .ZN(prince_inst_sbox_inst5_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst5_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst5_yxxx_inst_n52), .B(
        prince_inst_sbox_inst5_yxxx_inst_n51), .S(
        prince_inst_sbox_inst5_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst5_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n53), .A2(prince_inst_sin_x[23]), 
        .ZN(prince_inst_sbox_inst5_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst5_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n48), .A2(prince_inst_sin_y[20]), 
        .ZN(prince_inst_sbox_inst5_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n47), .A2(prince_inst_sin_x[23]), 
        .ZN(prince_inst_sbox_inst5_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U13 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sbox_inst5_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst5_yxxx_inst_n59), .B(
        prince_inst_sbox_inst5_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst5_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst5_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst5_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst5_yxxx_inst_U9 ( .A1(prince_inst_sin_x[21]), 
        .A2(prince_inst_sbox_inst5_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst5_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst5_yxxx_inst_U8 ( .A(prince_inst_sin_x[22]), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst5_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst5_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst5_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst5_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst5_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst5_yxxx_inst_U5 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sbox_inst5_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst5_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst5_yxxx_inst_U4 ( .A(prince_inst_sin_y[20]), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst5_yxxx_inst_U3 ( .A(prince_inst_sin_x[21]), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst5_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst5_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst5_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst5_yxxx_inst_U1 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst5_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst5_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst5_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst5_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst5_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n64), .A3(prince_inst_sin_y[23]), 
        .ZN(prince_inst_sbox_inst5_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst5_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n63), .A2(prince_inst_sin_y[22]), 
        .A3(prince_inst_sin_y[23]), .ZN(prince_inst_sbox_inst5_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst5_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst5_yxyy_inst_n62), .B(
        prince_inst_sbox_inst5_yxyy_inst_n61), .S(prince_inst_sin_y[20]), .Z(
        prince_inst_sbox_inst5_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst5_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst5_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst5_yxyy_inst_n64), .B(
        prince_inst_sbox_inst5_yxyy_inst_n60), .S(
        prince_inst_sbox_inst5_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst5_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst5_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst5_yxyy_inst_n62), .B(
        prince_inst_sbox_inst5_yxyy_inst_n54), .S(
        prince_inst_sbox_inst5_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst5_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst5_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst5_yxyy_inst_n53), .B(
        prince_inst_sbox_inst5_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst5_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst5_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst5_yxyy_inst_n68), .B(
        prince_inst_sbox_inst5_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst5_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U15 ( .A1(prince_inst_sin_y[23]), 
        .A2(prince_inst_sin_y[20]), .ZN(prince_inst_sbox_inst5_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst5_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst5_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst5_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst5_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst5_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst5_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst5_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst5_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n64), .A2(prince_inst_sin_y[22]), 
        .A3(prince_inst_sin_y[20]), .ZN(prince_inst_sbox_inst5_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst5_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U9 ( .A1(prince_inst_sin_y[23]), 
        .A2(prince_inst_sbox_inst5_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst5_yxyy_inst_U8 ( .A1(prince_inst_sin_y[22]), 
        .A2(prince_inst_sbox_inst5_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst5_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst5_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst5_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst5_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst5_yxyy_inst_U5 ( .A(prince_inst_sin_y[20]), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst5_yxyy_inst_U4 ( .A(prince_inst_sin_x[21]), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst5_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst5_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst5_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst5_yxyy_inst_U2 ( .A(prince_inst_sin_y[23]), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst5_yxyy_inst_U1 ( .A(prince_inst_sin_y[22]), .ZN(
        prince_inst_sbox_inst5_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst5_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U29 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sbox_inst5_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst5_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst5_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst5_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n75), .A2(prince_inst_sin_y[23]), 
        .A3(prince_inst_sbox_inst5_yyxy_inst_n70), .A4(prince_inst_sin_x[22]), 
        .ZN(prince_inst_sbox_inst5_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst5_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n69), .A3(prince_inst_sin_y[21]), 
        .A4(prince_inst_sbox_inst5_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst5_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst5_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst5_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst5_yyxy_inst_U23 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_x[22]), .A3(prince_inst_sin_y[20]), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst5_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n69), .A2(prince_inst_sin_y[21]), 
        .A3(prince_inst_sin_y[23]), .ZN(prince_inst_sbox_inst5_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst5_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n75), .A2(prince_inst_sin_x[22]), 
        .A3(prince_inst_sin_y[23]), .ZN(prince_inst_sbox_inst5_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst5_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst5_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst5_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n61), .A2(prince_inst_sin_x[22]), 
        .ZN(prince_inst_sbox_inst5_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst5_yyxy_inst_U18 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_y[23]), .A3(prince_inst_sbox_inst5_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst5_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst5_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst5_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst5_yyxy_inst_U16 ( .A1(prince_inst_sin_y[23]), 
        .A2(prince_inst_sbox_inst5_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst5_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst5_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst5_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n58), .A3(prince_inst_sin_y[20]), 
        .ZN(prince_inst_sbox_inst5_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst5_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst5_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst5_yyxy_inst_U13 ( .A1(prince_inst_sin_y[20]), 
        .A2(prince_inst_sbox_inst5_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst5_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst5_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst5_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst5_yyxy_inst_n54), .B(
        prince_inst_sbox_inst5_yyxy_inst_n55), .S(
        prince_inst_sbox_inst5_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst5_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst5_yyxy_inst_U9 ( .A(prince_inst_sin_x[22]), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n75), .A2(prince_inst_sin_y[23]), 
        .ZN(prince_inst_sbox_inst5_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst5_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst5_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst5_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U5 ( .A1(prince_inst_sin_x[22]), 
        .A2(prince_inst_sbox_inst5_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst5_yyxy_inst_U4 ( .A(prince_inst_sin_y[21]), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst5_yyxy_inst_U3 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sbox_inst5_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst5_yyxy_inst_U2 ( .A(prince_inst_sin_y[20]), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst5_yyxy_inst_U1 ( .A(prince_inst_sin_y[23]), .ZN(
        prince_inst_sbox_inst5_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst5_yyyx_inst_n58), .B(
        prince_inst_sbox_inst5_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst5_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst5_yyyx_inst_n56), .B(
        prince_inst_sbox_inst5_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst5_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst5_yyyx_inst_n54), .B(
        prince_inst_sbox_inst5_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst5_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst5_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst5_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst5_yyyx_inst_U21 ( .A1(prince_inst_sin_x[23]), 
        .A2(prince_inst_sbox_inst5_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst5_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst5_yyyx_inst_U20 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_y[22]), .A3(prince_inst_sbox_inst5_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst5_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst5_yyyx_inst_n50), .B(
        prince_inst_sbox_inst5_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst5_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst5_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n56), .A2(prince_inst_sin_y[22]), 
        .ZN(prince_inst_sbox_inst5_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst5_yyyx_inst_U17 ( .A1(prince_inst_sin_y[21]), 
        .A2(prince_inst_sin_y[20]), .A3(prince_inst_sin_y[22]), .ZN(
        prince_inst_sbox_inst5_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst5_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst5_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst5_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst5_yyyx_inst_U15 ( .A1(prince_inst_sin_x[23]), 
        .A2(prince_inst_sin_y[22]), .A3(prince_inst_sbox_inst5_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst5_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst5_yyyx_inst_U14 ( .A(prince_inst_sin_y[20]), 
        .ZN(prince_inst_sbox_inst5_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n58), .A2(prince_inst_sin_y[21]), 
        .ZN(prince_inst_sbox_inst5_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst5_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst5_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U11 ( .A1(prince_inst_sin_y[20]), 
        .A2(prince_inst_sbox_inst5_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst5_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst5_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst5_yyyx_inst_U9 ( .A1(prince_inst_sin_y[20]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst5_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst5_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst5_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst5_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n45), .A2(prince_inst_sin_y[20]), 
        .A3(prince_inst_sin_y[22]), .ZN(prince_inst_sbox_inst5_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst5_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst5_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst5_yyyx_inst_U4 ( .A1(prince_inst_sin_x[23]), 
        .A2(prince_inst_sin_y[22]), .ZN(prince_inst_sbox_inst5_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst5_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst5_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst5_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst5_yyyx_inst_U2 ( .A(prince_inst_sin_y[21]), .ZN(
        prince_inst_sbox_inst5_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst5_yyyx_inst_U1 ( .A1(prince_inst_sin_y[20]), 
        .A2(prince_inst_sin_x[23]), .ZN(prince_inst_sbox_inst5_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s00_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[0]), .B(prince_inst_sbox_inst5_s0_sh[0]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s01_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[1]), .B(prince_inst_sbox_inst5_s0_sh[1]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s02_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[2]), .B(prince_inst_sbox_inst5_s0_sh[2]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s03_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[3]), .B(prince_inst_sbox_inst5_s0_sh[3]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s04_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[4]), .B(prince_inst_sbox_inst5_s0_sh[4]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s05_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[5]), .B(prince_inst_sbox_inst5_s0_sh[5]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s06_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[6]), .B(prince_inst_sbox_inst5_s0_sh[6]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s07_U1 ( .A(
        prince_inst_sbox_inst5_t0_sh[7]), .B(prince_inst_sbox_inst5_s0_sh[7]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s10_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[0]), .B(prince_inst_sbox_inst5_s1_sh[0]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s11_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[1]), .B(prince_inst_sbox_inst5_s1_sh[1]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s12_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[2]), .B(prince_inst_sbox_inst5_s1_sh[2]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s13_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[3]), .B(prince_inst_sbox_inst5_s1_sh[3]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s14_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[4]), .B(prince_inst_sbox_inst5_s1_sh[4]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s15_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[5]), .B(prince_inst_sbox_inst5_s1_sh[5]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s16_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[6]), .B(prince_inst_sbox_inst5_s1_sh[6]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s17_U1 ( .A(
        prince_inst_sbox_inst5_t1_sh[7]), .B(prince_inst_sbox_inst5_s1_sh[7]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s20_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[0]), .B(prince_inst_sbox_inst5_s2_sh[0]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s21_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[1]), .B(prince_inst_sbox_inst5_s2_sh[1]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s22_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[2]), .B(prince_inst_sbox_inst5_s2_sh[2]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s23_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[3]), .B(prince_inst_sbox_inst5_s2_sh[3]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s24_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[4]), .B(prince_inst_sbox_inst5_s2_sh[4]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s25_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[5]), .B(prince_inst_sbox_inst5_s2_sh[5]), 
        .S(prince_inst_sbox_inst5_n8), .Z(prince_inst_sbox_inst5_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s26_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[6]), .B(prince_inst_sbox_inst5_s2_sh[6]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s27_U1 ( .A(
        prince_inst_sbox_inst5_t2_sh[7]), .B(prince_inst_sbox_inst5_s2_sh[7]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s30_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[0]), .B(prince_inst_sbox_inst5_s3_sh[0]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s31_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[1]), .B(prince_inst_sbox_inst5_s3_sh[1]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s32_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[2]), .B(prince_inst_sbox_inst5_s3_sh[2]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s33_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[3]), .B(prince_inst_sbox_inst5_s3_sh[3]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s34_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[4]), .B(prince_inst_sbox_inst5_s3_sh[4]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s35_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[5]), .B(prince_inst_sbox_inst5_s3_sh[5]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s36_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[6]), .B(prince_inst_sbox_inst5_s3_sh[6]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst5_mux_s37_U1 ( .A(
        prince_inst_sbox_inst5_t3_sh[7]), .B(prince_inst_sbox_inst5_s3_sh[7]), 
        .S(prince_inst_sbox_inst5_n9), .Z(prince_inst_sbox_inst5_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk0_U1 ( .A(r[16]), .B(
        prince_inst_sbox_inst5_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk1_U1 ( .A(r[17]), .B(
        prince_inst_sbox_inst5_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk2_U1 ( .A(r[18]), .B(
        prince_inst_sbox_inst5_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk3_U1 ( .A(r[19]), .B(
        prince_inst_sbox_inst5_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk4_U1 ( .A(r[16]), .B(
        prince_inst_sbox_inst5_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk5_U1 ( .A(r[17]), .B(
        prince_inst_sbox_inst5_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk6_U1 ( .A(r[18]), .B(
        prince_inst_sbox_inst5_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_msk7_U1 ( .A(r[19]), .B(
        prince_inst_sbox_inst5_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst5_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst5_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst5_c_inst0_ax_n5), .ZN(prince_inst_sout_x[20]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst5_c_inst0_y[1]), .B(
        prince_inst_sbox_inst5_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst5_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst5_c_inst0_y[2]), .B(
        prince_inst_sbox_inst5_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst5_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst5_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst5_c_inst0_ay_n5), .ZN(final_y[52]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst5_c_inst0_y[5]), .B(
        prince_inst_sbox_inst5_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst5_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst5_c_inst0_y[6]), .B(
        prince_inst_sbox_inst5_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst5_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk0_U1 ( .A(r[20]), .B(
        prince_inst_sbox_inst5_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk1_U1 ( .A(r[21]), .B(
        prince_inst_sbox_inst5_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk2_U1 ( .A(r[22]), .B(
        prince_inst_sbox_inst5_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk3_U1 ( .A(r[23]), .B(
        prince_inst_sbox_inst5_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk4_U1 ( .A(r[20]), .B(
        prince_inst_sbox_inst5_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk5_U1 ( .A(r[21]), .B(
        prince_inst_sbox_inst5_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk6_U1 ( .A(r[22]), .B(
        prince_inst_sbox_inst5_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_msk7_U1 ( .A(r[23]), .B(
        prince_inst_sbox_inst5_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst5_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst5_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst5_c_inst1_ax_n5), .ZN(prince_inst_sout_x[21]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst5_c_inst1_y[1]), .B(
        prince_inst_sbox_inst5_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst5_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst5_c_inst1_y[2]), .B(
        prince_inst_sbox_inst5_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst5_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst5_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst5_c_inst1_ay_n5), .ZN(final_y[53]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst5_c_inst1_y[5]), .B(
        prince_inst_sbox_inst5_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst5_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst5_c_inst1_y[6]), .B(
        prince_inst_sbox_inst5_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst5_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk0_U1 ( .A(r[24]), .B(
        prince_inst_sbox_inst5_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk1_U1 ( .A(r[25]), .B(
        prince_inst_sbox_inst5_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk2_U1 ( .A(r[26]), .B(
        prince_inst_sbox_inst5_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk3_U1 ( .A(r[27]), .B(
        prince_inst_sbox_inst5_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk4_U1 ( .A(r[24]), .B(
        prince_inst_sbox_inst5_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk5_U1 ( .A(r[25]), .B(
        prince_inst_sbox_inst5_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk6_U1 ( .A(r[26]), .B(
        prince_inst_sbox_inst5_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_msk7_U1 ( .A(r[27]), .B(
        prince_inst_sbox_inst5_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst5_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst5_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst5_c_inst2_ax_n5), .ZN(prince_inst_sout_x[22]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst5_c_inst2_y[1]), .B(
        prince_inst_sbox_inst5_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst5_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst5_c_inst2_y[2]), .B(
        prince_inst_sbox_inst5_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst5_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst5_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst5_c_inst2_ay_n5), .ZN(final_y[54]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst5_c_inst2_y[5]), .B(
        prince_inst_sbox_inst5_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst5_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst5_c_inst2_y[6]), .B(
        prince_inst_sbox_inst5_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst5_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk0_U1 ( .A(r[28]), .B(
        prince_inst_sbox_inst5_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk1_U1 ( .A(r[29]), .B(
        prince_inst_sbox_inst5_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk2_U1 ( .A(r[30]), .B(
        prince_inst_sbox_inst5_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk3_U1 ( .A(r[31]), .B(
        prince_inst_sbox_inst5_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk4_U1 ( .A(r[28]), .B(
        prince_inst_sbox_inst5_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk5_U1 ( .A(r[29]), .B(
        prince_inst_sbox_inst5_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk6_U1 ( .A(r[30]), .B(
        prince_inst_sbox_inst5_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_msk7_U1 ( .A(r[31]), .B(
        prince_inst_sbox_inst5_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst5_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst5_n6), .A3(
        prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst5_n11), .A2(prince_inst_sbox_inst5_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst5_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst5_n11), .ZN(
        prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst5_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst5_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst5_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst5_c_inst3_ax_n5), .ZN(prince_inst_sout_x[23]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst5_c_inst3_y[1]), .B(
        prince_inst_sbox_inst5_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst5_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst5_c_inst3_y[2]), .B(
        prince_inst_sbox_inst5_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst5_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst5_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst5_c_inst3_ay_n5), .ZN(final_y[55]) );
  XNOR2_X1 prince_inst_sbox_inst5_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst5_c_inst3_y[5]), .B(
        prince_inst_sbox_inst5_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst5_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst5_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst5_c_inst3_y[6]), .B(
        prince_inst_sbox_inst5_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst5_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst6_U7 ( .A(prince_inst_sbox_inst6_n12), .ZN(
        prince_inst_sbox_inst6_n11) );
  INV_X1 prince_inst_sbox_inst6_U6 ( .A(prince_inst_n30), .ZN(
        prince_inst_sbox_inst6_n10) );
  INV_X1 prince_inst_sbox_inst6_U5 ( .A(prince_inst_sbox_inst6_n10), .ZN(
        prince_inst_sbox_inst6_n8) );
  INV_X1 prince_inst_sbox_inst6_U4 ( .A(prince_inst_sbox_inst6_n10), .ZN(
        prince_inst_sbox_inst6_n9) );
  INV_X1 prince_inst_sbox_inst6_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst6_n12) );
  INV_X1 prince_inst_sbox_inst6_U2 ( .A(rst), .ZN(prince_inst_sbox_inst6_n7)
         );
  INV_X2 prince_inst_sbox_inst6_U1 ( .A(prince_inst_sbox_inst6_n7), .ZN(
        prince_inst_sbox_inst6_n6) );
  NAND3_X1 prince_inst_sbox_inst6_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n68), .A3(prince_inst_sin_x[24]), 
        .ZN(prince_inst_sbox_inst6_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U25 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sbox_inst6_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst6_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst6_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst6_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst6_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n67), .A2(prince_inst_sin_x[26]), 
        .A3(prince_inst_sin_x[24]), .A4(prince_inst_sin_y[27]), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst6_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n61), .A2(prince_inst_sin_x[25]), 
        .A3(prince_inst_sin_x[26]), .ZN(prince_inst_sbox_inst6_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst6_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n66), .A3(prince_inst_sin_x[25]), 
        .A4(prince_inst_sin_x[24]), .ZN(prince_inst_sbox_inst6_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst6_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst6_xxxy_inst_n59), .B(prince_inst_sin_y[27]), .Z(
        prince_inst_sbox_inst6_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U18 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sin_x[25]), .ZN(prince_inst_sbox_inst6_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst6_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst6_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n65), .A2(prince_inst_sin_x[26]), 
        .ZN(prince_inst_sbox_inst6_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst6_xxxy_inst_U15 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sin_y[27]), .A3(prince_inst_sbox_inst6_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst6_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst6_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst6_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst6_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst6_xxxy_inst_U13 ( .A(prince_inst_sin_x[24]), 
        .B(prince_inst_sin_x[25]), .S(prince_inst_sbox_inst6_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst6_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst6_xxxy_inst_U12 ( .A(prince_inst_sin_y[27]), 
        .ZN(prince_inst_sbox_inst6_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U11 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sin_x[24]), .ZN(prince_inst_sbox_inst6_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst6_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst6_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst6_xxxy_inst_n60), .B(
        prince_inst_sbox_inst6_xxxy_inst_n53), .S(
        prince_inst_sbox_inst6_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst6_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U8 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sbox_inst6_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U7 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sin_y[27]), .ZN(prince_inst_sbox_inst6_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst6_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst6_t1_sh[0]), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst6_xxxy_inst_U5 ( .A(prince_inst_sin_x[26]), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U4 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sbox_inst6_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst6_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst6_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst6_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst6_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst6_xxxy_inst_U2 ( .A(prince_inst_sin_x[24]), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst6_xxxy_inst_U1 ( .A(prince_inst_sin_x[25]), .ZN(
        prince_inst_sbox_inst6_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst6_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst6_t1_sh[1]), .B(
        prince_inst_sbox_inst6_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst6_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst6_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst6_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst6_xxyx_inst_n52), .B(
        prince_inst_sbox_inst6_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst6_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U23 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst6_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst6_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n48), .A2(prince_inst_sin_x[27]), 
        .A3(prince_inst_sin_x[24]), .ZN(prince_inst_sbox_inst6_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst6_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst6_xxyx_inst_U18 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sbox_inst6_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst6_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst6_xxyx_inst_U16 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sin_x[24]), .A3(prince_inst_sbox_inst6_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst6_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst6_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n46), .A2(prince_inst_sin_x[27]), 
        .A3(prince_inst_sin_x[25]), .ZN(prince_inst_sbox_inst6_xxyx_inst_n44)
         );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst6_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst6_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst6_xxyx_inst_n54), .B(
        prince_inst_sbox_inst6_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst6_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U12 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sin_y[26]), .ZN(prince_inst_sbox_inst6_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst6_xxyx_inst_U11 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sbox_inst6_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst6_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst6_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst6_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst6_xxyx_inst_U10 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst6_xxyx_inst_U9 ( .A1(prince_inst_sin_x[27]), 
        .A2(prince_inst_sbox_inst6_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst6_xxyx_inst_U8 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sbox_inst6_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst6_xxyx_inst_U7 ( .A(prince_inst_sin_y[26]), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst6_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst6_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst6_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n53), .A2(prince_inst_sin_x[25]), 
        .A3(prince_inst_sin_y[26]), .A4(prince_inst_sin_x[24]), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst6_xxyx_inst_U4 ( .A(prince_inst_sin_x[27]), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst6_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst6_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst6_xxyx_inst_n43), .A3(prince_inst_sin_x[27]), 
        .A4(prince_inst_sin_y[26]), .ZN(prince_inst_sbox_inst6_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst6_xxyx_inst_U2 ( .A(prince_inst_sin_x[24]), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst6_xxyx_inst_U1 ( .A(prince_inst_sin_x[25]), .ZN(
        prince_inst_sbox_inst6_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst6_xyxx_inst_n74), .B(
        prince_inst_sbox_inst6_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst6_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst6_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst6_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst6_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U26 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sbox_inst6_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U25 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst6_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst6_xyxx_inst_n72), .B(
        prince_inst_sbox_inst6_s0_sh[2]), .S(
        prince_inst_sbox_inst6_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst6_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst6_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n74), .A2(prince_inst_sin_x[27]), 
        .ZN(prince_inst_sbox_inst6_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst6_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U21 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sbox_inst6_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst6_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst6_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst6_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst6_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst6_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst6_xyxx_inst_U15 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_x[24]), .ZN(prince_inst_sbox_inst6_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst6_xyxx_inst_U13 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U12 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_x[26]), .ZN(prince_inst_sbox_inst6_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst6_xyxx_inst_n58), .B(
        prince_inst_sbox_inst6_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst6_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst6_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst6_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst6_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst6_xyxx_inst_U9 ( .A(prince_inst_sin_x[27]), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst6_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n54), .A2(prince_inst_sin_x[24]), 
        .ZN(prince_inst_sbox_inst6_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst6_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst6_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst6_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst6_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst6_xyxx_inst_U5 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sbox_inst6_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst6_xyxx_inst_U4 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst6_xyxx_inst_U3 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sbox_inst6_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst6_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst6_xyxx_inst_U2 ( .A(prince_inst_sin_y[25]), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst6_xyxx_inst_U1 ( .A(prince_inst_sin_x[26]), .ZN(
        prince_inst_sbox_inst6_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst6_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst6_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst6_xyyy_inst_n59), .B(
        prince_inst_sbox_inst6_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst6_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst6_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst6_xyyy_inst_U25 ( .A1(prince_inst_sin_y[26]), 
        .A2(prince_inst_sin_y[27]), .A3(prince_inst_sbox_inst6_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst6_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U24 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sbox_inst6_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U23 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sbox_inst6_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst6_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst6_xyyy_inst_U19 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sin_y[26]), .A3(prince_inst_sbox_inst6_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst6_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst6_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst6_xyyy_inst_n49), .B(
        prince_inst_sbox_inst6_xyyy_inst_n48), .S(
        prince_inst_sbox_inst6_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst6_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst6_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst6_xyyy_inst_U16 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sbox_inst6_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst6_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst6_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst6_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst6_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst6_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst6_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst6_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst6_xyyy_inst_U12 ( .A(prince_inst_sin_y[27]), 
        .ZN(prince_inst_sbox_inst6_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst6_xyyy_inst_U11 ( .A1(prince_inst_sin_y[27]), 
        .A2(prince_inst_sbox_inst6_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst6_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst6_t1_sh[3]), .B(
        prince_inst_sbox_inst6_xyyy_inst_n48), .S(
        prince_inst_sbox_inst6_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst6_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst6_xyyy_inst_U9 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sbox_inst6_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst6_xyyy_inst_U8 ( .A1(prince_inst_sin_x[24]), 
        .A2(prince_inst_sin_y[27]), .ZN(prince_inst_sbox_inst6_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst6_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst6_t1_sh[3]), .ZN(prince_inst_sbox_inst6_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst6_xyyy_inst_U6 ( .A1(prince_inst_sin_y[27]), 
        .A2(prince_inst_sbox_inst6_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst6_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst6_xyyy_inst_U4 ( .A(prince_inst_sin_y[25]), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst6_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst6_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst6_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst6_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst6_xyyy_inst_U2 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_x[24]), .ZN(prince_inst_sbox_inst6_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst6_xyyy_inst_U1 ( .A(prince_inst_sin_y[26]), .ZN(
        prince_inst_sbox_inst6_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst6_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U27 ( .A1(prince_inst_sin_y[24]), 
        .A2(prince_inst_sbox_inst6_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst6_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U24 ( .A1(prince_inst_sin_y[24]), 
        .A2(prince_inst_sbox_inst6_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst6_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U21 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst6_yxxx_inst_U19 ( .A(prince_inst_sin_x[27]), 
        .ZN(prince_inst_sbox_inst6_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst6_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst6_yxxx_inst_n52), .B(
        prince_inst_sbox_inst6_yxxx_inst_n51), .S(
        prince_inst_sbox_inst6_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst6_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n53), .A2(prince_inst_sin_x[27]), 
        .ZN(prince_inst_sbox_inst6_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst6_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n48), .A2(prince_inst_sin_y[24]), 
        .ZN(prince_inst_sbox_inst6_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n47), .A2(prince_inst_sin_x[27]), 
        .ZN(prince_inst_sbox_inst6_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U13 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sbox_inst6_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst6_yxxx_inst_n59), .B(
        prince_inst_sbox_inst6_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst6_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst6_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst6_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst6_yxxx_inst_U9 ( .A1(prince_inst_sin_x[25]), 
        .A2(prince_inst_sbox_inst6_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst6_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst6_yxxx_inst_U8 ( .A(prince_inst_sin_x[26]), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst6_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst6_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst6_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst6_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst6_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst6_yxxx_inst_U5 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sbox_inst6_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst6_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst6_yxxx_inst_U4 ( .A(prince_inst_sin_y[24]), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst6_yxxx_inst_U3 ( .A(prince_inst_sin_x[25]), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst6_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst6_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst6_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst6_yxxx_inst_U1 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst6_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst6_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst6_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst6_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst6_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n64), .A3(prince_inst_sin_y[27]), 
        .ZN(prince_inst_sbox_inst6_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst6_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n63), .A2(prince_inst_sin_y[26]), 
        .A3(prince_inst_sin_y[27]), .ZN(prince_inst_sbox_inst6_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst6_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst6_yxyy_inst_n62), .B(
        prince_inst_sbox_inst6_yxyy_inst_n61), .S(prince_inst_sin_y[24]), .Z(
        prince_inst_sbox_inst6_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst6_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst6_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst6_yxyy_inst_n64), .B(
        prince_inst_sbox_inst6_yxyy_inst_n60), .S(
        prince_inst_sbox_inst6_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst6_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst6_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst6_yxyy_inst_n62), .B(
        prince_inst_sbox_inst6_yxyy_inst_n54), .S(
        prince_inst_sbox_inst6_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst6_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst6_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst6_yxyy_inst_n53), .B(
        prince_inst_sbox_inst6_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst6_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst6_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst6_yxyy_inst_n68), .B(
        prince_inst_sbox_inst6_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst6_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U15 ( .A1(prince_inst_sin_y[27]), 
        .A2(prince_inst_sin_y[24]), .ZN(prince_inst_sbox_inst6_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst6_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst6_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst6_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst6_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst6_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst6_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst6_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst6_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n64), .A2(prince_inst_sin_y[26]), 
        .A3(prince_inst_sin_y[24]), .ZN(prince_inst_sbox_inst6_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst6_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U9 ( .A1(prince_inst_sin_y[27]), 
        .A2(prince_inst_sbox_inst6_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst6_yxyy_inst_U8 ( .A1(prince_inst_sin_y[26]), 
        .A2(prince_inst_sbox_inst6_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst6_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst6_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst6_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst6_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst6_yxyy_inst_U5 ( .A(prince_inst_sin_y[24]), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst6_yxyy_inst_U4 ( .A(prince_inst_sin_x[25]), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst6_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst6_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst6_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst6_yxyy_inst_U2 ( .A(prince_inst_sin_y[27]), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst6_yxyy_inst_U1 ( .A(prince_inst_sin_y[26]), .ZN(
        prince_inst_sbox_inst6_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst6_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U29 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sbox_inst6_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst6_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst6_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst6_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n75), .A2(prince_inst_sin_y[27]), 
        .A3(prince_inst_sbox_inst6_yyxy_inst_n70), .A4(prince_inst_sin_x[26]), 
        .ZN(prince_inst_sbox_inst6_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst6_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n69), .A3(prince_inst_sin_y[25]), 
        .A4(prince_inst_sbox_inst6_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst6_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst6_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst6_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst6_yyxy_inst_U23 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_x[26]), .A3(prince_inst_sin_y[24]), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst6_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n69), .A2(prince_inst_sin_y[25]), 
        .A3(prince_inst_sin_y[27]), .ZN(prince_inst_sbox_inst6_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst6_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n75), .A2(prince_inst_sin_x[26]), 
        .A3(prince_inst_sin_y[27]), .ZN(prince_inst_sbox_inst6_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst6_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst6_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst6_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n61), .A2(prince_inst_sin_x[26]), 
        .ZN(prince_inst_sbox_inst6_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst6_yyxy_inst_U18 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_y[27]), .A3(prince_inst_sbox_inst6_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst6_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst6_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst6_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst6_yyxy_inst_U16 ( .A1(prince_inst_sin_y[27]), 
        .A2(prince_inst_sbox_inst6_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst6_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst6_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst6_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n58), .A3(prince_inst_sin_y[24]), 
        .ZN(prince_inst_sbox_inst6_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst6_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst6_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst6_yyxy_inst_U13 ( .A1(prince_inst_sin_y[24]), 
        .A2(prince_inst_sbox_inst6_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst6_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst6_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst6_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst6_yyxy_inst_n54), .B(
        prince_inst_sbox_inst6_yyxy_inst_n55), .S(
        prince_inst_sbox_inst6_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst6_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst6_yyxy_inst_U9 ( .A(prince_inst_sin_x[26]), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n75), .A2(prince_inst_sin_y[27]), 
        .ZN(prince_inst_sbox_inst6_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst6_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst6_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst6_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U5 ( .A1(prince_inst_sin_x[26]), 
        .A2(prince_inst_sbox_inst6_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst6_yyxy_inst_U4 ( .A(prince_inst_sin_y[25]), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst6_yyxy_inst_U3 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sbox_inst6_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst6_yyxy_inst_U2 ( .A(prince_inst_sin_y[24]), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst6_yyxy_inst_U1 ( .A(prince_inst_sin_y[27]), .ZN(
        prince_inst_sbox_inst6_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst6_yyyx_inst_n58), .B(
        prince_inst_sbox_inst6_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst6_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst6_yyyx_inst_n56), .B(
        prince_inst_sbox_inst6_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst6_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst6_yyyx_inst_n54), .B(
        prince_inst_sbox_inst6_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst6_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst6_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst6_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst6_yyyx_inst_U21 ( .A1(prince_inst_sin_x[27]), 
        .A2(prince_inst_sbox_inst6_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst6_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst6_yyyx_inst_U20 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_y[26]), .A3(prince_inst_sbox_inst6_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst6_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst6_yyyx_inst_n50), .B(
        prince_inst_sbox_inst6_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst6_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst6_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n56), .A2(prince_inst_sin_y[26]), 
        .ZN(prince_inst_sbox_inst6_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst6_yyyx_inst_U17 ( .A1(prince_inst_sin_y[25]), 
        .A2(prince_inst_sin_y[24]), .A3(prince_inst_sin_y[26]), .ZN(
        prince_inst_sbox_inst6_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst6_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst6_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst6_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst6_yyyx_inst_U15 ( .A1(prince_inst_sin_x[27]), 
        .A2(prince_inst_sin_y[26]), .A3(prince_inst_sbox_inst6_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst6_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst6_yyyx_inst_U14 ( .A(prince_inst_sin_y[24]), 
        .ZN(prince_inst_sbox_inst6_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n58), .A2(prince_inst_sin_y[25]), 
        .ZN(prince_inst_sbox_inst6_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst6_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst6_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U11 ( .A1(prince_inst_sin_y[24]), 
        .A2(prince_inst_sbox_inst6_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst6_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst6_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst6_yyyx_inst_U9 ( .A1(prince_inst_sin_y[24]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst6_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst6_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst6_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst6_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n45), .A2(prince_inst_sin_y[24]), 
        .A3(prince_inst_sin_y[26]), .ZN(prince_inst_sbox_inst6_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst6_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst6_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst6_yyyx_inst_U4 ( .A1(prince_inst_sin_x[27]), 
        .A2(prince_inst_sin_y[26]), .ZN(prince_inst_sbox_inst6_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst6_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst6_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst6_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst6_yyyx_inst_U2 ( .A(prince_inst_sin_y[25]), .ZN(
        prince_inst_sbox_inst6_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst6_yyyx_inst_U1 ( .A1(prince_inst_sin_y[24]), 
        .A2(prince_inst_sin_x[27]), .ZN(prince_inst_sbox_inst6_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s00_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[0]), .B(prince_inst_sbox_inst6_s0_sh[0]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s01_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[1]), .B(prince_inst_sbox_inst6_s0_sh[1]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s02_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[2]), .B(prince_inst_sbox_inst6_s0_sh[2]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s03_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[3]), .B(prince_inst_sbox_inst6_s0_sh[3]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s04_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[4]), .B(prince_inst_sbox_inst6_s0_sh[4]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s05_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[5]), .B(prince_inst_sbox_inst6_s0_sh[5]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s06_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[6]), .B(prince_inst_sbox_inst6_s0_sh[6]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s07_U1 ( .A(
        prince_inst_sbox_inst6_t0_sh[7]), .B(prince_inst_sbox_inst6_s0_sh[7]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s10_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[0]), .B(prince_inst_sbox_inst6_s1_sh[0]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s11_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[1]), .B(prince_inst_sbox_inst6_s1_sh[1]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s12_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[2]), .B(prince_inst_sbox_inst6_s1_sh[2]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s13_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[3]), .B(prince_inst_sbox_inst6_s1_sh[3]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s14_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[4]), .B(prince_inst_sbox_inst6_s1_sh[4]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s15_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[5]), .B(prince_inst_sbox_inst6_s1_sh[5]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s16_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[6]), .B(prince_inst_sbox_inst6_s1_sh[6]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s17_U1 ( .A(
        prince_inst_sbox_inst6_t1_sh[7]), .B(prince_inst_sbox_inst6_s1_sh[7]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s20_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[0]), .B(prince_inst_sbox_inst6_s2_sh[0]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s21_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[1]), .B(prince_inst_sbox_inst6_s2_sh[1]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s22_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[2]), .B(prince_inst_sbox_inst6_s2_sh[2]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s23_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[3]), .B(prince_inst_sbox_inst6_s2_sh[3]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s24_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[4]), .B(prince_inst_sbox_inst6_s2_sh[4]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s25_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[5]), .B(prince_inst_sbox_inst6_s2_sh[5]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s26_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[6]), .B(prince_inst_sbox_inst6_s2_sh[6]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s27_U1 ( .A(
        prince_inst_sbox_inst6_t2_sh[7]), .B(prince_inst_sbox_inst6_s2_sh[7]), 
        .S(prince_inst_sbox_inst6_n8), .Z(prince_inst_sbox_inst6_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s30_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[0]), .B(prince_inst_sbox_inst6_s3_sh[0]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s31_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[1]), .B(prince_inst_sbox_inst6_s3_sh[1]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s32_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[2]), .B(prince_inst_sbox_inst6_s3_sh[2]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s33_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[3]), .B(prince_inst_sbox_inst6_s3_sh[3]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s34_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[4]), .B(prince_inst_sbox_inst6_s3_sh[4]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s35_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[5]), .B(prince_inst_sbox_inst6_s3_sh[5]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s36_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[6]), .B(prince_inst_sbox_inst6_s3_sh[6]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst6_mux_s37_U1 ( .A(
        prince_inst_sbox_inst6_t3_sh[7]), .B(prince_inst_sbox_inst6_s3_sh[7]), 
        .S(prince_inst_sbox_inst6_n9), .Z(prince_inst_sbox_inst6_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk0_U1 ( .A(r[32]), .B(
        prince_inst_sbox_inst6_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk1_U1 ( .A(r[33]), .B(
        prince_inst_sbox_inst6_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk2_U1 ( .A(r[34]), .B(
        prince_inst_sbox_inst6_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk3_U1 ( .A(r[35]), .B(
        prince_inst_sbox_inst6_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk4_U1 ( .A(r[32]), .B(
        prince_inst_sbox_inst6_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk5_U1 ( .A(r[33]), .B(
        prince_inst_sbox_inst6_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk6_U1 ( .A(r[34]), .B(
        prince_inst_sbox_inst6_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_msk7_U1 ( .A(r[35]), .B(
        prince_inst_sbox_inst6_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst6_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst6_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst6_c_inst0_ax_n5), .ZN(prince_inst_sout_x[24]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst6_c_inst0_y[1]), .B(
        prince_inst_sbox_inst6_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst6_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst6_c_inst0_y[2]), .B(
        prince_inst_sbox_inst6_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst6_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst6_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst6_c_inst0_ay_n5), .ZN(final_y[40]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst6_c_inst0_y[5]), .B(
        prince_inst_sbox_inst6_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst6_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst6_c_inst0_y[6]), .B(
        prince_inst_sbox_inst6_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst6_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk0_U1 ( .A(r[36]), .B(
        prince_inst_sbox_inst6_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk1_U1 ( .A(r[37]), .B(
        prince_inst_sbox_inst6_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk2_U1 ( .A(r[38]), .B(
        prince_inst_sbox_inst6_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk3_U1 ( .A(r[39]), .B(
        prince_inst_sbox_inst6_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk4_U1 ( .A(r[36]), .B(
        prince_inst_sbox_inst6_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk5_U1 ( .A(r[37]), .B(
        prince_inst_sbox_inst6_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk6_U1 ( .A(r[38]), .B(
        prince_inst_sbox_inst6_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_msk7_U1 ( .A(r[39]), .B(
        prince_inst_sbox_inst6_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst6_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst6_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst6_c_inst1_ax_n5), .ZN(prince_inst_sout_x[25]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst6_c_inst1_y[1]), .B(
        prince_inst_sbox_inst6_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst6_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst6_c_inst1_y[2]), .B(
        prince_inst_sbox_inst6_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst6_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst6_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst6_c_inst1_ay_n5), .ZN(final_y[41]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst6_c_inst1_y[5]), .B(
        prince_inst_sbox_inst6_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst6_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst6_c_inst1_y[6]), .B(
        prince_inst_sbox_inst6_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst6_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk0_U1 ( .A(r[40]), .B(
        prince_inst_sbox_inst6_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk1_U1 ( .A(r[41]), .B(
        prince_inst_sbox_inst6_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk2_U1 ( .A(r[42]), .B(
        prince_inst_sbox_inst6_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk3_U1 ( .A(r[43]), .B(
        prince_inst_sbox_inst6_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk4_U1 ( .A(r[40]), .B(
        prince_inst_sbox_inst6_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk5_U1 ( .A(r[41]), .B(
        prince_inst_sbox_inst6_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk6_U1 ( .A(r[42]), .B(
        prince_inst_sbox_inst6_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_msk7_U1 ( .A(r[43]), .B(
        prince_inst_sbox_inst6_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst6_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst6_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst6_c_inst2_ax_n5), .ZN(prince_inst_sout_x[26]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst6_c_inst2_y[1]), .B(
        prince_inst_sbox_inst6_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst6_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst6_c_inst2_y[2]), .B(
        prince_inst_sbox_inst6_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst6_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst6_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst6_c_inst2_ay_n5), .ZN(final_y[42]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst6_c_inst2_y[5]), .B(
        prince_inst_sbox_inst6_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst6_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst6_c_inst2_y[6]), .B(
        prince_inst_sbox_inst6_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst6_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk0_U1 ( .A(r[44]), .B(
        prince_inst_sbox_inst6_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk1_U1 ( .A(r[45]), .B(
        prince_inst_sbox_inst6_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk2_U1 ( .A(r[46]), .B(
        prince_inst_sbox_inst6_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk3_U1 ( .A(r[47]), .B(
        prince_inst_sbox_inst6_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk4_U1 ( .A(r[44]), .B(
        prince_inst_sbox_inst6_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk5_U1 ( .A(r[45]), .B(
        prince_inst_sbox_inst6_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk6_U1 ( .A(r[46]), .B(
        prince_inst_sbox_inst6_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_msk7_U1 ( .A(r[47]), .B(
        prince_inst_sbox_inst6_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst6_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst6_n6), .A3(
        prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst6_n11), .A2(prince_inst_sbox_inst6_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst6_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst6_n11), .ZN(
        prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst6_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst6_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst6_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst6_c_inst3_ax_n5), .ZN(prince_inst_sout_x[27]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst6_c_inst3_y[1]), .B(
        prince_inst_sbox_inst6_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst6_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst6_c_inst3_y[2]), .B(
        prince_inst_sbox_inst6_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst6_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst6_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst6_c_inst3_ay_n5), .ZN(final_y[43]) );
  XNOR2_X1 prince_inst_sbox_inst6_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst6_c_inst3_y[5]), .B(
        prince_inst_sbox_inst6_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst6_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst6_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst6_c_inst3_y[6]), .B(
        prince_inst_sbox_inst6_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst6_c_inst3_ay_n6) );
  INV_X1 prince_inst_sbox_inst7_U5 ( .A(prince_inst_n26), .ZN(
        prince_inst_sbox_inst7_n10) );
  INV_X1 prince_inst_sbox_inst7_U4 ( .A(prince_inst_sbox_inst7_n10), .ZN(
        prince_inst_sbox_inst7_n8) );
  INV_X1 prince_inst_sbox_inst7_U3 ( .A(prince_inst_sbox_inst7_n10), .ZN(
        prince_inst_sbox_inst7_n9) );
  INV_X1 prince_inst_sbox_inst7_U2 ( .A(rst), .ZN(prince_inst_sbox_inst7_n7)
         );
  INV_X2 prince_inst_sbox_inst7_U1 ( .A(prince_inst_sbox_inst7_n7), .ZN(
        prince_inst_sbox_inst7_n6) );
  NAND3_X1 prince_inst_sbox_inst7_xxxy_inst_U28 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n70), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n69), .A3(prince_inst_sin_x[28]), 
        .ZN(prince_inst_sbox_inst7_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n67), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n69) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U26 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n70) );
  NAND3_X1 prince_inst_sbox_inst7_xxxy_inst_U25 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n65), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n64), .A3(
        prince_inst_sbox_inst7_xxxy_inst_n63), .ZN(
        prince_inst_sbox_inst7_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst7_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n68), .A2(prince_inst_sin_x[30]), 
        .A3(prince_inst_sin_x[28]), .A4(prince_inst_sin_y[31]), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n63) );
  NAND3_X1 prince_inst_sbox_inst7_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n62), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n61), .A3(prince_inst_sin_x[30]), 
        .ZN(prince_inst_sbox_inst7_xxxy_inst_n64) );
  NAND4_X1 prince_inst_sbox_inst7_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n67), .A3(
        prince_inst_sbox_inst7_xxxy_inst_n61), .A4(prince_inst_sin_x[28]), 
        .ZN(prince_inst_sbox_inst7_xxxy_inst_n65) );
  XOR2_X1 prince_inst_sbox_inst7_xxxy_inst_U21 ( .A(
        prince_inst_sbox_inst7_xxxy_inst_n59), .B(prince_inst_sin_y[31]), .Z(
        prince_inst_sbox_inst7_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U20 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U19 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n58) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U18 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst7_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst7_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n66), .A2(prince_inst_sin_x[30]), 
        .ZN(prince_inst_sbox_inst7_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst7_xxxy_inst_U16 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sin_y[31]), .A3(prince_inst_sbox_inst7_xxxy_inst_n68), 
        .ZN(prince_inst_sbox_inst7_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst7_xxxy_inst_U15 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst7_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst7_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst7_xxxy_inst_U14 ( .A(prince_inst_sin_x[28]), 
        .B(prince_inst_sbox_inst7_xxxy_inst_n61), .S(
        prince_inst_sbox_inst7_xxxy_inst_n67), .Z(
        prince_inst_sbox_inst7_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst7_xxxy_inst_U13 ( .A(prince_inst_sin_y[31]), 
        .ZN(prince_inst_sbox_inst7_xxxy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U12 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n61), .A2(prince_inst_sin_x[28]), 
        .ZN(prince_inst_sbox_inst7_xxxy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U11 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst7_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst7_xxxy_inst_U10 ( .A(
        prince_inst_sbox_inst7_xxxy_inst_n60), .B(
        prince_inst_sbox_inst7_xxxy_inst_n53), .S(
        prince_inst_sbox_inst7_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst7_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U9 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sbox_inst7_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U8 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n61), .A2(prince_inst_sin_y[31]), 
        .ZN(prince_inst_sbox_inst7_xxxy_inst_n66) );
  INV_X1 prince_inst_sbox_inst7_xxxy_inst_U7 ( .A(
        prince_inst_sbox_inst7_xxxy_inst_n68), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst7_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst7_t1_sh[0]), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst7_xxxy_inst_U5 ( .A(prince_inst_sin_x[30]), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U4 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst7_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst7_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst7_xxxy_inst_n68), .A2(
        prince_inst_sbox_inst7_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst7_xxxy_inst_U2 ( .A(prince_inst_sin_x[28]), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n62) );
  INV_X1 prince_inst_sbox_inst7_xxxy_inst_U1 ( .A(prince_inst_sin_x[29]), .ZN(
        prince_inst_sbox_inst7_xxxy_inst_n68) );
  XOR2_X1 prince_inst_sbox_inst7_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst7_t1_sh[1]), .B(
        prince_inst_sbox_inst7_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst7_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst7_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst7_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst7_xxyx_inst_n52), .B(
        prince_inst_sbox_inst7_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst7_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U23 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst7_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst7_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n48), .A2(prince_inst_sin_x[31]), 
        .A3(prince_inst_sin_x[28]), .ZN(prince_inst_sbox_inst7_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst7_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst7_xxyx_inst_U18 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sbox_inst7_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst7_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst7_xxyx_inst_U16 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sin_x[28]), .A3(prince_inst_sbox_inst7_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst7_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst7_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n46), .A2(prince_inst_sin_x[31]), 
        .A3(prince_inst_sin_x[29]), .ZN(prince_inst_sbox_inst7_xxyx_inst_n44)
         );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst7_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst7_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst7_xxyx_inst_n54), .B(
        prince_inst_sbox_inst7_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst7_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U12 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sin_y[30]), .ZN(prince_inst_sbox_inst7_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst7_xxyx_inst_U11 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sbox_inst7_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst7_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst7_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst7_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst7_xxyx_inst_U10 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst7_xxyx_inst_U9 ( .A1(prince_inst_sin_x[31]), 
        .A2(prince_inst_sbox_inst7_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst7_xxyx_inst_U8 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sbox_inst7_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst7_xxyx_inst_U7 ( .A(prince_inst_sin_y[30]), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst7_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst7_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst7_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n53), .A2(prince_inst_sin_x[29]), 
        .A3(prince_inst_sin_y[30]), .A4(prince_inst_sin_x[28]), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst7_xxyx_inst_U4 ( .A(prince_inst_sin_x[31]), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst7_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst7_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst7_xxyx_inst_n43), .A3(prince_inst_sin_x[31]), 
        .A4(prince_inst_sin_y[30]), .ZN(prince_inst_sbox_inst7_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst7_xxyx_inst_U2 ( .A(prince_inst_sin_x[28]), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst7_xxyx_inst_U1 ( .A(prince_inst_sin_x[29]), .ZN(
        prince_inst_sbox_inst7_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst7_xyxx_inst_n74), .B(
        prince_inst_sbox_inst7_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst7_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst7_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst7_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst7_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U26 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sbox_inst7_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U25 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst7_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst7_xyxx_inst_n72), .B(
        prince_inst_sbox_inst7_s0_sh[2]), .S(
        prince_inst_sbox_inst7_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst7_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst7_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n74), .A2(prince_inst_sin_x[31]), 
        .ZN(prince_inst_sbox_inst7_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst7_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U21 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst7_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst7_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst7_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst7_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst7_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst7_xyxx_inst_U15 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_x[28]), .ZN(prince_inst_sbox_inst7_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst7_xyxx_inst_U13 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U12 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_x[30]), .ZN(prince_inst_sbox_inst7_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst7_xyxx_inst_n58), .B(
        prince_inst_sbox_inst7_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst7_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst7_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst7_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst7_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst7_xyxx_inst_U9 ( .A(prince_inst_sin_x[31]), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst7_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n54), .A2(prince_inst_sin_x[28]), 
        .ZN(prince_inst_sbox_inst7_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst7_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst7_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst7_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst7_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst7_xyxx_inst_U5 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst7_xyxx_inst_U4 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst7_xyxx_inst_U3 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sbox_inst7_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst7_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst7_xyxx_inst_U2 ( .A(prince_inst_sin_y[29]), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst7_xyxx_inst_U1 ( .A(prince_inst_sin_x[30]), .ZN(
        prince_inst_sbox_inst7_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst7_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst7_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst7_xyyy_inst_n59), .B(
        prince_inst_sbox_inst7_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst7_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst7_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst7_xyyy_inst_U25 ( .A1(prince_inst_sin_y[30]), 
        .A2(prince_inst_sin_y[31]), .A3(prince_inst_sbox_inst7_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst7_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U24 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sbox_inst7_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U23 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sbox_inst7_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst7_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst7_xyyy_inst_U19 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sin_y[30]), .A3(prince_inst_sbox_inst7_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst7_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst7_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst7_xyyy_inst_n49), .B(
        prince_inst_sbox_inst7_xyyy_inst_n48), .S(
        prince_inst_sbox_inst7_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst7_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst7_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst7_xyyy_inst_U16 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sbox_inst7_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst7_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst7_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst7_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst7_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst7_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst7_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst7_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst7_xyyy_inst_U12 ( .A(prince_inst_sin_y[31]), 
        .ZN(prince_inst_sbox_inst7_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst7_xyyy_inst_U11 ( .A1(prince_inst_sin_y[31]), 
        .A2(prince_inst_sbox_inst7_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst7_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst7_t1_sh[3]), .B(
        prince_inst_sbox_inst7_xyyy_inst_n48), .S(
        prince_inst_sbox_inst7_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst7_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst7_xyyy_inst_U9 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sbox_inst7_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst7_xyyy_inst_U8 ( .A1(prince_inst_sin_x[28]), 
        .A2(prince_inst_sin_y[31]), .ZN(prince_inst_sbox_inst7_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst7_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst7_t1_sh[3]), .ZN(prince_inst_sbox_inst7_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst7_xyyy_inst_U6 ( .A1(prince_inst_sin_y[31]), 
        .A2(prince_inst_sbox_inst7_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst7_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst7_xyyy_inst_U4 ( .A(prince_inst_sin_y[29]), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst7_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst7_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst7_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst7_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst7_xyyy_inst_U2 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_x[28]), .ZN(prince_inst_sbox_inst7_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst7_xyyy_inst_U1 ( .A(prince_inst_sin_y[30]), .ZN(
        prince_inst_sbox_inst7_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst7_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U27 ( .A1(prince_inst_sin_y[28]), 
        .A2(prince_inst_sbox_inst7_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst7_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U24 ( .A1(prince_inst_sin_y[28]), 
        .A2(prince_inst_sbox_inst7_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst7_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U21 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst7_yxxx_inst_U19 ( .A(prince_inst_sin_x[31]), 
        .ZN(prince_inst_sbox_inst7_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst7_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst7_yxxx_inst_n52), .B(
        prince_inst_sbox_inst7_yxxx_inst_n51), .S(
        prince_inst_sbox_inst7_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst7_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n53), .A2(prince_inst_sin_x[31]), 
        .ZN(prince_inst_sbox_inst7_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst7_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n48), .A2(prince_inst_sin_y[28]), 
        .ZN(prince_inst_sbox_inst7_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n47), .A2(prince_inst_sin_x[31]), 
        .ZN(prince_inst_sbox_inst7_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U13 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sbox_inst7_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst7_yxxx_inst_n59), .B(
        prince_inst_sbox_inst7_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst7_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst7_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst7_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst7_yxxx_inst_U9 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst7_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst7_yxxx_inst_U8 ( .A(
        prince_inst_sbox_inst7_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n51) );
  OR2_X1 prince_inst_sbox_inst7_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst7_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst7_yxxx_inst_U6 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sbox_inst7_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst7_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst7_yxxx_inst_U5 ( .A(prince_inst_sin_x[30]), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n55) );
  INV_X1 prince_inst_sbox_inst7_yxxx_inst_U4 ( .A(prince_inst_sin_y[28]), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst7_yxxx_inst_U3 ( .A1(
        prince_inst_sbox_inst7_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst7_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst7_yxxx_inst_U2 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_yxxx_inst_n45)
         );
  INV_X1 prince_inst_sbox_inst7_yxxx_inst_U1 ( .A(prince_inst_sin_x[29]), .ZN(
        prince_inst_sbox_inst7_yxxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n67), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n66), .ZN(
        prince_inst_sbox_inst7_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst7_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n66), .A3(
        prince_inst_sbox_inst7_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst7_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst7_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n64), .A2(prince_inst_sin_x[29]), 
        .A3(prince_inst_sin_y[31]), .ZN(prince_inst_sbox_inst7_yxyy_inst_n66)
         );
  NAND3_X1 prince_inst_sbox_inst7_yxyy_inst_U24 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n63), .A2(prince_inst_sin_y[30]), 
        .A3(prince_inst_sin_y[31]), .ZN(prince_inst_sbox_inst7_yxyy_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst7_yxyy_inst_U23 ( .A(
        prince_inst_sbox_inst7_yxyy_inst_n62), .B(
        prince_inst_sbox_inst7_yxyy_inst_n61), .S(prince_inst_sin_y[28]), .Z(
        prince_inst_sbox_inst7_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst7_yxyy_inst_U22 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n64), .A2(prince_inst_sin_x[29]), 
        .ZN(prince_inst_sbox_inst7_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst7_yxyy_inst_U21 ( .A(prince_inst_sin_x[29]), 
        .B(prince_inst_sbox_inst7_yxyy_inst_n60), .S(
        prince_inst_sbox_inst7_yxyy_inst_n64), .Z(
        prince_inst_sbox_inst7_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U18 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst7_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst7_yxyy_inst_n62), .B(
        prince_inst_sbox_inst7_yxyy_inst_n54), .S(
        prince_inst_sbox_inst7_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst7_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst7_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst7_yxyy_inst_n53), .B(
        prince_inst_sbox_inst7_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst7_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst7_yxyy_inst_U15 ( .A(
        prince_inst_sbox_inst7_yxyy_inst_n67), .B(
        prince_inst_sbox_inst7_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst7_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U14 ( .A1(prince_inst_sin_y[31]), 
        .A2(prince_inst_sin_y[28]), .ZN(prince_inst_sbox_inst7_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst7_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst7_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst7_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst7_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst7_yxyy_inst_U12 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst7_yxyy_inst_U11 ( .A(
        prince_inst_sbox_inst7_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst7_yxyy_inst_U10 ( .A1(prince_inst_sin_x[29]), 
        .A2(prince_inst_sin_y[30]), .A3(prince_inst_sin_y[28]), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U9 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst7_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U8 ( .A1(prince_inst_sin_y[31]), 
        .A2(prince_inst_sbox_inst7_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst7_yxyy_inst_U7 ( .A1(prince_inst_sin_y[30]), 
        .A2(prince_inst_sin_x[29]), .ZN(prince_inst_sbox_inst7_yxyy_inst_n49)
         );
  OR3_X1 prince_inst_sbox_inst7_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst7_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst7_yxyy_inst_U5 ( .A(prince_inst_sin_y[28]), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst7_yxyy_inst_U4 ( .A(prince_inst_sin_x[29]), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst7_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst7_yxyy_inst_n64), .A2(
        prince_inst_sbox_inst7_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst7_yxyy_inst_U2 ( .A(prince_inst_sin_y[31]), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst7_yxyy_inst_U1 ( .A(prince_inst_sin_y[30]), .ZN(
        prince_inst_sbox_inst7_yxyy_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst7_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U29 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst7_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst7_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst7_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n75), .A2(prince_inst_sin_y[31]), 
        .A3(prince_inst_sbox_inst7_yyxy_inst_n70), .A4(prince_inst_sin_x[30]), 
        .ZN(prince_inst_sbox_inst7_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst7_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n69), .A3(prince_inst_sin_y[29]), 
        .A4(prince_inst_sbox_inst7_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst7_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst7_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst7_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst7_yyxy_inst_U23 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_x[30]), .A3(prince_inst_sin_y[28]), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst7_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n69), .A2(prince_inst_sin_y[29]), 
        .A3(prince_inst_sin_y[31]), .ZN(prince_inst_sbox_inst7_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst7_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n75), .A2(prince_inst_sin_x[30]), 
        .A3(prince_inst_sin_y[31]), .ZN(prince_inst_sbox_inst7_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst7_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst7_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst7_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n61), .A2(prince_inst_sin_x[30]), 
        .ZN(prince_inst_sbox_inst7_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst7_yyxy_inst_U18 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_y[31]), .A3(prince_inst_sbox_inst7_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst7_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst7_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst7_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst7_yyxy_inst_U16 ( .A1(prince_inst_sin_y[31]), 
        .A2(prince_inst_sbox_inst7_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst7_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst7_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst7_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n58), .A3(prince_inst_sin_y[28]), 
        .ZN(prince_inst_sbox_inst7_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst7_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst7_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst7_yyxy_inst_U13 ( .A1(prince_inst_sin_y[28]), 
        .A2(prince_inst_sbox_inst7_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst7_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst7_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst7_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst7_yyxy_inst_n54), .B(
        prince_inst_sbox_inst7_yyxy_inst_n55), .S(
        prince_inst_sbox_inst7_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst7_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst7_yyxy_inst_U9 ( .A(prince_inst_sin_x[30]), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n75), .A2(prince_inst_sin_y[31]), 
        .ZN(prince_inst_sbox_inst7_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst7_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst7_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst7_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U5 ( .A1(prince_inst_sin_x[30]), 
        .A2(prince_inst_sbox_inst7_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst7_yyxy_inst_U4 ( .A(prince_inst_sin_y[29]), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst7_yyxy_inst_U3 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sbox_inst7_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst7_yyxy_inst_U2 ( .A(prince_inst_sin_y[28]), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst7_yyxy_inst_U1 ( .A(prince_inst_sin_y[31]), .ZN(
        prince_inst_sbox_inst7_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst7_yyyx_inst_n58), .B(
        prince_inst_sbox_inst7_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst7_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst7_yyyx_inst_n56), .B(
        prince_inst_sbox_inst7_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst7_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst7_yyyx_inst_n54), .B(
        prince_inst_sbox_inst7_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst7_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst7_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst7_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst7_yyyx_inst_U21 ( .A1(prince_inst_sin_x[31]), 
        .A2(prince_inst_sbox_inst7_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst7_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst7_yyyx_inst_U20 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_y[30]), .A3(prince_inst_sbox_inst7_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst7_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst7_yyyx_inst_n50), .B(
        prince_inst_sbox_inst7_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst7_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst7_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n56), .A2(prince_inst_sin_y[30]), 
        .ZN(prince_inst_sbox_inst7_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst7_yyyx_inst_U17 ( .A1(prince_inst_sin_y[29]), 
        .A2(prince_inst_sin_y[28]), .A3(prince_inst_sin_y[30]), .ZN(
        prince_inst_sbox_inst7_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst7_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst7_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst7_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst7_yyyx_inst_U15 ( .A1(prince_inst_sin_x[31]), 
        .A2(prince_inst_sin_y[30]), .A3(prince_inst_sbox_inst7_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst7_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst7_yyyx_inst_U14 ( .A(prince_inst_sin_y[28]), 
        .ZN(prince_inst_sbox_inst7_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n58), .A2(prince_inst_sin_y[29]), 
        .ZN(prince_inst_sbox_inst7_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst7_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst7_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U11 ( .A1(prince_inst_sin_y[28]), 
        .A2(prince_inst_sbox_inst7_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst7_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst7_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst7_yyyx_inst_U9 ( .A1(prince_inst_sin_y[28]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst7_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst7_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst7_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst7_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n45), .A2(prince_inst_sin_y[28]), 
        .A3(prince_inst_sin_y[30]), .ZN(prince_inst_sbox_inst7_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst7_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst7_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst7_yyyx_inst_U4 ( .A1(prince_inst_sin_x[31]), 
        .A2(prince_inst_sin_y[30]), .ZN(prince_inst_sbox_inst7_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst7_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst7_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst7_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst7_yyyx_inst_U2 ( .A(prince_inst_sin_y[29]), .ZN(
        prince_inst_sbox_inst7_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst7_yyyx_inst_U1 ( .A1(prince_inst_sin_y[28]), 
        .A2(prince_inst_sin_x[31]), .ZN(prince_inst_sbox_inst7_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s00_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[0]), .B(prince_inst_sbox_inst7_s0_sh[0]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s01_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[1]), .B(prince_inst_sbox_inst7_s0_sh[1]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s02_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[2]), .B(prince_inst_sbox_inst7_s0_sh[2]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s03_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[3]), .B(prince_inst_sbox_inst7_s0_sh[3]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s04_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[4]), .B(prince_inst_sbox_inst7_s0_sh[4]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s05_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[5]), .B(prince_inst_sbox_inst7_s0_sh[5]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s06_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[6]), .B(prince_inst_sbox_inst7_s0_sh[6]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s07_U1 ( .A(
        prince_inst_sbox_inst7_t0_sh[7]), .B(prince_inst_sbox_inst7_s0_sh[7]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s10_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[0]), .B(prince_inst_sbox_inst7_s1_sh[0]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s11_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[1]), .B(prince_inst_sbox_inst7_s1_sh[1]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s12_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[2]), .B(prince_inst_sbox_inst7_s1_sh[2]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s13_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[3]), .B(prince_inst_sbox_inst7_s1_sh[3]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s14_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[4]), .B(prince_inst_sbox_inst7_s1_sh[4]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s15_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[5]), .B(prince_inst_sbox_inst7_s1_sh[5]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s16_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[6]), .B(prince_inst_sbox_inst7_s1_sh[6]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s17_U1 ( .A(
        prince_inst_sbox_inst7_t1_sh[7]), .B(prince_inst_sbox_inst7_s1_sh[7]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s20_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[0]), .B(prince_inst_sbox_inst7_s2_sh[0]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s21_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[1]), .B(prince_inst_sbox_inst7_s2_sh[1]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s22_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[2]), .B(prince_inst_sbox_inst7_s2_sh[2]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s23_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[3]), .B(prince_inst_sbox_inst7_s2_sh[3]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s24_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[4]), .B(prince_inst_sbox_inst7_s2_sh[4]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s25_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[5]), .B(prince_inst_sbox_inst7_s2_sh[5]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s26_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[6]), .B(prince_inst_sbox_inst7_s2_sh[6]), 
        .S(prince_inst_sbox_inst7_n8), .Z(prince_inst_sbox_inst7_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s27_U1 ( .A(
        prince_inst_sbox_inst7_t2_sh[7]), .B(prince_inst_sbox_inst7_s2_sh[7]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s30_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[0]), .B(prince_inst_sbox_inst7_s3_sh[0]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s31_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[1]), .B(prince_inst_sbox_inst7_s3_sh[1]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s32_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[2]), .B(prince_inst_sbox_inst7_s3_sh[2]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s33_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[3]), .B(prince_inst_sbox_inst7_s3_sh[3]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s34_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[4]), .B(prince_inst_sbox_inst7_s3_sh[4]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s35_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[5]), .B(prince_inst_sbox_inst7_s3_sh[5]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s36_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[6]), .B(prince_inst_sbox_inst7_s3_sh[6]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst7_mux_s37_U1 ( .A(
        prince_inst_sbox_inst7_t3_sh[7]), .B(prince_inst_sbox_inst7_s3_sh[7]), 
        .S(prince_inst_sbox_inst7_n9), .Z(prince_inst_sbox_inst7_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk0_U1 ( .A(r[48]), .B(
        prince_inst_sbox_inst7_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk1_U1 ( .A(r[49]), .B(
        prince_inst_sbox_inst7_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[1]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk2_U1 ( .A(r[50]), .B(
        prince_inst_sbox_inst7_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[2]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk3_U1 ( .A(r[51]), .B(
        prince_inst_sbox_inst7_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[3]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk4_U1 ( .A(r[48]), .B(
        prince_inst_sbox_inst7_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk5_U1 ( .A(r[49]), .B(
        prince_inst_sbox_inst7_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[5]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk6_U1 ( .A(r[50]), .B(
        prince_inst_sbox_inst7_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[6]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_msk7_U1 ( .A(r[51]), .B(
        prince_inst_sbox_inst7_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst7_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst0_y[7]), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst7_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst7_c_inst0_ax_n5), .ZN(prince_inst_sout_x[28]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst7_c_inst0_y[1]), .B(
        prince_inst_sbox_inst7_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst7_c_inst0_y[2]), .B(
        prince_inst_sbox_inst7_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst7_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst7_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst7_c_inst0_ay_n5), .ZN(final_y[28]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst7_c_inst0_y[5]), .B(
        prince_inst_sbox_inst7_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst7_c_inst0_y[6]), .B(
        prince_inst_sbox_inst7_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst7_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk0_U1 ( .A(r[52]), .B(
        prince_inst_sbox_inst7_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk1_U1 ( .A(r[53]), .B(
        prince_inst_sbox_inst7_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[1]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk2_U1 ( .A(r[54]), .B(
        prince_inst_sbox_inst7_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[2]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk3_U1 ( .A(r[55]), .B(
        prince_inst_sbox_inst7_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[3]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk4_U1 ( .A(r[52]), .B(
        prince_inst_sbox_inst7_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk5_U1 ( .A(r[53]), .B(
        prince_inst_sbox_inst7_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[5]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk6_U1 ( .A(r[54]), .B(
        prince_inst_sbox_inst7_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[6]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_msk7_U1 ( .A(r[55]), .B(
        prince_inst_sbox_inst7_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst7_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst1_y[7]), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst7_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst7_c_inst1_ax_n5), .ZN(prince_inst_sout_x[29]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst7_c_inst1_y[1]), .B(
        prince_inst_sbox_inst7_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst7_c_inst1_y[2]), .B(
        prince_inst_sbox_inst7_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst7_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst7_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst7_c_inst1_ay_n5), .ZN(final_y[29]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst7_c_inst1_y[5]), .B(
        prince_inst_sbox_inst7_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst7_c_inst1_y[6]), .B(
        prince_inst_sbox_inst7_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst7_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk0_U1 ( .A(r[56]), .B(
        prince_inst_sbox_inst7_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk1_U1 ( .A(r[57]), .B(
        prince_inst_sbox_inst7_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[1]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk2_U1 ( .A(r[58]), .B(
        prince_inst_sbox_inst7_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[2]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk3_U1 ( .A(r[59]), .B(
        prince_inst_sbox_inst7_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[3]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk4_U1 ( .A(r[56]), .B(
        prince_inst_sbox_inst7_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk5_U1 ( .A(r[57]), .B(
        prince_inst_sbox_inst7_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[5]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk6_U1 ( .A(r[58]), .B(
        prince_inst_sbox_inst7_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[6]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_msk7_U1 ( .A(r[59]), .B(
        prince_inst_sbox_inst7_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst7_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst2_y[7]), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst7_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst7_c_inst2_ax_n5), .ZN(prince_inst_sout_x[30]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst7_c_inst2_y[1]), .B(
        prince_inst_sbox_inst7_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst7_c_inst2_y[2]), .B(
        prince_inst_sbox_inst7_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst7_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst7_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst7_c_inst2_ay_n5), .ZN(final_y[30]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst7_c_inst2_y[5]), .B(
        prince_inst_sbox_inst7_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst7_c_inst2_y[6]), .B(
        prince_inst_sbox_inst7_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst7_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk0_U1 ( .A(r[60]), .B(
        prince_inst_sbox_inst7_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk1_U1 ( .A(r[61]), .B(
        prince_inst_sbox_inst7_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[1]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk2_U1 ( .A(r[62]), .B(
        prince_inst_sbox_inst7_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[2]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk3_U1 ( .A(r[63]), .B(
        prince_inst_sbox_inst7_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[3]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk4_U1 ( .A(r[60]), .B(
        prince_inst_sbox_inst7_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk5_U1 ( .A(r[61]), .B(
        prince_inst_sbox_inst7_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[5]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk6_U1 ( .A(r[62]), .B(
        prince_inst_sbox_inst7_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[6]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_msk7_U1 ( .A(r[63]), .B(
        prince_inst_sbox_inst7_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst7_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst7_n6), .A3(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_U5 ( .A1(en_sig), .A2(
        prince_inst_sbox_inst7_c_inst3_y[7]), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst7_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst7_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst7_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst7_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst7_c_inst3_ax_n5), .ZN(prince_inst_sout_x[31]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst7_c_inst3_y[1]), .B(
        prince_inst_sbox_inst7_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst7_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst7_c_inst3_y[2]), .B(
        prince_inst_sbox_inst7_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst7_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst7_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst7_c_inst3_ay_n5), .ZN(final_y[31]) );
  XNOR2_X1 prince_inst_sbox_inst7_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst7_c_inst3_y[5]), .B(
        prince_inst_sbox_inst7_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst7_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst7_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst7_c_inst3_y[6]), .B(
        prince_inst_sbox_inst7_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst7_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst8_U5 ( .A(prince_inst_sbox_inst8_n10), .ZN(
        prince_inst_sbox_inst8_n9) );
  INV_X1 prince_inst_sbox_inst8_U4 ( .A(prince_inst_n27), .ZN(
        prince_inst_sbox_inst8_n8) );
  INV_X1 prince_inst_sbox_inst8_U3 ( .A(prince_inst_sbox_inst8_n8), .ZN(
        prince_inst_sbox_inst8_n6) );
  INV_X1 prince_inst_sbox_inst8_U2 ( .A(prince_inst_sbox_inst8_n8), .ZN(
        prince_inst_sbox_inst8_n7) );
  INV_X1 prince_inst_sbox_inst8_U1 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst8_n10) );
  NAND3_X1 prince_inst_sbox_inst8_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n68), .A3(prince_inst_sin_x[32]), 
        .ZN(prince_inst_sbox_inst8_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U25 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sbox_inst8_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst8_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst8_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst8_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst8_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n67), .A2(prince_inst_sin_x[34]), 
        .A3(prince_inst_sin_x[32]), .A4(prince_inst_sin_y[35]), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst8_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n61), .A2(prince_inst_sin_x[33]), 
        .A3(prince_inst_sin_x[34]), .ZN(prince_inst_sbox_inst8_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst8_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n66), .A3(prince_inst_sin_x[33]), 
        .A4(prince_inst_sin_x[32]), .ZN(prince_inst_sbox_inst8_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst8_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst8_xxxy_inst_n59), .B(prince_inst_sin_y[35]), .Z(
        prince_inst_sbox_inst8_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U18 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sin_x[33]), .ZN(prince_inst_sbox_inst8_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst8_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst8_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n65), .A2(prince_inst_sin_x[34]), 
        .ZN(prince_inst_sbox_inst8_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst8_xxxy_inst_U15 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sin_y[35]), .A3(prince_inst_sbox_inst8_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst8_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst8_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst8_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst8_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst8_xxxy_inst_U13 ( .A(prince_inst_sin_x[32]), 
        .B(prince_inst_sin_x[33]), .S(prince_inst_sbox_inst8_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst8_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst8_xxxy_inst_U12 ( .A(prince_inst_sin_y[35]), 
        .ZN(prince_inst_sbox_inst8_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U11 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sin_x[32]), .ZN(prince_inst_sbox_inst8_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst8_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst8_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst8_xxxy_inst_n60), .B(
        prince_inst_sbox_inst8_xxxy_inst_n53), .S(
        prince_inst_sbox_inst8_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst8_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U8 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sbox_inst8_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U7 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sin_y[35]), .ZN(prince_inst_sbox_inst8_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst8_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst8_t1_sh[0]), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst8_xxxy_inst_U5 ( .A(prince_inst_sin_x[34]), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U4 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sbox_inst8_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst8_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst8_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst8_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst8_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst8_xxxy_inst_U2 ( .A(prince_inst_sin_x[32]), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst8_xxxy_inst_U1 ( .A(prince_inst_sin_x[33]), .ZN(
        prince_inst_sbox_inst8_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst8_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst8_t1_sh[1]), .B(
        prince_inst_sbox_inst8_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst8_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst8_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst8_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst8_xxyx_inst_n52), .B(
        prince_inst_sbox_inst8_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst8_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U23 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst8_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst8_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n48), .A2(prince_inst_sin_x[35]), 
        .A3(prince_inst_sin_x[32]), .ZN(prince_inst_sbox_inst8_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n45), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst8_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst8_xxyx_inst_U18 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n46), .A2(prince_inst_sin_x[35]), 
        .A3(prince_inst_sin_x[33]), .ZN(prince_inst_sbox_inst8_xxyx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst8_t2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst8_xxyx_inst_U16 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sin_x[32]), .A3(prince_inst_sbox_inst8_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst8_xxyx_inst_n44) );
  OR2_X1 prince_inst_sbox_inst8_xxyx_inst_U15 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sbox_inst8_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst8_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst8_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst8_xxyx_inst_n54), .B(
        prince_inst_sbox_inst8_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst8_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U12 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sin_y[34]), .ZN(prince_inst_sbox_inst8_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst8_xxyx_inst_U11 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sbox_inst8_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst8_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst8_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst8_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst8_xxyx_inst_U10 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst8_xxyx_inst_U9 ( .A1(prince_inst_sin_x[35]), 
        .A2(prince_inst_sbox_inst8_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst8_xxyx_inst_U8 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sbox_inst8_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst8_xxyx_inst_U7 ( .A(prince_inst_sin_y[34]), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst8_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst8_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst8_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n53), .A2(prince_inst_sin_x[33]), 
        .A3(prince_inst_sin_y[34]), .A4(prince_inst_sin_x[32]), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst8_xxyx_inst_U4 ( .A(prince_inst_sin_x[35]), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst8_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst8_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst8_xxyx_inst_n43), .A3(prince_inst_sin_x[35]), 
        .A4(prince_inst_sin_y[34]), .ZN(prince_inst_sbox_inst8_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst8_xxyx_inst_U2 ( .A(prince_inst_sin_x[32]), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst8_xxyx_inst_U1 ( .A(prince_inst_sin_x[33]), .ZN(
        prince_inst_sbox_inst8_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst8_xyxx_inst_n74), .B(
        prince_inst_sbox_inst8_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst8_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst8_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst8_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst8_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U26 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sbox_inst8_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U25 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst8_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst8_xyxx_inst_n72), .B(
        prince_inst_sbox_inst8_s0_sh[2]), .S(
        prince_inst_sbox_inst8_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst8_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst8_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n74), .A2(prince_inst_sin_x[35]), 
        .ZN(prince_inst_sbox_inst8_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst8_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U21 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sbox_inst8_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst8_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst8_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst8_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst8_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst8_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst8_xyxx_inst_U15 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_x[32]), .ZN(prince_inst_sbox_inst8_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst8_xyxx_inst_U13 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U12 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_x[34]), .ZN(prince_inst_sbox_inst8_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst8_xyxx_inst_n58), .B(
        prince_inst_sbox_inst8_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst8_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst8_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst8_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst8_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst8_xyxx_inst_U9 ( .A(prince_inst_sin_x[35]), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst8_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n54), .A2(prince_inst_sin_x[32]), 
        .ZN(prince_inst_sbox_inst8_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst8_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst8_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst8_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst8_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst8_xyxx_inst_U5 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sbox_inst8_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst8_xyxx_inst_U4 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst8_xyxx_inst_U3 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sbox_inst8_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst8_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst8_xyxx_inst_U2 ( .A(prince_inst_sin_y[33]), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst8_xyxx_inst_U1 ( .A(prince_inst_sin_x[34]), .ZN(
        prince_inst_sbox_inst8_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst8_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst8_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst8_xyyy_inst_n59), .B(
        prince_inst_sbox_inst8_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst8_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst8_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst8_xyyy_inst_U25 ( .A1(prince_inst_sin_y[34]), 
        .A2(prince_inst_sin_y[35]), .A3(prince_inst_sbox_inst8_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst8_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U24 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sbox_inst8_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U23 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sbox_inst8_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst8_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst8_xyyy_inst_U19 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sin_y[34]), .A3(prince_inst_sbox_inst8_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst8_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst8_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst8_xyyy_inst_n49), .B(
        prince_inst_sbox_inst8_xyyy_inst_n48), .S(
        prince_inst_sbox_inst8_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst8_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst8_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst8_xyyy_inst_U16 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sbox_inst8_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst8_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst8_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst8_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst8_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst8_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst8_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst8_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst8_xyyy_inst_U12 ( .A(prince_inst_sin_y[35]), 
        .ZN(prince_inst_sbox_inst8_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst8_xyyy_inst_U11 ( .A1(prince_inst_sin_y[35]), 
        .A2(prince_inst_sbox_inst8_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst8_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst8_t1_sh[3]), .B(
        prince_inst_sbox_inst8_xyyy_inst_n48), .S(
        prince_inst_sbox_inst8_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst8_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst8_xyyy_inst_U9 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sbox_inst8_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst8_xyyy_inst_U8 ( .A1(prince_inst_sin_x[32]), 
        .A2(prince_inst_sin_y[35]), .ZN(prince_inst_sbox_inst8_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst8_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst8_t1_sh[3]), .ZN(prince_inst_sbox_inst8_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst8_xyyy_inst_U6 ( .A1(prince_inst_sin_y[35]), 
        .A2(prince_inst_sbox_inst8_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst8_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst8_xyyy_inst_U4 ( .A(prince_inst_sin_y[33]), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst8_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst8_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst8_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst8_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst8_xyyy_inst_U2 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_x[32]), .ZN(prince_inst_sbox_inst8_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst8_xyyy_inst_U1 ( .A(prince_inst_sin_y[34]), .ZN(
        prince_inst_sbox_inst8_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst8_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U27 ( .A1(prince_inst_sin_y[32]), 
        .A2(prince_inst_sbox_inst8_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst8_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U24 ( .A1(prince_inst_sin_y[32]), 
        .A2(prince_inst_sbox_inst8_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst8_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U21 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst8_yxxx_inst_U19 ( .A(prince_inst_sin_x[35]), 
        .ZN(prince_inst_sbox_inst8_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst8_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst8_yxxx_inst_n52), .B(
        prince_inst_sbox_inst8_yxxx_inst_n51), .S(
        prince_inst_sbox_inst8_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst8_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n53), .A2(prince_inst_sin_x[35]), 
        .ZN(prince_inst_sbox_inst8_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst8_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n48), .A2(prince_inst_sin_y[32]), 
        .ZN(prince_inst_sbox_inst8_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n47), .A2(prince_inst_sin_x[35]), 
        .ZN(prince_inst_sbox_inst8_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U13 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sbox_inst8_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst8_yxxx_inst_n59), .B(
        prince_inst_sbox_inst8_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst8_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst8_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst8_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst8_yxxx_inst_U9 ( .A1(prince_inst_sin_x[33]), 
        .A2(prince_inst_sbox_inst8_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst8_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst8_yxxx_inst_U8 ( .A(prince_inst_sin_x[34]), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst8_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst8_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst8_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst8_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst8_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst8_yxxx_inst_U5 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sbox_inst8_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst8_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst8_yxxx_inst_U4 ( .A(prince_inst_sin_y[32]), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst8_yxxx_inst_U3 ( .A(prince_inst_sin_x[33]), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst8_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst8_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst8_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst8_yxxx_inst_U1 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst8_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst8_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst8_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst8_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst8_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n64), .A3(prince_inst_sin_y[35]), 
        .ZN(prince_inst_sbox_inst8_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst8_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n63), .A2(prince_inst_sin_y[34]), 
        .A3(prince_inst_sin_y[35]), .ZN(prince_inst_sbox_inst8_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst8_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst8_yxyy_inst_n62), .B(
        prince_inst_sbox_inst8_yxyy_inst_n61), .S(prince_inst_sin_y[32]), .Z(
        prince_inst_sbox_inst8_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst8_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst8_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst8_yxyy_inst_n64), .B(
        prince_inst_sbox_inst8_yxyy_inst_n60), .S(
        prince_inst_sbox_inst8_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst8_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst8_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst8_yxyy_inst_n62), .B(
        prince_inst_sbox_inst8_yxyy_inst_n54), .S(
        prince_inst_sbox_inst8_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst8_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst8_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst8_yxyy_inst_n53), .B(
        prince_inst_sbox_inst8_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst8_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst8_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst8_yxyy_inst_n68), .B(
        prince_inst_sbox_inst8_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst8_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U15 ( .A1(prince_inst_sin_y[35]), 
        .A2(prince_inst_sin_y[32]), .ZN(prince_inst_sbox_inst8_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst8_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst8_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst8_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst8_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst8_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst8_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst8_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst8_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n64), .A2(prince_inst_sin_y[34]), 
        .A3(prince_inst_sin_y[32]), .ZN(prince_inst_sbox_inst8_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst8_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U9 ( .A1(prince_inst_sin_y[35]), 
        .A2(prince_inst_sbox_inst8_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst8_yxyy_inst_U8 ( .A1(prince_inst_sin_y[34]), 
        .A2(prince_inst_sbox_inst8_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst8_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst8_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst8_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst8_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst8_yxyy_inst_U5 ( .A(prince_inst_sin_y[32]), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst8_yxyy_inst_U4 ( .A(prince_inst_sin_x[33]), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst8_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst8_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst8_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst8_yxyy_inst_U2 ( .A(prince_inst_sin_y[35]), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst8_yxyy_inst_U1 ( .A(prince_inst_sin_y[34]), .ZN(
        prince_inst_sbox_inst8_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst8_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U29 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sbox_inst8_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst8_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst8_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst8_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n75), .A2(prince_inst_sin_y[35]), 
        .A3(prince_inst_sbox_inst8_yyxy_inst_n70), .A4(prince_inst_sin_x[34]), 
        .ZN(prince_inst_sbox_inst8_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst8_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n69), .A3(prince_inst_sin_y[33]), 
        .A4(prince_inst_sbox_inst8_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst8_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst8_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst8_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst8_yyxy_inst_U23 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_x[34]), .A3(prince_inst_sin_y[32]), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst8_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n69), .A2(prince_inst_sin_y[33]), 
        .A3(prince_inst_sin_y[35]), .ZN(prince_inst_sbox_inst8_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst8_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n75), .A2(prince_inst_sin_x[34]), 
        .A3(prince_inst_sin_y[35]), .ZN(prince_inst_sbox_inst8_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst8_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst8_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst8_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n61), .A2(prince_inst_sin_x[34]), 
        .ZN(prince_inst_sbox_inst8_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst8_yyxy_inst_U18 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_y[35]), .A3(prince_inst_sbox_inst8_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst8_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst8_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst8_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst8_yyxy_inst_U16 ( .A1(prince_inst_sin_y[35]), 
        .A2(prince_inst_sbox_inst8_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst8_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst8_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst8_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n58), .A3(prince_inst_sin_y[32]), 
        .ZN(prince_inst_sbox_inst8_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst8_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst8_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst8_yyxy_inst_U13 ( .A1(prince_inst_sin_y[32]), 
        .A2(prince_inst_sbox_inst8_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst8_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst8_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst8_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst8_yyxy_inst_n54), .B(
        prince_inst_sbox_inst8_yyxy_inst_n55), .S(
        prince_inst_sbox_inst8_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst8_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst8_yyxy_inst_U9 ( .A(prince_inst_sin_x[34]), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n75), .A2(prince_inst_sin_y[35]), 
        .ZN(prince_inst_sbox_inst8_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst8_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst8_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst8_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U5 ( .A1(prince_inst_sin_x[34]), 
        .A2(prince_inst_sbox_inst8_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst8_yyxy_inst_U4 ( .A(prince_inst_sin_y[33]), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst8_yyxy_inst_U3 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sbox_inst8_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst8_yyxy_inst_U2 ( .A(prince_inst_sin_y[32]), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst8_yyxy_inst_U1 ( .A(prince_inst_sin_y[35]), .ZN(
        prince_inst_sbox_inst8_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst8_yyyx_inst_n58), .B(
        prince_inst_sbox_inst8_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst8_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst8_yyyx_inst_n56), .B(
        prince_inst_sbox_inst8_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst8_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst8_yyyx_inst_n54), .B(
        prince_inst_sbox_inst8_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst8_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst8_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst8_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst8_yyyx_inst_U21 ( .A1(prince_inst_sin_x[35]), 
        .A2(prince_inst_sbox_inst8_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst8_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst8_yyyx_inst_U20 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_y[34]), .A3(prince_inst_sbox_inst8_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst8_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst8_yyyx_inst_n50), .B(
        prince_inst_sbox_inst8_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst8_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst8_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n56), .A2(prince_inst_sin_y[34]), 
        .ZN(prince_inst_sbox_inst8_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst8_yyyx_inst_U17 ( .A1(prince_inst_sin_y[33]), 
        .A2(prince_inst_sin_y[32]), .A3(prince_inst_sin_y[34]), .ZN(
        prince_inst_sbox_inst8_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst8_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst8_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst8_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst8_yyyx_inst_U15 ( .A1(prince_inst_sin_x[35]), 
        .A2(prince_inst_sin_y[34]), .A3(prince_inst_sbox_inst8_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst8_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst8_yyyx_inst_U14 ( .A(prince_inst_sin_y[32]), 
        .ZN(prince_inst_sbox_inst8_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n58), .A2(prince_inst_sin_y[33]), 
        .ZN(prince_inst_sbox_inst8_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst8_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst8_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U11 ( .A1(prince_inst_sin_y[32]), 
        .A2(prince_inst_sbox_inst8_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst8_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst8_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst8_yyyx_inst_U9 ( .A1(prince_inst_sin_y[32]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst8_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst8_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst8_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst8_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n45), .A2(prince_inst_sin_y[32]), 
        .A3(prince_inst_sin_y[34]), .ZN(prince_inst_sbox_inst8_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst8_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst8_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst8_yyyx_inst_U4 ( .A1(prince_inst_sin_x[35]), 
        .A2(prince_inst_sin_y[34]), .ZN(prince_inst_sbox_inst8_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst8_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst8_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst8_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst8_yyyx_inst_U2 ( .A(prince_inst_sin_y[33]), .ZN(
        prince_inst_sbox_inst8_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst8_yyyx_inst_U1 ( .A1(prince_inst_sin_y[32]), 
        .A2(prince_inst_sin_x[35]), .ZN(prince_inst_sbox_inst8_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s00_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[0]), .B(prince_inst_sbox_inst8_s0_sh[0]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s01_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[1]), .B(prince_inst_sbox_inst8_s0_sh[1]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s02_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[2]), .B(prince_inst_sbox_inst8_s0_sh[2]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s03_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[3]), .B(prince_inst_sbox_inst8_s0_sh[3]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s04_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[4]), .B(prince_inst_sbox_inst8_s0_sh[4]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s05_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[5]), .B(prince_inst_sbox_inst8_s0_sh[5]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s06_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[6]), .B(prince_inst_sbox_inst8_s0_sh[6]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s07_U1 ( .A(
        prince_inst_sbox_inst8_t0_sh[7]), .B(prince_inst_sbox_inst8_s0_sh[7]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s10_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[0]), .B(prince_inst_sbox_inst8_s1_sh[0]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s11_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[1]), .B(prince_inst_sbox_inst8_s1_sh[1]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s12_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[2]), .B(prince_inst_sbox_inst8_s1_sh[2]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s13_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[3]), .B(prince_inst_sbox_inst8_s1_sh[3]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s14_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[4]), .B(prince_inst_sbox_inst8_s1_sh[4]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s15_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[5]), .B(prince_inst_sbox_inst8_s1_sh[5]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s16_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[6]), .B(prince_inst_sbox_inst8_s1_sh[6]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s17_U1 ( .A(
        prince_inst_sbox_inst8_t1_sh[7]), .B(prince_inst_sbox_inst8_s1_sh[7]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s20_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[0]), .B(prince_inst_sbox_inst8_s2_sh[0]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s21_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[1]), .B(prince_inst_sbox_inst8_s2_sh[1]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s22_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[2]), .B(prince_inst_sbox_inst8_s2_sh[2]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s23_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[3]), .B(prince_inst_sbox_inst8_s2_sh[3]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s24_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[4]), .B(prince_inst_sbox_inst8_s2_sh[4]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s25_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[5]), .B(prince_inst_sbox_inst8_s2_sh[5]), 
        .S(prince_inst_sbox_inst8_n6), .Z(prince_inst_sbox_inst8_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s26_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[6]), .B(prince_inst_sbox_inst8_s2_sh[6]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s27_U1 ( .A(
        prince_inst_sbox_inst8_t2_sh[7]), .B(prince_inst_sbox_inst8_s2_sh[7]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s30_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[0]), .B(prince_inst_sbox_inst8_s3_sh[0]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s31_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[1]), .B(prince_inst_sbox_inst8_s3_sh[1]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s32_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[2]), .B(prince_inst_sbox_inst8_s3_sh[2]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s33_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[3]), .B(prince_inst_sbox_inst8_s3_sh[3]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s34_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[4]), .B(prince_inst_sbox_inst8_s3_sh[4]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s35_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[5]), .B(prince_inst_sbox_inst8_s3_sh[5]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s36_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[6]), .B(prince_inst_sbox_inst8_s3_sh[6]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst8_mux_s37_U1 ( .A(
        prince_inst_sbox_inst8_t3_sh[7]), .B(prince_inst_sbox_inst8_s3_sh[7]), 
        .S(prince_inst_sbox_inst8_n7), .Z(prince_inst_sbox_inst8_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk0_U1 ( .A(r[64]), .B(
        prince_inst_sbox_inst8_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk1_U1 ( .A(r[65]), .B(
        prince_inst_sbox_inst8_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk2_U1 ( .A(r[66]), .B(
        prince_inst_sbox_inst8_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk3_U1 ( .A(r[67]), .B(
        prince_inst_sbox_inst8_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk4_U1 ( .A(r[64]), .B(
        prince_inst_sbox_inst8_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk5_U1 ( .A(r[65]), .B(
        prince_inst_sbox_inst8_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk6_U1 ( .A(r[66]), .B(
        prince_inst_sbox_inst8_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_msk7_U1 ( .A(r[67]), .B(
        prince_inst_sbox_inst8_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst8_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst8_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst8_c_inst0_ax_n5), .ZN(prince_inst_sout_x[32]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst8_c_inst0_y[1]), .B(
        prince_inst_sbox_inst8_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst8_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst8_c_inst0_y[2]), .B(
        prince_inst_sbox_inst8_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst8_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst8_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst8_c_inst0_ay_n5), .ZN(final_y[16]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst8_c_inst0_y[5]), .B(
        prince_inst_sbox_inst8_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst8_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst8_c_inst0_y[6]), .B(
        prince_inst_sbox_inst8_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst8_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk0_U1 ( .A(r[68]), .B(
        prince_inst_sbox_inst8_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk1_U1 ( .A(r[69]), .B(
        prince_inst_sbox_inst8_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk2_U1 ( .A(r[70]), .B(
        prince_inst_sbox_inst8_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk3_U1 ( .A(r[71]), .B(
        prince_inst_sbox_inst8_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk4_U1 ( .A(r[68]), .B(
        prince_inst_sbox_inst8_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk5_U1 ( .A(r[69]), .B(
        prince_inst_sbox_inst8_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk6_U1 ( .A(r[70]), .B(
        prince_inst_sbox_inst8_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_msk7_U1 ( .A(r[71]), .B(
        prince_inst_sbox_inst8_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst8_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst8_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst8_c_inst1_ax_n5), .ZN(prince_inst_sout_x[33]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst8_c_inst1_y[1]), .B(
        prince_inst_sbox_inst8_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst8_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst8_c_inst1_y[2]), .B(
        prince_inst_sbox_inst8_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst8_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst8_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst8_c_inst1_ay_n5), .ZN(final_y[17]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst8_c_inst1_y[5]), .B(
        prince_inst_sbox_inst8_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst8_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst8_c_inst1_y[6]), .B(
        prince_inst_sbox_inst8_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst8_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk0_U1 ( .A(r[72]), .B(
        prince_inst_sbox_inst8_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk1_U1 ( .A(r[73]), .B(
        prince_inst_sbox_inst8_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk2_U1 ( .A(r[74]), .B(
        prince_inst_sbox_inst8_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk3_U1 ( .A(r[75]), .B(
        prince_inst_sbox_inst8_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk4_U1 ( .A(r[72]), .B(
        prince_inst_sbox_inst8_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk5_U1 ( .A(r[73]), .B(
        prince_inst_sbox_inst8_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk6_U1 ( .A(r[74]), .B(
        prince_inst_sbox_inst8_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_msk7_U1 ( .A(r[75]), .B(
        prince_inst_sbox_inst8_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst8_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst8_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst8_c_inst2_ax_n5), .ZN(prince_inst_sout_x[34]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst8_c_inst2_y[1]), .B(
        prince_inst_sbox_inst8_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst8_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst8_c_inst2_y[2]), .B(
        prince_inst_sbox_inst8_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst8_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst8_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst8_c_inst2_ay_n5), .ZN(final_y[18]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst8_c_inst2_y[5]), .B(
        prince_inst_sbox_inst8_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst8_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst8_c_inst2_y[6]), .B(
        prince_inst_sbox_inst8_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst8_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk0_U1 ( .A(r[76]), .B(
        prince_inst_sbox_inst8_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk1_U1 ( .A(r[77]), .B(
        prince_inst_sbox_inst8_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk2_U1 ( .A(r[78]), .B(
        prince_inst_sbox_inst8_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk3_U1 ( .A(r[79]), .B(
        prince_inst_sbox_inst8_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk4_U1 ( .A(r[76]), .B(
        prince_inst_sbox_inst8_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk5_U1 ( .A(r[77]), .B(
        prince_inst_sbox_inst8_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk6_U1 ( .A(r[78]), .B(
        prince_inst_sbox_inst8_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_msk7_U1 ( .A(r[79]), .B(
        prince_inst_sbox_inst8_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst8_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst8_n9), .A2(prince_inst_sbox_inst8_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst8_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst8_n9), .ZN(
        prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst8_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst8_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst8_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst8_c_inst3_ax_n5), .ZN(prince_inst_sout_x[35]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst8_c_inst3_y[1]), .B(
        prince_inst_sbox_inst8_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst8_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst8_c_inst3_y[2]), .B(
        prince_inst_sbox_inst8_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst8_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst8_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst8_c_inst3_ay_n5), .ZN(final_y[19]) );
  XNOR2_X1 prince_inst_sbox_inst8_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst8_c_inst3_y[5]), .B(
        prince_inst_sbox_inst8_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst8_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst8_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst8_c_inst3_y[6]), .B(
        prince_inst_sbox_inst8_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst8_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst9_U5 ( .A(prince_inst_sbox_inst9_n10), .ZN(
        prince_inst_sbox_inst9_n9) );
  INV_X1 prince_inst_sbox_inst9_U4 ( .A(prince_inst_n28), .ZN(
        prince_inst_sbox_inst9_n8) );
  INV_X1 prince_inst_sbox_inst9_U3 ( .A(prince_inst_sbox_inst9_n8), .ZN(
        prince_inst_sbox_inst9_n6) );
  INV_X1 prince_inst_sbox_inst9_U2 ( .A(prince_inst_sbox_inst9_n8), .ZN(
        prince_inst_sbox_inst9_n7) );
  INV_X1 prince_inst_sbox_inst9_U1 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst9_n10) );
  NAND3_X1 prince_inst_sbox_inst9_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n68), .A3(prince_inst_sin_x[36]), 
        .ZN(prince_inst_sbox_inst9_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U25 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sbox_inst9_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst9_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst9_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst9_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst9_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n67), .A2(prince_inst_sin_x[38]), 
        .A3(prince_inst_sin_x[36]), .A4(prince_inst_sin_y[39]), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst9_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n61), .A2(prince_inst_sin_x[37]), 
        .A3(prince_inst_sin_x[38]), .ZN(prince_inst_sbox_inst9_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst9_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n66), .A3(prince_inst_sin_x[37]), 
        .A4(prince_inst_sin_x[36]), .ZN(prince_inst_sbox_inst9_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst9_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst9_xxxy_inst_n59), .B(prince_inst_sin_y[39]), .Z(
        prince_inst_sbox_inst9_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U18 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sin_x[37]), .ZN(prince_inst_sbox_inst9_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst9_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst9_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n65), .A2(prince_inst_sin_x[38]), 
        .ZN(prince_inst_sbox_inst9_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst9_xxxy_inst_U15 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sin_y[39]), .A3(prince_inst_sbox_inst9_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst9_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst9_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst9_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst9_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst9_xxxy_inst_U13 ( .A(prince_inst_sin_x[36]), 
        .B(prince_inst_sin_x[37]), .S(prince_inst_sbox_inst9_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst9_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst9_xxxy_inst_U12 ( .A(prince_inst_sin_y[39]), 
        .ZN(prince_inst_sbox_inst9_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U11 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sin_x[36]), .ZN(prince_inst_sbox_inst9_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst9_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst9_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst9_xxxy_inst_n60), .B(
        prince_inst_sbox_inst9_xxxy_inst_n53), .S(
        prince_inst_sbox_inst9_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst9_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U8 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sbox_inst9_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U7 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sin_y[39]), .ZN(prince_inst_sbox_inst9_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst9_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst9_t1_sh[0]), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst9_xxxy_inst_U5 ( .A(prince_inst_sin_x[38]), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U4 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sbox_inst9_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst9_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst9_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst9_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst9_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst9_xxxy_inst_U2 ( .A(prince_inst_sin_x[36]), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst9_xxxy_inst_U1 ( .A(prince_inst_sin_x[37]), .ZN(
        prince_inst_sbox_inst9_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst9_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst9_t1_sh[1]), .B(
        prince_inst_sbox_inst9_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst9_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst9_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst9_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst9_xxyx_inst_n52), .B(
        prince_inst_sbox_inst9_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst9_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U23 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst9_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst9_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n48), .A2(prince_inst_sin_x[39]), 
        .A3(prince_inst_sin_x[36]), .ZN(prince_inst_sbox_inst9_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n45), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst9_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst9_xxyx_inst_U18 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n46), .A2(prince_inst_sin_x[39]), 
        .A3(prince_inst_sin_x[37]), .ZN(prince_inst_sbox_inst9_xxyx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst9_t2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst9_xxyx_inst_U16 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sin_x[36]), .A3(prince_inst_sbox_inst9_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst9_xxyx_inst_n44) );
  OR2_X1 prince_inst_sbox_inst9_xxyx_inst_U15 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sbox_inst9_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst9_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst9_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst9_xxyx_inst_n54), .B(
        prince_inst_sbox_inst9_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst9_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U12 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sin_y[38]), .ZN(prince_inst_sbox_inst9_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst9_xxyx_inst_U11 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sbox_inst9_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst9_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst9_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst9_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst9_xxyx_inst_U10 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst9_xxyx_inst_U9 ( .A1(prince_inst_sin_x[39]), 
        .A2(prince_inst_sbox_inst9_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst9_xxyx_inst_U8 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sbox_inst9_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst9_xxyx_inst_U7 ( .A(prince_inst_sin_y[38]), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst9_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst9_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst9_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n53), .A2(prince_inst_sin_x[37]), 
        .A3(prince_inst_sin_y[38]), .A4(prince_inst_sin_x[36]), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst9_xxyx_inst_U4 ( .A(prince_inst_sin_x[39]), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst9_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst9_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst9_xxyx_inst_n43), .A3(prince_inst_sin_x[39]), 
        .A4(prince_inst_sin_y[38]), .ZN(prince_inst_sbox_inst9_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst9_xxyx_inst_U2 ( .A(prince_inst_sin_x[36]), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst9_xxyx_inst_U1 ( .A(prince_inst_sin_x[37]), .ZN(
        prince_inst_sbox_inst9_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst9_xyxx_inst_n74), .B(
        prince_inst_sbox_inst9_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst9_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst9_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst9_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst9_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U26 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sbox_inst9_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U25 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst9_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst9_xyxx_inst_n72), .B(
        prince_inst_sbox_inst9_s0_sh[2]), .S(
        prince_inst_sbox_inst9_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst9_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst9_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n74), .A2(prince_inst_sin_x[39]), 
        .ZN(prince_inst_sbox_inst9_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst9_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U21 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sbox_inst9_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst9_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst9_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst9_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst9_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst9_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst9_xyxx_inst_U15 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_x[36]), .ZN(prince_inst_sbox_inst9_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst9_xyxx_inst_U13 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U12 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_x[38]), .ZN(prince_inst_sbox_inst9_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst9_xyxx_inst_n58), .B(
        prince_inst_sbox_inst9_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst9_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst9_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst9_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst9_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst9_xyxx_inst_U9 ( .A(prince_inst_sin_x[39]), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst9_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n54), .A2(prince_inst_sin_x[36]), 
        .ZN(prince_inst_sbox_inst9_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst9_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst9_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst9_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst9_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst9_xyxx_inst_U5 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sbox_inst9_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst9_xyxx_inst_U4 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst9_xyxx_inst_U3 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sbox_inst9_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst9_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst9_xyxx_inst_U2 ( .A(prince_inst_sin_y[37]), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst9_xyxx_inst_U1 ( .A(prince_inst_sin_x[38]), .ZN(
        prince_inst_sbox_inst9_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst9_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst9_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst9_xyyy_inst_n59), .B(
        prince_inst_sbox_inst9_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst9_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst9_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst9_xyyy_inst_U25 ( .A1(prince_inst_sin_y[38]), 
        .A2(prince_inst_sin_y[39]), .A3(prince_inst_sbox_inst9_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst9_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U24 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sbox_inst9_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U23 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sbox_inst9_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst9_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst9_xyyy_inst_U19 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sin_y[38]), .A3(prince_inst_sbox_inst9_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst9_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst9_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst9_xyyy_inst_n49), .B(
        prince_inst_sbox_inst9_xyyy_inst_n48), .S(
        prince_inst_sbox_inst9_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst9_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst9_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst9_xyyy_inst_U16 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sbox_inst9_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst9_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst9_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst9_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst9_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst9_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst9_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst9_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst9_xyyy_inst_U12 ( .A(prince_inst_sin_y[39]), 
        .ZN(prince_inst_sbox_inst9_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst9_xyyy_inst_U11 ( .A1(prince_inst_sin_y[39]), 
        .A2(prince_inst_sbox_inst9_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst9_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst9_t1_sh[3]), .B(
        prince_inst_sbox_inst9_xyyy_inst_n48), .S(
        prince_inst_sbox_inst9_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst9_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst9_xyyy_inst_U9 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sbox_inst9_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst9_xyyy_inst_U8 ( .A1(prince_inst_sin_x[36]), 
        .A2(prince_inst_sin_y[39]), .ZN(prince_inst_sbox_inst9_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst9_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst9_t1_sh[3]), .ZN(prince_inst_sbox_inst9_s1_sh[3])
         );
  NAND2_X1 prince_inst_sbox_inst9_xyyy_inst_U6 ( .A1(prince_inst_sin_y[39]), 
        .A2(prince_inst_sbox_inst9_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst9_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst9_xyyy_inst_U4 ( .A(prince_inst_sin_y[37]), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst9_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst9_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst9_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst9_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst9_xyyy_inst_U2 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_x[36]), .ZN(prince_inst_sbox_inst9_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst9_xyyy_inst_U1 ( .A(prince_inst_sin_y[38]), .ZN(
        prince_inst_sbox_inst9_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst9_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U27 ( .A1(prince_inst_sin_y[36]), 
        .A2(prince_inst_sbox_inst9_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst9_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U24 ( .A1(prince_inst_sin_y[36]), 
        .A2(prince_inst_sbox_inst9_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst9_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U21 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst9_yxxx_inst_U19 ( .A(prince_inst_sin_x[39]), 
        .ZN(prince_inst_sbox_inst9_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst9_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst9_yxxx_inst_n52), .B(
        prince_inst_sbox_inst9_yxxx_inst_n51), .S(
        prince_inst_sbox_inst9_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst9_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n53), .A2(prince_inst_sin_x[39]), 
        .ZN(prince_inst_sbox_inst9_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst9_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n48), .A2(prince_inst_sin_y[36]), 
        .ZN(prince_inst_sbox_inst9_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n47), .A2(prince_inst_sin_x[39]), 
        .ZN(prince_inst_sbox_inst9_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U13 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sbox_inst9_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst9_yxxx_inst_n59), .B(
        prince_inst_sbox_inst9_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst9_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst9_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst9_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst9_yxxx_inst_U9 ( .A1(prince_inst_sin_x[37]), 
        .A2(prince_inst_sbox_inst9_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst9_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst9_yxxx_inst_U8 ( .A(prince_inst_sin_x[38]), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst9_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst9_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst9_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst9_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst9_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst9_yxxx_inst_U5 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sbox_inst9_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst9_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst9_yxxx_inst_U4 ( .A(prince_inst_sin_y[36]), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst9_yxxx_inst_U3 ( .A(prince_inst_sin_x[37]), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst9_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst9_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst9_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst9_yxxx_inst_U1 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst9_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst9_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst9_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst9_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst9_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n64), .A3(prince_inst_sin_y[39]), 
        .ZN(prince_inst_sbox_inst9_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst9_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n63), .A2(prince_inst_sin_y[38]), 
        .A3(prince_inst_sin_y[39]), .ZN(prince_inst_sbox_inst9_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst9_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst9_yxyy_inst_n62), .B(
        prince_inst_sbox_inst9_yxyy_inst_n61), .S(prince_inst_sin_y[36]), .Z(
        prince_inst_sbox_inst9_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst9_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst9_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst9_yxyy_inst_n64), .B(
        prince_inst_sbox_inst9_yxyy_inst_n60), .S(
        prince_inst_sbox_inst9_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst9_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst9_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst9_yxyy_inst_n62), .B(
        prince_inst_sbox_inst9_yxyy_inst_n54), .S(
        prince_inst_sbox_inst9_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst9_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst9_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst9_yxyy_inst_n53), .B(
        prince_inst_sbox_inst9_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst9_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst9_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst9_yxyy_inst_n68), .B(
        prince_inst_sbox_inst9_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst9_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U15 ( .A1(prince_inst_sin_y[39]), 
        .A2(prince_inst_sin_y[36]), .ZN(prince_inst_sbox_inst9_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst9_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst9_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst9_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst9_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst9_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst9_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst9_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst9_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n64), .A2(prince_inst_sin_y[38]), 
        .A3(prince_inst_sin_y[36]), .ZN(prince_inst_sbox_inst9_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst9_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U9 ( .A1(prince_inst_sin_y[39]), 
        .A2(prince_inst_sbox_inst9_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst9_yxyy_inst_U8 ( .A1(prince_inst_sin_y[38]), 
        .A2(prince_inst_sbox_inst9_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst9_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst9_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst9_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst9_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst9_yxyy_inst_U5 ( .A(prince_inst_sin_y[36]), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst9_yxyy_inst_U4 ( .A(prince_inst_sin_x[37]), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst9_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst9_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst9_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst9_yxyy_inst_U2 ( .A(prince_inst_sin_y[39]), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst9_yxyy_inst_U1 ( .A(prince_inst_sin_y[38]), .ZN(
        prince_inst_sbox_inst9_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst9_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U29 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sbox_inst9_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst9_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst9_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst9_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n75), .A2(prince_inst_sin_y[39]), 
        .A3(prince_inst_sbox_inst9_yyxy_inst_n70), .A4(prince_inst_sin_x[38]), 
        .ZN(prince_inst_sbox_inst9_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst9_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n69), .A3(prince_inst_sin_y[37]), 
        .A4(prince_inst_sbox_inst9_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst9_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst9_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst9_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst9_yyxy_inst_U23 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_x[38]), .A3(prince_inst_sin_y[36]), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst9_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n69), .A2(prince_inst_sin_y[37]), 
        .A3(prince_inst_sin_y[39]), .ZN(prince_inst_sbox_inst9_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst9_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n75), .A2(prince_inst_sin_x[38]), 
        .A3(prince_inst_sin_y[39]), .ZN(prince_inst_sbox_inst9_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst9_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst9_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst9_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n61), .A2(prince_inst_sin_x[38]), 
        .ZN(prince_inst_sbox_inst9_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst9_yyxy_inst_U18 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_y[39]), .A3(prince_inst_sbox_inst9_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst9_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst9_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst9_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst9_yyxy_inst_U16 ( .A1(prince_inst_sin_y[39]), 
        .A2(prince_inst_sbox_inst9_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst9_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst9_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst9_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n58), .A3(prince_inst_sin_y[36]), 
        .ZN(prince_inst_sbox_inst9_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst9_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst9_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst9_yyxy_inst_U13 ( .A1(prince_inst_sin_y[36]), 
        .A2(prince_inst_sbox_inst9_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst9_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst9_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst9_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst9_yyxy_inst_n54), .B(
        prince_inst_sbox_inst9_yyxy_inst_n55), .S(
        prince_inst_sbox_inst9_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst9_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst9_yyxy_inst_U9 ( .A(prince_inst_sin_x[38]), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n75), .A2(prince_inst_sin_y[39]), 
        .ZN(prince_inst_sbox_inst9_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst9_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst9_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst9_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U5 ( .A1(prince_inst_sin_x[38]), 
        .A2(prince_inst_sbox_inst9_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst9_yyxy_inst_U4 ( .A(prince_inst_sin_y[37]), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst9_yyxy_inst_U3 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sbox_inst9_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst9_yyxy_inst_U2 ( .A(prince_inst_sin_y[36]), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst9_yyxy_inst_U1 ( .A(prince_inst_sin_y[39]), .ZN(
        prince_inst_sbox_inst9_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst9_yyyx_inst_n58), .B(
        prince_inst_sbox_inst9_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst9_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst9_yyyx_inst_n56), .B(
        prince_inst_sbox_inst9_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst9_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst9_yyyx_inst_n54), .B(
        prince_inst_sbox_inst9_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst9_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst9_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst9_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst9_yyyx_inst_U21 ( .A1(prince_inst_sin_x[39]), 
        .A2(prince_inst_sbox_inst9_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst9_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst9_yyyx_inst_U20 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_y[38]), .A3(prince_inst_sbox_inst9_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst9_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst9_yyyx_inst_n50), .B(
        prince_inst_sbox_inst9_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst9_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst9_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n56), .A2(prince_inst_sin_y[38]), 
        .ZN(prince_inst_sbox_inst9_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst9_yyyx_inst_U17 ( .A1(prince_inst_sin_y[37]), 
        .A2(prince_inst_sin_y[36]), .A3(prince_inst_sin_y[38]), .ZN(
        prince_inst_sbox_inst9_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst9_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst9_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst9_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst9_yyyx_inst_U15 ( .A1(prince_inst_sin_x[39]), 
        .A2(prince_inst_sin_y[38]), .A3(prince_inst_sbox_inst9_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst9_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst9_yyyx_inst_U14 ( .A(prince_inst_sin_y[36]), 
        .ZN(prince_inst_sbox_inst9_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n58), .A2(prince_inst_sin_y[37]), 
        .ZN(prince_inst_sbox_inst9_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst9_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst9_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U11 ( .A1(prince_inst_sin_y[36]), 
        .A2(prince_inst_sbox_inst9_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst9_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst9_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst9_yyyx_inst_U9 ( .A1(prince_inst_sin_y[36]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst9_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst9_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst9_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst9_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n45), .A2(prince_inst_sin_y[36]), 
        .A3(prince_inst_sin_y[38]), .ZN(prince_inst_sbox_inst9_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst9_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst9_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst9_yyyx_inst_U4 ( .A1(prince_inst_sin_x[39]), 
        .A2(prince_inst_sin_y[38]), .ZN(prince_inst_sbox_inst9_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst9_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst9_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst9_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst9_yyyx_inst_U2 ( .A(prince_inst_sin_y[37]), .ZN(
        prince_inst_sbox_inst9_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst9_yyyx_inst_U1 ( .A1(prince_inst_sin_y[36]), 
        .A2(prince_inst_sin_x[39]), .ZN(prince_inst_sbox_inst9_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s00_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[0]), .B(prince_inst_sbox_inst9_s0_sh[0]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh0_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s01_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[1]), .B(prince_inst_sbox_inst9_s0_sh[1]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh0_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s02_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[2]), .B(prince_inst_sbox_inst9_s0_sh[2]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh0_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s03_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[3]), .B(prince_inst_sbox_inst9_s0_sh[3]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh0_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s04_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[4]), .B(prince_inst_sbox_inst9_s0_sh[4]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh0_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s05_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[5]), .B(prince_inst_sbox_inst9_s0_sh[5]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh0_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s06_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[6]), .B(prince_inst_sbox_inst9_s0_sh[6]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh0_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s07_U1 ( .A(
        prince_inst_sbox_inst9_t0_sh[7]), .B(prince_inst_sbox_inst9_s0_sh[7]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh0_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s10_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[0]), .B(prince_inst_sbox_inst9_s1_sh[0]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh1_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s11_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[1]), .B(prince_inst_sbox_inst9_s1_sh[1]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh1_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s12_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[2]), .B(prince_inst_sbox_inst9_s1_sh[2]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh1_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s13_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[3]), .B(prince_inst_sbox_inst9_s1_sh[3]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh1_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s14_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[4]), .B(prince_inst_sbox_inst9_s1_sh[4]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh1_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s15_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[5]), .B(prince_inst_sbox_inst9_s1_sh[5]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh1_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s16_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[6]), .B(prince_inst_sbox_inst9_s1_sh[6]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh1_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s17_U1 ( .A(
        prince_inst_sbox_inst9_t1_sh[7]), .B(prince_inst_sbox_inst9_s1_sh[7]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh1_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s20_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[0]), .B(prince_inst_sbox_inst9_s2_sh[0]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh2_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s21_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[1]), .B(prince_inst_sbox_inst9_s2_sh[1]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh2_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s22_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[2]), .B(prince_inst_sbox_inst9_s2_sh[2]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh2_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s23_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[3]), .B(prince_inst_sbox_inst9_s2_sh[3]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh2_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s24_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[4]), .B(prince_inst_sbox_inst9_s2_sh[4]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh2_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s25_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[5]), .B(prince_inst_sbox_inst9_s2_sh[5]), 
        .S(prince_inst_sbox_inst9_n6), .Z(prince_inst_sbox_inst9_sh2_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s26_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[6]), .B(prince_inst_sbox_inst9_s2_sh[6]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh2_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s27_U1 ( .A(
        prince_inst_sbox_inst9_t2_sh[7]), .B(prince_inst_sbox_inst9_s2_sh[7]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh2_tmp[7])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s30_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[0]), .B(prince_inst_sbox_inst9_s3_sh[0]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[0])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s31_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[1]), .B(prince_inst_sbox_inst9_s3_sh[1]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[1])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s32_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[2]), .B(prince_inst_sbox_inst9_s3_sh[2]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[2])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s33_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[3]), .B(prince_inst_sbox_inst9_s3_sh[3]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[3])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s34_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[4]), .B(prince_inst_sbox_inst9_s3_sh[4]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[4])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s35_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[5]), .B(prince_inst_sbox_inst9_s3_sh[5]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[5])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s36_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[6]), .B(prince_inst_sbox_inst9_s3_sh[6]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[6])
         );
  MUX2_X1 prince_inst_sbox_inst9_mux_s37_U1 ( .A(
        prince_inst_sbox_inst9_t3_sh[7]), .B(prince_inst_sbox_inst9_s3_sh[7]), 
        .S(prince_inst_sbox_inst9_n7), .Z(prince_inst_sbox_inst9_sh3_tmp[7])
         );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk0_U1 ( .A(r[80]), .B(
        prince_inst_sbox_inst9_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk1_U1 ( .A(r[81]), .B(
        prince_inst_sbox_inst9_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk2_U1 ( .A(r[82]), .B(
        prince_inst_sbox_inst9_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk3_U1 ( .A(r[83]), .B(
        prince_inst_sbox_inst9_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk4_U1 ( .A(r[80]), .B(
        prince_inst_sbox_inst9_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk5_U1 ( .A(r[81]), .B(
        prince_inst_sbox_inst9_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk6_U1 ( .A(r[82]), .B(
        prince_inst_sbox_inst9_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_msk7_U1 ( .A(r[83]), .B(
        prince_inst_sbox_inst9_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst9_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst9_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst9_c_inst0_ax_n5), .ZN(prince_inst_sout_x[36]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst9_c_inst0_y[1]), .B(
        prince_inst_sbox_inst9_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst9_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst9_c_inst0_y[2]), .B(
        prince_inst_sbox_inst9_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst9_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst9_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst9_c_inst0_ay_n5), .ZN(final_y[4]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst9_c_inst0_y[5]), .B(
        prince_inst_sbox_inst9_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst9_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst9_c_inst0_y[6]), .B(
        prince_inst_sbox_inst9_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst9_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk0_U1 ( .A(r[84]), .B(
        prince_inst_sbox_inst9_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk1_U1 ( .A(r[85]), .B(
        prince_inst_sbox_inst9_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk2_U1 ( .A(r[86]), .B(
        prince_inst_sbox_inst9_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk3_U1 ( .A(r[87]), .B(
        prince_inst_sbox_inst9_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk4_U1 ( .A(r[84]), .B(
        prince_inst_sbox_inst9_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk5_U1 ( .A(r[85]), .B(
        prince_inst_sbox_inst9_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk6_U1 ( .A(r[86]), .B(
        prince_inst_sbox_inst9_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_msk7_U1 ( .A(r[87]), .B(
        prince_inst_sbox_inst9_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst9_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst9_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst9_c_inst1_ax_n5), .ZN(prince_inst_sout_x[37]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst9_c_inst1_y[1]), .B(
        prince_inst_sbox_inst9_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst9_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst9_c_inst1_y[2]), .B(
        prince_inst_sbox_inst9_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst9_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst9_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst9_c_inst1_ay_n5), .ZN(final_y[5]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst9_c_inst1_y[5]), .B(
        prince_inst_sbox_inst9_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst9_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst9_c_inst1_y[6]), .B(
        prince_inst_sbox_inst9_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst9_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk0_U1 ( .A(r[88]), .B(
        prince_inst_sbox_inst9_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk1_U1 ( .A(r[89]), .B(
        prince_inst_sbox_inst9_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk2_U1 ( .A(r[90]), .B(
        prince_inst_sbox_inst9_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk3_U1 ( .A(r[91]), .B(
        prince_inst_sbox_inst9_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk4_U1 ( .A(r[88]), .B(
        prince_inst_sbox_inst9_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk5_U1 ( .A(r[89]), .B(
        prince_inst_sbox_inst9_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk6_U1 ( .A(r[90]), .B(
        prince_inst_sbox_inst9_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_msk7_U1 ( .A(r[91]), .B(
        prince_inst_sbox_inst9_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst9_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst9_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst9_c_inst2_ax_n5), .ZN(prince_inst_sout_x[38]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst9_c_inst2_y[1]), .B(
        prince_inst_sbox_inst9_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst9_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst9_c_inst2_y[2]), .B(
        prince_inst_sbox_inst9_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst9_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst9_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst9_c_inst2_ay_n5), .ZN(final_y[6]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst9_c_inst2_y[5]), .B(
        prince_inst_sbox_inst9_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst9_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst9_c_inst2_y[6]), .B(
        prince_inst_sbox_inst9_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst9_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk0_U1 ( .A(r[92]), .B(
        prince_inst_sbox_inst9_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk1_U1 ( .A(r[93]), .B(
        prince_inst_sbox_inst9_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk2_U1 ( .A(r[94]), .B(
        prince_inst_sbox_inst9_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk3_U1 ( .A(r[95]), .B(
        prince_inst_sbox_inst9_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk4_U1 ( .A(r[92]), .B(
        prince_inst_sbox_inst9_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk5_U1 ( .A(r[93]), .B(
        prince_inst_sbox_inst9_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk6_U1 ( .A(r[94]), .B(
        prince_inst_sbox_inst9_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_msk7_U1 ( .A(r[95]), .B(
        prince_inst_sbox_inst9_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst9_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst9_n9), .A2(prince_inst_sbox_inst9_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst9_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst9_n9), .ZN(
        prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst9_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst9_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst9_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst9_c_inst3_ax_n5), .ZN(prince_inst_sout_x[39]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst9_c_inst3_y[1]), .B(
        prince_inst_sbox_inst9_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst9_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst9_c_inst3_y[2]), .B(
        prince_inst_sbox_inst9_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst9_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst9_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst9_c_inst3_ay_n5), .ZN(final_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst9_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst9_c_inst3_y[5]), .B(
        prince_inst_sbox_inst9_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst9_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst9_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst9_c_inst3_y[6]), .B(
        prince_inst_sbox_inst9_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst9_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst10_U5 ( .A(prince_inst_sbox_inst10_n11), .ZN(
        prince_inst_sbox_inst10_n10) );
  INV_X1 prince_inst_sbox_inst10_U4 ( .A(prince_inst_n29), .ZN(
        prince_inst_sbox_inst10_n9) );
  INV_X1 prince_inst_sbox_inst10_U3 ( .A(prince_inst_sbox_inst10_n9), .ZN(
        prince_inst_sbox_inst10_n7) );
  INV_X1 prince_inst_sbox_inst10_U2 ( .A(prince_inst_sbox_inst10_n9), .ZN(
        prince_inst_sbox_inst10_n8) );
  INV_X1 prince_inst_sbox_inst10_U1 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst10_n11) );
  NAND3_X1 prince_inst_sbox_inst10_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n68), .A3(prince_inst_sin_x[40]), 
        .ZN(prince_inst_sbox_inst10_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst10_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U25 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sbox_inst10_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst10_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst10_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst10_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst10_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst10_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n67), .A2(prince_inst_sin_x[42]), 
        .A3(prince_inst_sin_x[40]), .A4(prince_inst_sin_y[43]), .ZN(
        prince_inst_sbox_inst10_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst10_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n61), .A2(prince_inst_sin_x[41]), 
        .A3(prince_inst_sin_x[42]), .ZN(prince_inst_sbox_inst10_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst10_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n66), .A3(prince_inst_sin_x[41]), 
        .A4(prince_inst_sin_x[40]), .ZN(prince_inst_sbox_inst10_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst10_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst10_xxxy_inst_n59), .B(prince_inst_sin_y[43]), .Z(
        prince_inst_sbox_inst10_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst10_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U18 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sin_x[41]), .ZN(prince_inst_sbox_inst10_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst10_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst10_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n65), .A2(prince_inst_sin_x[42]), 
        .ZN(prince_inst_sbox_inst10_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst10_xxxy_inst_U15 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sin_y[43]), .A3(prince_inst_sbox_inst10_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst10_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst10_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst10_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst10_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst10_xxxy_inst_U13 ( .A(prince_inst_sin_x[40]), 
        .B(prince_inst_sin_x[41]), .S(prince_inst_sbox_inst10_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst10_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst10_xxxy_inst_U12 ( .A(prince_inst_sin_y[43]), 
        .ZN(prince_inst_sbox_inst10_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U11 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sin_x[40]), .ZN(prince_inst_sbox_inst10_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst10_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst10_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst10_xxxy_inst_n60), .B(
        prince_inst_sbox_inst10_xxxy_inst_n53), .S(
        prince_inst_sbox_inst10_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst10_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U8 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sbox_inst10_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst10_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U7 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sin_y[43]), .ZN(prince_inst_sbox_inst10_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst10_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst10_t1_sh[0]), .ZN(
        prince_inst_sbox_inst10_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst10_xxxy_inst_U5 ( .A(prince_inst_sin_x[42]), 
        .ZN(prince_inst_sbox_inst10_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U4 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sbox_inst10_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst10_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst10_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst10_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst10_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst10_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst10_xxxy_inst_U2 ( .A(prince_inst_sin_x[40]), 
        .ZN(prince_inst_sbox_inst10_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst10_xxxy_inst_U1 ( .A(prince_inst_sin_x[41]), 
        .ZN(prince_inst_sbox_inst10_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst10_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst10_t1_sh[1]), .B(
        prince_inst_sbox_inst10_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst10_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst10_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst10_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst10_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst10_xxyx_inst_n52), .B(
        prince_inst_sbox_inst10_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst10_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U23 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst10_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst10_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n48), .A2(prince_inst_sin_x[43]), 
        .A3(prince_inst_sin_x[40]), .ZN(prince_inst_sbox_inst10_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst10_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst10_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst10_xxyx_inst_U18 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sbox_inst10_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst10_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst10_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst10_xxyx_inst_U16 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sin_x[40]), .A3(prince_inst_sbox_inst10_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst10_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst10_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n46), .A2(prince_inst_sin_x[43]), 
        .A3(prince_inst_sin_x[41]), .ZN(prince_inst_sbox_inst10_xxyx_inst_n44)
         );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst10_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst10_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst10_xxyx_inst_n54), .B(
        prince_inst_sbox_inst10_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst10_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U12 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sin_y[42]), .ZN(prince_inst_sbox_inst10_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst10_xxyx_inst_U11 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sbox_inst10_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst10_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst10_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst10_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst10_xxyx_inst_U10 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst10_xxyx_inst_U9 ( .A1(prince_inst_sin_x[43]), 
        .A2(prince_inst_sbox_inst10_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst10_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst10_xxyx_inst_U8 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sbox_inst10_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst10_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst10_xxyx_inst_U7 ( .A(prince_inst_sin_y[42]), 
        .ZN(prince_inst_sbox_inst10_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst10_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst10_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst10_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n53), .A2(prince_inst_sin_x[41]), 
        .A3(prince_inst_sin_y[42]), .A4(prince_inst_sin_x[40]), .ZN(
        prince_inst_sbox_inst10_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst10_xxyx_inst_U4 ( .A(prince_inst_sin_x[43]), 
        .ZN(prince_inst_sbox_inst10_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst10_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst10_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst10_xxyx_inst_n43), .A3(prince_inst_sin_x[43]), 
        .A4(prince_inst_sin_y[42]), .ZN(prince_inst_sbox_inst10_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst10_xxyx_inst_U2 ( .A(prince_inst_sin_x[40]), 
        .ZN(prince_inst_sbox_inst10_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst10_xxyx_inst_U1 ( .A(prince_inst_sin_x[41]), 
        .ZN(prince_inst_sbox_inst10_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst10_xyxx_inst_n74), .B(
        prince_inst_sbox_inst10_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst10_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst10_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst10_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst10_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U26 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sbox_inst10_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U25 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst10_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst10_xyxx_inst_n72), .B(
        prince_inst_sbox_inst10_s0_sh[2]), .S(
        prince_inst_sbox_inst10_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst10_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst10_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n74), .A2(prince_inst_sin_x[43]), 
        .ZN(prince_inst_sbox_inst10_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst10_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U21 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sbox_inst10_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst10_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst10_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst10_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst10_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst10_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst10_xyxx_inst_U15 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_x[40]), .ZN(prince_inst_sbox_inst10_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst10_xyxx_inst_U13 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U12 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_x[42]), .ZN(prince_inst_sbox_inst10_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst10_xyxx_inst_n58), .B(
        prince_inst_sbox_inst10_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst10_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst10_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst10_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst10_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst10_xyxx_inst_U9 ( .A(prince_inst_sin_x[43]), 
        .ZN(prince_inst_sbox_inst10_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst10_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n54), .A2(prince_inst_sin_x[40]), 
        .ZN(prince_inst_sbox_inst10_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst10_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst10_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst10_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst10_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst10_xyxx_inst_U5 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sbox_inst10_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst10_xyxx_inst_U4 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst10_xyxx_inst_U3 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sbox_inst10_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst10_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst10_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst10_xyxx_inst_U2 ( .A(prince_inst_sin_y[41]), 
        .ZN(prince_inst_sbox_inst10_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst10_xyxx_inst_U1 ( .A(prince_inst_sin_x[42]), 
        .ZN(prince_inst_sbox_inst10_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst10_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst10_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst10_xyyy_inst_n59), .B(
        prince_inst_sbox_inst10_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst10_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst10_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst10_xyyy_inst_U25 ( .A1(prince_inst_sin_y[42]), 
        .A2(prince_inst_sin_y[43]), .A3(prince_inst_sbox_inst10_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst10_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U24 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sbox_inst10_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U23 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sbox_inst10_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst10_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst10_xyyy_inst_U19 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sin_y[42]), .A3(prince_inst_sbox_inst10_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst10_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst10_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst10_xyyy_inst_n49), .B(
        prince_inst_sbox_inst10_xyyy_inst_n48), .S(
        prince_inst_sbox_inst10_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst10_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst10_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst10_xyyy_inst_U16 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sbox_inst10_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst10_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst10_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst10_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst10_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst10_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst10_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst10_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst10_xyyy_inst_U12 ( .A(prince_inst_sin_y[43]), 
        .ZN(prince_inst_sbox_inst10_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst10_xyyy_inst_U11 ( .A1(prince_inst_sin_y[43]), 
        .A2(prince_inst_sbox_inst10_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst10_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst10_t1_sh[3]), .B(
        prince_inst_sbox_inst10_xyyy_inst_n48), .S(
        prince_inst_sbox_inst10_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst10_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst10_xyyy_inst_U9 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sbox_inst10_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst10_xyyy_inst_U8 ( .A1(prince_inst_sin_x[40]), 
        .A2(prince_inst_sin_y[43]), .ZN(prince_inst_sbox_inst10_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst10_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst10_t1_sh[3]), .ZN(
        prince_inst_sbox_inst10_s1_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst10_xyyy_inst_U6 ( .A1(prince_inst_sin_y[43]), 
        .A2(prince_inst_sbox_inst10_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst10_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst10_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst10_xyyy_inst_U4 ( .A(prince_inst_sin_y[41]), 
        .ZN(prince_inst_sbox_inst10_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst10_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst10_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst10_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst10_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst10_xyyy_inst_U2 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_x[40]), .ZN(prince_inst_sbox_inst10_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst10_xyyy_inst_U1 ( .A(prince_inst_sin_y[42]), 
        .ZN(prince_inst_sbox_inst10_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst10_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U27 ( .A1(prince_inst_sin_y[40]), 
        .A2(prince_inst_sbox_inst10_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst10_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U24 ( .A1(prince_inst_sin_y[40]), 
        .A2(prince_inst_sbox_inst10_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst10_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U21 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst10_yxxx_inst_U19 ( .A(prince_inst_sin_x[43]), 
        .ZN(prince_inst_sbox_inst10_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst10_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst10_yxxx_inst_n52), .B(
        prince_inst_sbox_inst10_yxxx_inst_n51), .S(
        prince_inst_sbox_inst10_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst10_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n53), .A2(prince_inst_sin_x[43]), 
        .ZN(prince_inst_sbox_inst10_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst10_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n48), .A2(prince_inst_sin_y[40]), 
        .ZN(prince_inst_sbox_inst10_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n47), .A2(prince_inst_sin_x[43]), 
        .ZN(prince_inst_sbox_inst10_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U13 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sbox_inst10_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst10_yxxx_inst_n59), .B(
        prince_inst_sbox_inst10_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst10_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst10_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst10_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst10_yxxx_inst_U9 ( .A1(prince_inst_sin_x[41]), 
        .A2(prince_inst_sbox_inst10_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst10_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst10_yxxx_inst_U8 ( .A(prince_inst_sin_x[42]), 
        .ZN(prince_inst_sbox_inst10_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst10_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst10_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst10_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst10_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst10_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst10_yxxx_inst_U5 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sbox_inst10_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst10_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst10_yxxx_inst_U4 ( .A(prince_inst_sin_y[40]), 
        .ZN(prince_inst_sbox_inst10_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst10_yxxx_inst_U3 ( .A(prince_inst_sin_x[41]), 
        .ZN(prince_inst_sbox_inst10_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst10_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst10_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst10_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst10_yxxx_inst_U1 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst10_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst10_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst10_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst10_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst10_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n64), .A3(prince_inst_sin_y[43]), 
        .ZN(prince_inst_sbox_inst10_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst10_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n63), .A2(prince_inst_sin_y[42]), 
        .A3(prince_inst_sin_y[43]), .ZN(prince_inst_sbox_inst10_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst10_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst10_yxyy_inst_n62), .B(
        prince_inst_sbox_inst10_yxyy_inst_n61), .S(prince_inst_sin_y[40]), .Z(
        prince_inst_sbox_inst10_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst10_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst10_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst10_yxyy_inst_n64), .B(
        prince_inst_sbox_inst10_yxyy_inst_n60), .S(
        prince_inst_sbox_inst10_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst10_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst10_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst10_yxyy_inst_n62), .B(
        prince_inst_sbox_inst10_yxyy_inst_n54), .S(
        prince_inst_sbox_inst10_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst10_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst10_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst10_yxyy_inst_n53), .B(
        prince_inst_sbox_inst10_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst10_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst10_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst10_yxyy_inst_n68), .B(
        prince_inst_sbox_inst10_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst10_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U15 ( .A1(prince_inst_sin_y[43]), 
        .A2(prince_inst_sin_y[40]), .ZN(prince_inst_sbox_inst10_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst10_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst10_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst10_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst10_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst10_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst10_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst10_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst10_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n64), .A2(prince_inst_sin_y[42]), 
        .A3(prince_inst_sin_y[40]), .ZN(prince_inst_sbox_inst10_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst10_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U9 ( .A1(prince_inst_sin_y[43]), 
        .A2(prince_inst_sbox_inst10_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst10_yxyy_inst_U8 ( .A1(prince_inst_sin_y[42]), 
        .A2(prince_inst_sbox_inst10_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst10_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst10_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst10_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst10_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst10_yxyy_inst_U5 ( .A(prince_inst_sin_y[40]), 
        .ZN(prince_inst_sbox_inst10_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst10_yxyy_inst_U4 ( .A(prince_inst_sin_x[41]), 
        .ZN(prince_inst_sbox_inst10_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst10_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst10_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst10_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst10_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst10_yxyy_inst_U2 ( .A(prince_inst_sin_y[43]), 
        .ZN(prince_inst_sbox_inst10_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst10_yxyy_inst_U1 ( .A(prince_inst_sin_y[42]), 
        .ZN(prince_inst_sbox_inst10_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst10_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U29 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sbox_inst10_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst10_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst10_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst10_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n75), .A2(prince_inst_sin_y[43]), 
        .A3(prince_inst_sbox_inst10_yyxy_inst_n70), .A4(prince_inst_sin_x[42]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst10_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n69), .A3(prince_inst_sin_y[41]), 
        .A4(prince_inst_sbox_inst10_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst10_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst10_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst10_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst10_yyxy_inst_U23 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_x[42]), .A3(prince_inst_sin_y[40]), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst10_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n69), .A2(prince_inst_sin_y[41]), 
        .A3(prince_inst_sin_y[43]), .ZN(prince_inst_sbox_inst10_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst10_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n75), .A2(prince_inst_sin_x[42]), 
        .A3(prince_inst_sin_y[43]), .ZN(prince_inst_sbox_inst10_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst10_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst10_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst10_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n61), .A2(prince_inst_sin_x[42]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst10_yyxy_inst_U18 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_y[43]), .A3(prince_inst_sbox_inst10_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst10_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst10_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst10_yyxy_inst_U16 ( .A1(prince_inst_sin_y[43]), 
        .A2(prince_inst_sbox_inst10_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst10_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst10_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst10_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n58), .A3(prince_inst_sin_y[40]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst10_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst10_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst10_yyxy_inst_U13 ( .A1(prince_inst_sin_y[40]), 
        .A2(prince_inst_sbox_inst10_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst10_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst10_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst10_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst10_yyxy_inst_n54), .B(
        prince_inst_sbox_inst10_yyxy_inst_n55), .S(
        prince_inst_sbox_inst10_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst10_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst10_yyxy_inst_U9 ( .A(prince_inst_sin_x[42]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n75), .A2(prince_inst_sin_y[43]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst10_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst10_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst10_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U5 ( .A1(prince_inst_sin_x[42]), 
        .A2(prince_inst_sbox_inst10_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst10_yyxy_inst_U4 ( .A(prince_inst_sin_y[41]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst10_yyxy_inst_U3 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sbox_inst10_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst10_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst10_yyxy_inst_U2 ( .A(prince_inst_sin_y[40]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst10_yyxy_inst_U1 ( .A(prince_inst_sin_y[43]), 
        .ZN(prince_inst_sbox_inst10_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst10_yyyx_inst_n58), .B(
        prince_inst_sbox_inst10_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst10_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst10_yyyx_inst_n56), .B(
        prince_inst_sbox_inst10_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst10_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst10_yyyx_inst_n54), .B(
        prince_inst_sbox_inst10_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst10_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst10_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst10_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst10_yyyx_inst_U21 ( .A1(prince_inst_sin_x[43]), 
        .A2(prince_inst_sbox_inst10_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst10_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst10_yyyx_inst_U20 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_y[42]), .A3(prince_inst_sbox_inst10_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst10_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst10_yyyx_inst_n50), .B(
        prince_inst_sbox_inst10_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst10_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst10_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n56), .A2(prince_inst_sin_y[42]), 
        .ZN(prince_inst_sbox_inst10_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst10_yyyx_inst_U17 ( .A1(prince_inst_sin_y[41]), 
        .A2(prince_inst_sin_y[40]), .A3(prince_inst_sin_y[42]), .ZN(
        prince_inst_sbox_inst10_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst10_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst10_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst10_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst10_yyyx_inst_U15 ( .A1(prince_inst_sin_x[43]), 
        .A2(prince_inst_sin_y[42]), .A3(prince_inst_sbox_inst10_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst10_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst10_yyyx_inst_U14 ( .A(prince_inst_sin_y[40]), 
        .ZN(prince_inst_sbox_inst10_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n58), .A2(prince_inst_sin_y[41]), 
        .ZN(prince_inst_sbox_inst10_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst10_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst10_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U11 ( .A1(prince_inst_sin_y[40]), 
        .A2(prince_inst_sbox_inst10_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst10_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst10_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst10_yyyx_inst_U9 ( .A1(prince_inst_sin_y[40]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst10_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst10_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst10_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst10_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n45), .A2(prince_inst_sin_y[40]), 
        .A3(prince_inst_sin_y[42]), .ZN(prince_inst_sbox_inst10_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst10_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst10_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst10_yyyx_inst_U4 ( .A1(prince_inst_sin_x[43]), 
        .A2(prince_inst_sin_y[42]), .ZN(prince_inst_sbox_inst10_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst10_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst10_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst10_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst10_yyyx_inst_U2 ( .A(prince_inst_sin_y[41]), 
        .ZN(prince_inst_sbox_inst10_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst10_yyyx_inst_U1 ( .A1(prince_inst_sin_y[40]), 
        .A2(prince_inst_sin_x[43]), .ZN(prince_inst_sbox_inst10_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst10_mux_s00_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[0]), .B(prince_inst_sbox_inst10_s0_sh[0]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh0_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s01_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[1]), .B(prince_inst_sbox_inst10_s0_sh[1]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh0_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s02_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[2]), .B(prince_inst_sbox_inst10_s0_sh[2]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh0_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s03_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[3]), .B(prince_inst_sbox_inst10_s0_sh[3]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh0_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s04_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[4]), .B(prince_inst_sbox_inst10_s0_sh[4]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh0_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s05_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[5]), .B(prince_inst_sbox_inst10_s0_sh[5]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh0_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s06_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[6]), .B(prince_inst_sbox_inst10_s0_sh[6]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh0_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s07_U1 ( .A(
        prince_inst_sbox_inst10_t0_sh[7]), .B(prince_inst_sbox_inst10_s0_sh[7]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh0_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s10_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[0]), .B(prince_inst_sbox_inst10_s1_sh[0]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh1_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s11_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[1]), .B(prince_inst_sbox_inst10_s1_sh[1]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh1_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s12_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[2]), .B(prince_inst_sbox_inst10_s1_sh[2]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh1_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s13_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[3]), .B(prince_inst_sbox_inst10_s1_sh[3]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh1_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s14_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[4]), .B(prince_inst_sbox_inst10_s1_sh[4]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh1_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s15_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[5]), .B(prince_inst_sbox_inst10_s1_sh[5]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh1_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s16_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[6]), .B(prince_inst_sbox_inst10_s1_sh[6]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh1_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s17_U1 ( .A(
        prince_inst_sbox_inst10_t1_sh[7]), .B(prince_inst_sbox_inst10_s1_sh[7]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh1_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s20_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[0]), .B(prince_inst_sbox_inst10_s2_sh[0]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh2_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s21_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[1]), .B(prince_inst_sbox_inst10_s2_sh[1]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh2_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s22_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[2]), .B(prince_inst_sbox_inst10_s2_sh[2]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh2_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s23_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[3]), .B(prince_inst_sbox_inst10_s2_sh[3]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh2_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s24_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[4]), .B(prince_inst_sbox_inst10_s2_sh[4]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh2_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s25_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[5]), .B(prince_inst_sbox_inst10_s2_sh[5]), .S(prince_inst_n29), .Z(prince_inst_sbox_inst10_sh2_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s26_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[6]), .B(prince_inst_sbox_inst10_s2_sh[6]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh2_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s27_U1 ( .A(
        prince_inst_sbox_inst10_t2_sh[7]), .B(prince_inst_sbox_inst10_s2_sh[7]), .S(prince_inst_sbox_inst10_n7), .Z(prince_inst_sbox_inst10_sh2_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s30_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[0]), .B(prince_inst_sbox_inst10_s3_sh[0]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s31_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[1]), .B(prince_inst_sbox_inst10_s3_sh[1]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s32_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[2]), .B(prince_inst_sbox_inst10_s3_sh[2]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s33_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[3]), .B(prince_inst_sbox_inst10_s3_sh[3]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s34_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[4]), .B(prince_inst_sbox_inst10_s3_sh[4]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s35_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[5]), .B(prince_inst_sbox_inst10_s3_sh[5]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s36_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[6]), .B(prince_inst_sbox_inst10_s3_sh[6]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst10_mux_s37_U1 ( .A(
        prince_inst_sbox_inst10_t3_sh[7]), .B(prince_inst_sbox_inst10_s3_sh[7]), .S(prince_inst_sbox_inst10_n8), .Z(prince_inst_sbox_inst10_sh3_tmp[7]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk0_U1 ( .A(r[96]), .B(
        prince_inst_sbox_inst10_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[0]), .ZN(prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk1_U1 ( .A(r[97]), .B(
        prince_inst_sbox_inst10_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[1]), .ZN(prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk2_U1 ( .A(r[98]), .B(
        prince_inst_sbox_inst10_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[2]), .ZN(prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk3_U1 ( .A(r[99]), .B(
        prince_inst_sbox_inst10_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[3]), .ZN(prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk4_U1 ( .A(r[96]), .B(
        prince_inst_sbox_inst10_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[4]), .ZN(prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk5_U1 ( .A(r[97]), .B(
        prince_inst_sbox_inst10_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[5]), .ZN(prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk6_U1 ( .A(r[98]), .B(
        prince_inst_sbox_inst10_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[6]), .ZN(prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_msk7_U1 ( .A(r[99]), .B(
        prince_inst_sbox_inst10_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst10_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst0_y[7]), .ZN(prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst10_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst10_c_inst0_ax_n5), .ZN(prince_inst_sout_x[40]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst10_c_inst0_y[1]), .B(
        prince_inst_sbox_inst10_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst10_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst10_c_inst0_y[2]), .B(
        prince_inst_sbox_inst10_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst10_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst10_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst10_c_inst0_ay_n5), .ZN(final_y[56]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst10_c_inst0_y[5]), .B(
        prince_inst_sbox_inst10_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst10_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst10_c_inst0_y[6]), .B(
        prince_inst_sbox_inst10_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst10_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk0_U1 ( .A(r[100]), .B(
        prince_inst_sbox_inst10_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[0]), .ZN(prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk1_U1 ( .A(r[101]), .B(
        prince_inst_sbox_inst10_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[1]), .ZN(prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk2_U1 ( .A(r[102]), .B(
        prince_inst_sbox_inst10_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[2]), .ZN(prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk3_U1 ( .A(r[103]), .B(
        prince_inst_sbox_inst10_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[3]), .ZN(prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk4_U1 ( .A(r[100]), .B(
        prince_inst_sbox_inst10_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[4]), .ZN(prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk5_U1 ( .A(r[101]), .B(
        prince_inst_sbox_inst10_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[5]), .ZN(prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk6_U1 ( .A(r[102]), .B(
        prince_inst_sbox_inst10_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[6]), .ZN(prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_msk7_U1 ( .A(r[103]), .B(
        prince_inst_sbox_inst10_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst10_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst1_y[7]), .ZN(prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst10_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst10_c_inst1_ax_n5), .ZN(prince_inst_sout_x[41]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst10_c_inst1_y[1]), .B(
        prince_inst_sbox_inst10_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst10_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst10_c_inst1_y[2]), .B(
        prince_inst_sbox_inst10_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst10_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst10_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst10_c_inst1_ay_n5), .ZN(final_y[57]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst10_c_inst1_y[5]), .B(
        prince_inst_sbox_inst10_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst10_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst10_c_inst1_y[6]), .B(
        prince_inst_sbox_inst10_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst10_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk0_U1 ( .A(r[104]), .B(
        prince_inst_sbox_inst10_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[0]), .ZN(prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk1_U1 ( .A(r[105]), .B(
        prince_inst_sbox_inst10_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[1]), .ZN(prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk2_U1 ( .A(r[106]), .B(
        prince_inst_sbox_inst10_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[2]), .ZN(prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk3_U1 ( .A(r[107]), .B(
        prince_inst_sbox_inst10_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[3]), .ZN(prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk4_U1 ( .A(r[104]), .B(
        prince_inst_sbox_inst10_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[4]), .ZN(prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk5_U1 ( .A(r[105]), .B(
        prince_inst_sbox_inst10_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[5]), .ZN(prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk6_U1 ( .A(r[106]), .B(
        prince_inst_sbox_inst10_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[6]), .ZN(prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_msk7_U1 ( .A(r[107]), .B(
        prince_inst_sbox_inst10_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst10_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst2_y[7]), .ZN(prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst10_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst10_c_inst2_ax_n5), .ZN(prince_inst_sout_x[42]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst10_c_inst2_y[1]), .B(
        prince_inst_sbox_inst10_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst10_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst10_c_inst2_y[2]), .B(
        prince_inst_sbox_inst10_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst10_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst10_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst10_c_inst2_ay_n5), .ZN(final_y[58]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst10_c_inst2_y[5]), .B(
        prince_inst_sbox_inst10_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst10_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst10_c_inst2_y[6]), .B(
        prince_inst_sbox_inst10_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst10_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk0_U1 ( .A(r[108]), .B(
        prince_inst_sbox_inst10_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[0]), .ZN(prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk1_U1 ( .A(r[109]), .B(
        prince_inst_sbox_inst10_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[1]), .ZN(prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk2_U1 ( .A(r[110]), .B(
        prince_inst_sbox_inst10_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[2]), .ZN(prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk3_U1 ( .A(r[111]), .B(
        prince_inst_sbox_inst10_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[3]), .ZN(prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk4_U1 ( .A(r[108]), .B(
        prince_inst_sbox_inst10_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[4]), .ZN(prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk5_U1 ( .A(r[109]), .B(
        prince_inst_sbox_inst10_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[5]), .ZN(prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk6_U1 ( .A(r[110]), .B(
        prince_inst_sbox_inst10_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[6]), .ZN(prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_msk7_U1 ( .A(r[111]), .B(
        prince_inst_sbox_inst10_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst10_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst10_n10), .A2(prince_inst_sbox_inst10_c_inst3_y[7]), .ZN(prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst10_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst10_n10), .ZN(
        prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst10_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst10_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst10_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst10_c_inst3_ax_n5), .ZN(prince_inst_sout_x[43]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst10_c_inst3_y[1]), .B(
        prince_inst_sbox_inst10_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst10_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst10_c_inst3_y[2]), .B(
        prince_inst_sbox_inst10_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst10_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst10_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst10_c_inst3_ay_n5), .ZN(final_y[59]) );
  XNOR2_X1 prince_inst_sbox_inst10_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst10_c_inst3_y[5]), .B(
        prince_inst_sbox_inst10_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst10_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst10_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst10_c_inst3_y[6]), .B(
        prince_inst_sbox_inst10_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst10_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst11_U7 ( .A(prince_inst_sbox_inst11_n13), .ZN(
        prince_inst_sbox_inst11_n12) );
  INV_X1 prince_inst_sbox_inst11_U6 ( .A(prince_inst_n33), .ZN(
        prince_inst_sbox_inst11_n11) );
  INV_X1 prince_inst_sbox_inst11_U5 ( .A(prince_inst_sbox_inst11_n11), .ZN(
        prince_inst_sbox_inst11_n9) );
  INV_X1 prince_inst_sbox_inst11_U4 ( .A(prince_inst_sbox_inst11_n11), .ZN(
        prince_inst_sbox_inst11_n10) );
  INV_X1 prince_inst_sbox_inst11_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst11_n13) );
  INV_X1 prince_inst_sbox_inst11_U2 ( .A(rst), .ZN(prince_inst_sbox_inst11_n8)
         );
  INV_X2 prince_inst_sbox_inst11_U1 ( .A(prince_inst_sbox_inst11_n8), .ZN(
        prince_inst_sbox_inst11_n7) );
  NAND3_X1 prince_inst_sbox_inst11_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n68), .A3(prince_inst_sin_x[44]), 
        .ZN(prince_inst_sbox_inst11_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst11_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U25 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sbox_inst11_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst11_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst11_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst11_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst11_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst11_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n67), .A2(prince_inst_sin_x[46]), 
        .A3(prince_inst_sin_x[44]), .A4(prince_inst_sin_y[47]), .ZN(
        prince_inst_sbox_inst11_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst11_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n61), .A2(prince_inst_sin_x[45]), 
        .A3(prince_inst_sin_x[46]), .ZN(prince_inst_sbox_inst11_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst11_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n66), .A3(prince_inst_sin_x[45]), 
        .A4(prince_inst_sin_x[44]), .ZN(prince_inst_sbox_inst11_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst11_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst11_xxxy_inst_n59), .B(prince_inst_sin_y[47]), .Z(
        prince_inst_sbox_inst11_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst11_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U18 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sin_x[45]), .ZN(prince_inst_sbox_inst11_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst11_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst11_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n65), .A2(prince_inst_sin_x[46]), 
        .ZN(prince_inst_sbox_inst11_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst11_xxxy_inst_U15 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sin_y[47]), .A3(prince_inst_sbox_inst11_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst11_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst11_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst11_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst11_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst11_xxxy_inst_U13 ( .A(prince_inst_sin_x[44]), 
        .B(prince_inst_sin_x[45]), .S(prince_inst_sbox_inst11_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst11_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst11_xxxy_inst_U12 ( .A(prince_inst_sin_y[47]), 
        .ZN(prince_inst_sbox_inst11_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U11 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sin_x[44]), .ZN(prince_inst_sbox_inst11_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst11_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst11_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst11_xxxy_inst_n60), .B(
        prince_inst_sbox_inst11_xxxy_inst_n53), .S(
        prince_inst_sbox_inst11_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst11_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U8 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sbox_inst11_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst11_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U7 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sin_y[47]), .ZN(prince_inst_sbox_inst11_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst11_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst11_t1_sh[0]), .ZN(
        prince_inst_sbox_inst11_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst11_xxxy_inst_U5 ( .A(prince_inst_sin_x[46]), 
        .ZN(prince_inst_sbox_inst11_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U4 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sbox_inst11_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst11_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst11_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst11_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst11_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst11_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst11_xxxy_inst_U2 ( .A(prince_inst_sin_x[44]), 
        .ZN(prince_inst_sbox_inst11_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst11_xxxy_inst_U1 ( .A(prince_inst_sin_x[45]), 
        .ZN(prince_inst_sbox_inst11_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst11_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst11_t1_sh[1]), .B(
        prince_inst_sbox_inst11_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst11_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst11_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst11_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst11_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst11_xxyx_inst_n52), .B(
        prince_inst_sbox_inst11_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst11_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U23 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst11_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst11_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n48), .A2(prince_inst_sin_x[47]), 
        .A3(prince_inst_sin_x[44]), .ZN(prince_inst_sbox_inst11_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst11_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst11_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst11_xxyx_inst_U18 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sbox_inst11_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst11_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst11_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst11_xxyx_inst_U16 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sin_x[44]), .A3(prince_inst_sbox_inst11_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst11_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst11_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n46), .A2(prince_inst_sin_x[47]), 
        .A3(prince_inst_sin_x[45]), .ZN(prince_inst_sbox_inst11_xxyx_inst_n44)
         );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst11_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst11_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst11_xxyx_inst_n54), .B(
        prince_inst_sbox_inst11_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst11_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U12 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sin_y[46]), .ZN(prince_inst_sbox_inst11_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst11_xxyx_inst_U11 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sbox_inst11_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst11_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst11_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst11_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst11_xxyx_inst_U10 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst11_xxyx_inst_U9 ( .A1(prince_inst_sin_x[47]), 
        .A2(prince_inst_sbox_inst11_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst11_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst11_xxyx_inst_U8 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sbox_inst11_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst11_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst11_xxyx_inst_U7 ( .A(prince_inst_sin_y[46]), 
        .ZN(prince_inst_sbox_inst11_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst11_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst11_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst11_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n53), .A2(prince_inst_sin_x[45]), 
        .A3(prince_inst_sin_y[46]), .A4(prince_inst_sin_x[44]), .ZN(
        prince_inst_sbox_inst11_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst11_xxyx_inst_U4 ( .A(prince_inst_sin_x[47]), 
        .ZN(prince_inst_sbox_inst11_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst11_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst11_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst11_xxyx_inst_n43), .A3(prince_inst_sin_x[47]), 
        .A4(prince_inst_sin_y[46]), .ZN(prince_inst_sbox_inst11_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst11_xxyx_inst_U2 ( .A(prince_inst_sin_x[44]), 
        .ZN(prince_inst_sbox_inst11_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst11_xxyx_inst_U1 ( .A(prince_inst_sin_x[45]), 
        .ZN(prince_inst_sbox_inst11_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst11_xyxx_inst_n74), .B(
        prince_inst_sbox_inst11_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst11_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst11_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst11_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst11_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U26 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sbox_inst11_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U25 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst11_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst11_xyxx_inst_n72), .B(
        prince_inst_sbox_inst11_s0_sh[2]), .S(
        prince_inst_sbox_inst11_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst11_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst11_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n74), .A2(prince_inst_sin_x[47]), 
        .ZN(prince_inst_sbox_inst11_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst11_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U21 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sbox_inst11_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst11_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst11_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst11_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst11_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst11_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst11_xyxx_inst_U15 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_x[44]), .ZN(prince_inst_sbox_inst11_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst11_xyxx_inst_U13 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U12 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_x[46]), .ZN(prince_inst_sbox_inst11_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst11_xyxx_inst_n58), .B(
        prince_inst_sbox_inst11_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst11_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst11_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst11_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst11_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst11_xyxx_inst_U9 ( .A(prince_inst_sin_x[47]), 
        .ZN(prince_inst_sbox_inst11_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst11_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n54), .A2(prince_inst_sin_x[44]), 
        .ZN(prince_inst_sbox_inst11_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst11_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst11_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst11_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst11_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst11_xyxx_inst_U5 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sbox_inst11_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst11_xyxx_inst_U4 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst11_xyxx_inst_U3 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sbox_inst11_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst11_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst11_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst11_xyxx_inst_U2 ( .A(prince_inst_sin_y[45]), 
        .ZN(prince_inst_sbox_inst11_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst11_xyxx_inst_U1 ( .A(prince_inst_sin_x[46]), 
        .ZN(prince_inst_sbox_inst11_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst11_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst11_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst11_xyyy_inst_n59), .B(
        prince_inst_sbox_inst11_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst11_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst11_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst11_xyyy_inst_U25 ( .A1(prince_inst_sin_y[46]), 
        .A2(prince_inst_sin_y[47]), .A3(prince_inst_sbox_inst11_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst11_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U24 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sbox_inst11_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U23 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sbox_inst11_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst11_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst11_xyyy_inst_U19 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sin_y[46]), .A3(prince_inst_sbox_inst11_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst11_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst11_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst11_xyyy_inst_n49), .B(
        prince_inst_sbox_inst11_xyyy_inst_n48), .S(
        prince_inst_sbox_inst11_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst11_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst11_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst11_xyyy_inst_U16 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sbox_inst11_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst11_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst11_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst11_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst11_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst11_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst11_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst11_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst11_xyyy_inst_U12 ( .A(prince_inst_sin_y[47]), 
        .ZN(prince_inst_sbox_inst11_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst11_xyyy_inst_U11 ( .A1(prince_inst_sin_y[47]), 
        .A2(prince_inst_sbox_inst11_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst11_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst11_t1_sh[3]), .B(
        prince_inst_sbox_inst11_xyyy_inst_n48), .S(
        prince_inst_sbox_inst11_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst11_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst11_xyyy_inst_U9 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sbox_inst11_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst11_xyyy_inst_U8 ( .A1(prince_inst_sin_x[44]), 
        .A2(prince_inst_sin_y[47]), .ZN(prince_inst_sbox_inst11_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst11_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst11_t1_sh[3]), .ZN(
        prince_inst_sbox_inst11_s1_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst11_xyyy_inst_U6 ( .A1(prince_inst_sin_y[47]), 
        .A2(prince_inst_sbox_inst11_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst11_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst11_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst11_xyyy_inst_U4 ( .A(prince_inst_sin_y[45]), 
        .ZN(prince_inst_sbox_inst11_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst11_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst11_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst11_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst11_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst11_xyyy_inst_U2 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_x[44]), .ZN(prince_inst_sbox_inst11_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst11_xyyy_inst_U1 ( .A(prince_inst_sin_y[46]), 
        .ZN(prince_inst_sbox_inst11_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst11_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U27 ( .A1(prince_inst_sin_y[44]), 
        .A2(prince_inst_sbox_inst11_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst11_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U24 ( .A1(prince_inst_sin_y[44]), 
        .A2(prince_inst_sbox_inst11_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst11_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U21 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst11_yxxx_inst_U19 ( .A(prince_inst_sin_x[47]), 
        .ZN(prince_inst_sbox_inst11_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst11_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst11_yxxx_inst_n52), .B(
        prince_inst_sbox_inst11_yxxx_inst_n51), .S(
        prince_inst_sbox_inst11_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst11_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n53), .A2(prince_inst_sin_x[47]), 
        .ZN(prince_inst_sbox_inst11_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst11_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n48), .A2(prince_inst_sin_y[44]), 
        .ZN(prince_inst_sbox_inst11_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n47), .A2(prince_inst_sin_x[47]), 
        .ZN(prince_inst_sbox_inst11_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U13 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sbox_inst11_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst11_yxxx_inst_n59), .B(
        prince_inst_sbox_inst11_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst11_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst11_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst11_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst11_yxxx_inst_U9 ( .A1(prince_inst_sin_x[45]), 
        .A2(prince_inst_sbox_inst11_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst11_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst11_yxxx_inst_U8 ( .A(prince_inst_sin_x[46]), 
        .ZN(prince_inst_sbox_inst11_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst11_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst11_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst11_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst11_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst11_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst11_yxxx_inst_U5 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sbox_inst11_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst11_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst11_yxxx_inst_U4 ( .A(prince_inst_sin_y[44]), 
        .ZN(prince_inst_sbox_inst11_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst11_yxxx_inst_U3 ( .A(prince_inst_sin_x[45]), 
        .ZN(prince_inst_sbox_inst11_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst11_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst11_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst11_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst11_yxxx_inst_U1 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst11_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst11_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst11_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst11_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst11_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n64), .A3(prince_inst_sin_y[47]), 
        .ZN(prince_inst_sbox_inst11_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst11_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n63), .A2(prince_inst_sin_y[46]), 
        .A3(prince_inst_sin_y[47]), .ZN(prince_inst_sbox_inst11_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst11_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst11_yxyy_inst_n62), .B(
        prince_inst_sbox_inst11_yxyy_inst_n61), .S(prince_inst_sin_y[44]), .Z(
        prince_inst_sbox_inst11_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst11_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst11_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst11_yxyy_inst_n64), .B(
        prince_inst_sbox_inst11_yxyy_inst_n60), .S(
        prince_inst_sbox_inst11_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst11_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst11_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst11_yxyy_inst_n62), .B(
        prince_inst_sbox_inst11_yxyy_inst_n54), .S(
        prince_inst_sbox_inst11_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst11_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst11_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst11_yxyy_inst_n53), .B(
        prince_inst_sbox_inst11_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst11_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst11_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst11_yxyy_inst_n68), .B(
        prince_inst_sbox_inst11_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst11_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U15 ( .A1(prince_inst_sin_y[47]), 
        .A2(prince_inst_sin_y[44]), .ZN(prince_inst_sbox_inst11_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst11_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst11_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst11_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst11_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst11_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst11_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst11_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst11_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n64), .A2(prince_inst_sin_y[46]), 
        .A3(prince_inst_sin_y[44]), .ZN(prince_inst_sbox_inst11_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst11_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U9 ( .A1(prince_inst_sin_y[47]), 
        .A2(prince_inst_sbox_inst11_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst11_yxyy_inst_U8 ( .A1(prince_inst_sin_y[46]), 
        .A2(prince_inst_sbox_inst11_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst11_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst11_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst11_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst11_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst11_yxyy_inst_U5 ( .A(prince_inst_sin_y[44]), 
        .ZN(prince_inst_sbox_inst11_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst11_yxyy_inst_U4 ( .A(prince_inst_sin_x[45]), 
        .ZN(prince_inst_sbox_inst11_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst11_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst11_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst11_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst11_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst11_yxyy_inst_U2 ( .A(prince_inst_sin_y[47]), 
        .ZN(prince_inst_sbox_inst11_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst11_yxyy_inst_U1 ( .A(prince_inst_sin_y[46]), 
        .ZN(prince_inst_sbox_inst11_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst11_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U29 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sbox_inst11_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst11_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst11_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst11_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n75), .A2(prince_inst_sin_y[47]), 
        .A3(prince_inst_sbox_inst11_yyxy_inst_n70), .A4(prince_inst_sin_x[46]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst11_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n69), .A3(prince_inst_sin_y[45]), 
        .A4(prince_inst_sbox_inst11_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst11_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst11_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst11_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst11_yyxy_inst_U23 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_x[46]), .A3(prince_inst_sin_y[44]), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst11_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n69), .A2(prince_inst_sin_y[45]), 
        .A3(prince_inst_sin_y[47]), .ZN(prince_inst_sbox_inst11_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst11_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n75), .A2(prince_inst_sin_x[46]), 
        .A3(prince_inst_sin_y[47]), .ZN(prince_inst_sbox_inst11_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst11_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst11_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst11_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n61), .A2(prince_inst_sin_x[46]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst11_yyxy_inst_U18 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_y[47]), .A3(prince_inst_sbox_inst11_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst11_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst11_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst11_yyxy_inst_U16 ( .A1(prince_inst_sin_y[47]), 
        .A2(prince_inst_sbox_inst11_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst11_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst11_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst11_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n58), .A3(prince_inst_sin_y[44]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst11_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst11_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst11_yyxy_inst_U13 ( .A1(prince_inst_sin_y[44]), 
        .A2(prince_inst_sbox_inst11_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst11_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst11_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst11_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst11_yyxy_inst_n54), .B(
        prince_inst_sbox_inst11_yyxy_inst_n55), .S(
        prince_inst_sbox_inst11_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst11_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst11_yyxy_inst_U9 ( .A(prince_inst_sin_x[46]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n75), .A2(prince_inst_sin_y[47]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst11_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst11_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst11_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U5 ( .A1(prince_inst_sin_x[46]), 
        .A2(prince_inst_sbox_inst11_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst11_yyxy_inst_U4 ( .A(prince_inst_sin_y[45]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst11_yyxy_inst_U3 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sbox_inst11_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst11_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst11_yyxy_inst_U2 ( .A(prince_inst_sin_y[44]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst11_yyxy_inst_U1 ( .A(prince_inst_sin_y[47]), 
        .ZN(prince_inst_sbox_inst11_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst11_yyyx_inst_n58), .B(
        prince_inst_sbox_inst11_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst11_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst11_yyyx_inst_n56), .B(
        prince_inst_sbox_inst11_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst11_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst11_yyyx_inst_n54), .B(
        prince_inst_sbox_inst11_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst11_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst11_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst11_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst11_yyyx_inst_U21 ( .A1(prince_inst_sin_x[47]), 
        .A2(prince_inst_sbox_inst11_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst11_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst11_yyyx_inst_U20 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_y[46]), .A3(prince_inst_sbox_inst11_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst11_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst11_yyyx_inst_n50), .B(
        prince_inst_sbox_inst11_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst11_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst11_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n56), .A2(prince_inst_sin_y[46]), 
        .ZN(prince_inst_sbox_inst11_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst11_yyyx_inst_U17 ( .A1(prince_inst_sin_y[45]), 
        .A2(prince_inst_sin_y[44]), .A3(prince_inst_sin_y[46]), .ZN(
        prince_inst_sbox_inst11_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst11_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst11_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst11_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst11_yyyx_inst_U15 ( .A1(prince_inst_sin_x[47]), 
        .A2(prince_inst_sin_y[46]), .A3(prince_inst_sbox_inst11_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst11_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst11_yyyx_inst_U14 ( .A(prince_inst_sin_y[44]), 
        .ZN(prince_inst_sbox_inst11_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n58), .A2(prince_inst_sin_y[45]), 
        .ZN(prince_inst_sbox_inst11_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst11_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst11_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U11 ( .A1(prince_inst_sin_y[44]), 
        .A2(prince_inst_sbox_inst11_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst11_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst11_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst11_yyyx_inst_U9 ( .A1(prince_inst_sin_y[44]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst11_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst11_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst11_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst11_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n45), .A2(prince_inst_sin_y[44]), 
        .A3(prince_inst_sin_y[46]), .ZN(prince_inst_sbox_inst11_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst11_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst11_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst11_yyyx_inst_U4 ( .A1(prince_inst_sin_x[47]), 
        .A2(prince_inst_sin_y[46]), .ZN(prince_inst_sbox_inst11_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst11_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst11_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst11_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst11_yyyx_inst_U2 ( .A(prince_inst_sin_y[45]), 
        .ZN(prince_inst_sbox_inst11_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst11_yyyx_inst_U1 ( .A1(prince_inst_sin_y[44]), 
        .A2(prince_inst_sin_x[47]), .ZN(prince_inst_sbox_inst11_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst11_mux_s00_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[0]), .B(prince_inst_sbox_inst11_s0_sh[0]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh0_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s01_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[1]), .B(prince_inst_sbox_inst11_s0_sh[1]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh0_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s02_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[2]), .B(prince_inst_sbox_inst11_s0_sh[2]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh0_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s03_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[3]), .B(prince_inst_sbox_inst11_s0_sh[3]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh0_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s04_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[4]), .B(prince_inst_sbox_inst11_s0_sh[4]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh0_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s05_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[5]), .B(prince_inst_sbox_inst11_s0_sh[5]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh0_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s06_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[6]), .B(prince_inst_sbox_inst11_s0_sh[6]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh0_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s07_U1 ( .A(
        prince_inst_sbox_inst11_t0_sh[7]), .B(prince_inst_sbox_inst11_s0_sh[7]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh0_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s10_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[0]), .B(prince_inst_sbox_inst11_s1_sh[0]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh1_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s11_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[1]), .B(prince_inst_sbox_inst11_s1_sh[1]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh1_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s12_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[2]), .B(prince_inst_sbox_inst11_s1_sh[2]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh1_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s13_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[3]), .B(prince_inst_sbox_inst11_s1_sh[3]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh1_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s14_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[4]), .B(prince_inst_sbox_inst11_s1_sh[4]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh1_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s15_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[5]), .B(prince_inst_sbox_inst11_s1_sh[5]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh1_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s16_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[6]), .B(prince_inst_sbox_inst11_s1_sh[6]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh1_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s17_U1 ( .A(
        prince_inst_sbox_inst11_t1_sh[7]), .B(prince_inst_sbox_inst11_s1_sh[7]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh1_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s20_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[0]), .B(prince_inst_sbox_inst11_s2_sh[0]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh2_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s21_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[1]), .B(prince_inst_sbox_inst11_s2_sh[1]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh2_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s22_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[2]), .B(prince_inst_sbox_inst11_s2_sh[2]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh2_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s23_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[3]), .B(prince_inst_sbox_inst11_s2_sh[3]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh2_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s24_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[4]), .B(prince_inst_sbox_inst11_s2_sh[4]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh2_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s25_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[5]), .B(prince_inst_sbox_inst11_s2_sh[5]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh2_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s26_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[6]), .B(prince_inst_sbox_inst11_s2_sh[6]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh2_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s27_U1 ( .A(
        prince_inst_sbox_inst11_t2_sh[7]), .B(prince_inst_sbox_inst11_s2_sh[7]), .S(prince_inst_sbox_inst11_n9), .Z(prince_inst_sbox_inst11_sh2_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s30_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[0]), .B(prince_inst_sbox_inst11_s3_sh[0]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s31_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[1]), .B(prince_inst_sbox_inst11_s3_sh[1]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s32_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[2]), .B(prince_inst_sbox_inst11_s3_sh[2]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s33_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[3]), .B(prince_inst_sbox_inst11_s3_sh[3]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s34_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[4]), .B(prince_inst_sbox_inst11_s3_sh[4]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s35_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[5]), .B(prince_inst_sbox_inst11_s3_sh[5]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s36_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[6]), .B(prince_inst_sbox_inst11_s3_sh[6]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst11_mux_s37_U1 ( .A(
        prince_inst_sbox_inst11_t3_sh[7]), .B(prince_inst_sbox_inst11_s3_sh[7]), .S(prince_inst_sbox_inst11_n10), .Z(prince_inst_sbox_inst11_sh3_tmp[7]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk0_U1 ( .A(r[112]), .B(
        prince_inst_sbox_inst11_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[0]), .ZN(prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk1_U1 ( .A(r[113]), .B(
        prince_inst_sbox_inst11_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[1]), .ZN(prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk2_U1 ( .A(r[114]), .B(
        prince_inst_sbox_inst11_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[2]), .ZN(prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk3_U1 ( .A(r[115]), .B(
        prince_inst_sbox_inst11_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[3]), .ZN(prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk4_U1 ( .A(r[112]), .B(
        prince_inst_sbox_inst11_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[4]), .ZN(prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk5_U1 ( .A(r[113]), .B(
        prince_inst_sbox_inst11_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[5]), .ZN(prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk6_U1 ( .A(r[114]), .B(
        prince_inst_sbox_inst11_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[6]), .ZN(prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_msk7_U1 ( .A(r[115]), .B(
        prince_inst_sbox_inst11_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst11_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst0_y[7]), .ZN(prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst11_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst11_c_inst0_ax_n5), .ZN(prince_inst_sout_x[44]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst11_c_inst0_y[1]), .B(
        prince_inst_sbox_inst11_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst11_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst11_c_inst0_y[2]), .B(
        prince_inst_sbox_inst11_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst11_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst11_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst11_c_inst0_ay_n5), .ZN(final_y[44]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst11_c_inst0_y[5]), .B(
        prince_inst_sbox_inst11_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst11_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst11_c_inst0_y[6]), .B(
        prince_inst_sbox_inst11_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst11_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk0_U1 ( .A(r[116]), .B(
        prince_inst_sbox_inst11_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[0]), .ZN(prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk1_U1 ( .A(r[117]), .B(
        prince_inst_sbox_inst11_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[1]), .ZN(prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk2_U1 ( .A(r[118]), .B(
        prince_inst_sbox_inst11_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[2]), .ZN(prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk3_U1 ( .A(r[119]), .B(
        prince_inst_sbox_inst11_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[3]), .ZN(prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk4_U1 ( .A(r[116]), .B(
        prince_inst_sbox_inst11_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[4]), .ZN(prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk5_U1 ( .A(r[117]), .B(
        prince_inst_sbox_inst11_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[5]), .ZN(prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk6_U1 ( .A(r[118]), .B(
        prince_inst_sbox_inst11_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[6]), .ZN(prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_msk7_U1 ( .A(r[119]), .B(
        prince_inst_sbox_inst11_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst11_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst1_y[7]), .ZN(prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst11_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst11_c_inst1_ax_n5), .ZN(prince_inst_sout_x[45]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst11_c_inst1_y[1]), .B(
        prince_inst_sbox_inst11_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst11_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst11_c_inst1_y[2]), .B(
        prince_inst_sbox_inst11_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst11_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst11_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst11_c_inst1_ay_n5), .ZN(final_y[45]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst11_c_inst1_y[5]), .B(
        prince_inst_sbox_inst11_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst11_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst11_c_inst1_y[6]), .B(
        prince_inst_sbox_inst11_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst11_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk0_U1 ( .A(r[120]), .B(
        prince_inst_sbox_inst11_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[0]), .ZN(prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk1_U1 ( .A(r[121]), .B(
        prince_inst_sbox_inst11_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[1]), .ZN(prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk2_U1 ( .A(r[122]), .B(
        prince_inst_sbox_inst11_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[2]), .ZN(prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk3_U1 ( .A(r[123]), .B(
        prince_inst_sbox_inst11_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[3]), .ZN(prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk4_U1 ( .A(r[120]), .B(
        prince_inst_sbox_inst11_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[4]), .ZN(prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk5_U1 ( .A(r[121]), .B(
        prince_inst_sbox_inst11_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[5]), .ZN(prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk6_U1 ( .A(r[122]), .B(
        prince_inst_sbox_inst11_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[6]), .ZN(prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_msk7_U1 ( .A(r[123]), .B(
        prince_inst_sbox_inst11_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst11_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst2_y[7]), .ZN(prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst11_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst11_c_inst2_ax_n5), .ZN(prince_inst_sout_x[46]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst11_c_inst2_y[1]), .B(
        prince_inst_sbox_inst11_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst11_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst11_c_inst2_y[2]), .B(
        prince_inst_sbox_inst11_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst11_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst11_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst11_c_inst2_ay_n5), .ZN(final_y[46]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst11_c_inst2_y[5]), .B(
        prince_inst_sbox_inst11_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst11_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst11_c_inst2_y[6]), .B(
        prince_inst_sbox_inst11_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst11_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk0_U1 ( .A(r[124]), .B(
        prince_inst_sbox_inst11_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[0]), .ZN(prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk1_U1 ( .A(r[125]), .B(
        prince_inst_sbox_inst11_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[1]), .ZN(prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk2_U1 ( .A(r[126]), .B(
        prince_inst_sbox_inst11_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[2]), .ZN(prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk3_U1 ( .A(r[127]), .B(
        prince_inst_sbox_inst11_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[3]), .ZN(prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk4_U1 ( .A(r[124]), .B(
        prince_inst_sbox_inst11_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[4]), .ZN(prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk5_U1 ( .A(r[125]), .B(
        prince_inst_sbox_inst11_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[5]), .ZN(prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk6_U1 ( .A(r[126]), .B(
        prince_inst_sbox_inst11_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[6]), .ZN(prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_msk7_U1 ( .A(r[127]), .B(
        prince_inst_sbox_inst11_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst11_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst11_n7), .A3(
        prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst11_n12), .A2(prince_inst_sbox_inst11_c_inst3_y[7]), .ZN(prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst11_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst11_n12), .ZN(
        prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst11_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst11_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst11_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst11_c_inst3_ax_n5), .ZN(prince_inst_sout_x[47]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst11_c_inst3_y[1]), .B(
        prince_inst_sbox_inst11_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst11_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst11_c_inst3_y[2]), .B(
        prince_inst_sbox_inst11_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst11_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst11_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst11_c_inst3_ay_n5), .ZN(final_y[47]) );
  XNOR2_X1 prince_inst_sbox_inst11_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst11_c_inst3_y[5]), .B(
        prince_inst_sbox_inst11_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst11_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst11_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst11_c_inst3_y[6]), .B(
        prince_inst_sbox_inst11_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst11_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst12_U7 ( .A(prince_inst_sbox_inst12_n13), .ZN(
        prince_inst_sbox_inst12_n12) );
  INV_X1 prince_inst_sbox_inst12_U6 ( .A(prince_inst_n33), .ZN(
        prince_inst_sbox_inst12_n11) );
  INV_X1 prince_inst_sbox_inst12_U5 ( .A(prince_inst_sbox_inst12_n11), .ZN(
        prince_inst_sbox_inst12_n9) );
  INV_X1 prince_inst_sbox_inst12_U4 ( .A(prince_inst_sbox_inst12_n11), .ZN(
        prince_inst_sbox_inst12_n10) );
  INV_X1 prince_inst_sbox_inst12_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst12_n13) );
  INV_X1 prince_inst_sbox_inst12_U2 ( .A(rst), .ZN(prince_inst_sbox_inst12_n8)
         );
  INV_X2 prince_inst_sbox_inst12_U1 ( .A(prince_inst_sbox_inst12_n8), .ZN(
        prince_inst_sbox_inst12_n7) );
  NAND3_X1 prince_inst_sbox_inst12_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n68), .A3(prince_inst_sin_x[48]), 
        .ZN(prince_inst_sbox_inst12_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst12_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U25 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sbox_inst12_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst12_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst12_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst12_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst12_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst12_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n67), .A2(prince_inst_sin_x[50]), 
        .A3(prince_inst_sin_x[48]), .A4(prince_inst_sin_y[51]), .ZN(
        prince_inst_sbox_inst12_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst12_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n61), .A2(prince_inst_sin_x[49]), 
        .A3(prince_inst_sin_x[50]), .ZN(prince_inst_sbox_inst12_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst12_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n66), .A3(prince_inst_sin_x[49]), 
        .A4(prince_inst_sin_x[48]), .ZN(prince_inst_sbox_inst12_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst12_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst12_xxxy_inst_n59), .B(prince_inst_sin_y[51]), .Z(
        prince_inst_sbox_inst12_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst12_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U18 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sin_x[49]), .ZN(prince_inst_sbox_inst12_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst12_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst12_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n65), .A2(prince_inst_sin_x[50]), 
        .ZN(prince_inst_sbox_inst12_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst12_xxxy_inst_U15 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sin_y[51]), .A3(prince_inst_sbox_inst12_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst12_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst12_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst12_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst12_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst12_xxxy_inst_U13 ( .A(prince_inst_sin_x[48]), 
        .B(prince_inst_sin_x[49]), .S(prince_inst_sbox_inst12_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst12_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst12_xxxy_inst_U12 ( .A(prince_inst_sin_y[51]), 
        .ZN(prince_inst_sbox_inst12_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U11 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sin_x[48]), .ZN(prince_inst_sbox_inst12_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst12_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst12_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst12_xxxy_inst_n60), .B(
        prince_inst_sbox_inst12_xxxy_inst_n53), .S(
        prince_inst_sbox_inst12_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst12_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U8 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sbox_inst12_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst12_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U7 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sin_y[51]), .ZN(prince_inst_sbox_inst12_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst12_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst12_t1_sh[0]), .ZN(
        prince_inst_sbox_inst12_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst12_xxxy_inst_U5 ( .A(prince_inst_sin_x[50]), 
        .ZN(prince_inst_sbox_inst12_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U4 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sbox_inst12_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst12_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst12_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst12_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst12_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst12_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst12_xxxy_inst_U2 ( .A(prince_inst_sin_x[48]), 
        .ZN(prince_inst_sbox_inst12_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst12_xxxy_inst_U1 ( .A(prince_inst_sin_x[49]), 
        .ZN(prince_inst_sbox_inst12_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst12_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst12_t1_sh[1]), .B(
        prince_inst_sbox_inst12_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst12_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst12_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst12_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst12_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst12_xxyx_inst_n52), .B(
        prince_inst_sbox_inst12_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst12_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U23 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst12_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst12_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n48), .A2(prince_inst_sin_x[51]), 
        .A3(prince_inst_sin_x[48]), .ZN(prince_inst_sbox_inst12_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst12_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n45), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst12_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst12_xxyx_inst_U18 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n46), .A2(prince_inst_sin_x[51]), 
        .A3(prince_inst_sin_x[49]), .ZN(prince_inst_sbox_inst12_xxyx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst12_t2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst12_xxyx_inst_U16 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sin_x[48]), .A3(prince_inst_sbox_inst12_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst12_xxyx_inst_n44) );
  OR2_X1 prince_inst_sbox_inst12_xxyx_inst_U15 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sbox_inst12_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst12_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst12_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst12_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst12_xxyx_inst_n54), .B(
        prince_inst_sbox_inst12_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst12_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U12 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sin_y[50]), .ZN(prince_inst_sbox_inst12_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst12_xxyx_inst_U11 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sbox_inst12_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst12_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst12_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst12_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst12_xxyx_inst_U10 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst12_xxyx_inst_U9 ( .A1(prince_inst_sin_x[51]), 
        .A2(prince_inst_sbox_inst12_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst12_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst12_xxyx_inst_U8 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sbox_inst12_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst12_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst12_xxyx_inst_U7 ( .A(prince_inst_sin_y[50]), 
        .ZN(prince_inst_sbox_inst12_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst12_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst12_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst12_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n53), .A2(prince_inst_sin_x[49]), 
        .A3(prince_inst_sin_y[50]), .A4(prince_inst_sin_x[48]), .ZN(
        prince_inst_sbox_inst12_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst12_xxyx_inst_U4 ( .A(prince_inst_sin_x[51]), 
        .ZN(prince_inst_sbox_inst12_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst12_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst12_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst12_xxyx_inst_n43), .A3(prince_inst_sin_x[51]), 
        .A4(prince_inst_sin_y[50]), .ZN(prince_inst_sbox_inst12_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst12_xxyx_inst_U2 ( .A(prince_inst_sin_x[48]), 
        .ZN(prince_inst_sbox_inst12_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst12_xxyx_inst_U1 ( .A(prince_inst_sin_x[49]), 
        .ZN(prince_inst_sbox_inst12_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst12_xyxx_inst_n74), .B(
        prince_inst_sbox_inst12_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst12_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst12_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst12_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst12_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U26 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sbox_inst12_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U25 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst12_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst12_xyxx_inst_n72), .B(
        prince_inst_sbox_inst12_s0_sh[2]), .S(
        prince_inst_sbox_inst12_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst12_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst12_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n74), .A2(prince_inst_sin_x[51]), 
        .ZN(prince_inst_sbox_inst12_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst12_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U21 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sbox_inst12_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst12_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst12_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst12_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst12_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst12_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst12_xyxx_inst_U15 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_x[48]), .ZN(prince_inst_sbox_inst12_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst12_xyxx_inst_U13 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U12 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_x[50]), .ZN(prince_inst_sbox_inst12_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst12_xyxx_inst_n58), .B(
        prince_inst_sbox_inst12_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst12_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst12_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst12_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst12_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst12_xyxx_inst_U9 ( .A(prince_inst_sin_x[51]), 
        .ZN(prince_inst_sbox_inst12_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst12_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n54), .A2(prince_inst_sin_x[48]), 
        .ZN(prince_inst_sbox_inst12_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst12_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst12_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst12_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst12_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst12_xyxx_inst_U5 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sbox_inst12_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst12_xyxx_inst_U4 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst12_xyxx_inst_U3 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sbox_inst12_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst12_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst12_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst12_xyxx_inst_U2 ( .A(prince_inst_sin_y[49]), 
        .ZN(prince_inst_sbox_inst12_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst12_xyxx_inst_U1 ( .A(prince_inst_sin_x[50]), 
        .ZN(prince_inst_sbox_inst12_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst12_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst12_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst12_xyyy_inst_n59), .B(
        prince_inst_sbox_inst12_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst12_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst12_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst12_xyyy_inst_U25 ( .A1(prince_inst_sin_y[50]), 
        .A2(prince_inst_sin_y[51]), .A3(prince_inst_sbox_inst12_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst12_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U24 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sbox_inst12_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U23 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sbox_inst12_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst12_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst12_xyyy_inst_U19 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sin_y[50]), .A3(prince_inst_sbox_inst12_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst12_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst12_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst12_xyyy_inst_n49), .B(
        prince_inst_sbox_inst12_xyyy_inst_n48), .S(
        prince_inst_sbox_inst12_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst12_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst12_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst12_xyyy_inst_U16 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sbox_inst12_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst12_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst12_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst12_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst12_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst12_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst12_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst12_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst12_xyyy_inst_U12 ( .A(prince_inst_sin_y[51]), 
        .ZN(prince_inst_sbox_inst12_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst12_xyyy_inst_U11 ( .A1(prince_inst_sin_y[51]), 
        .A2(prince_inst_sbox_inst12_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst12_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst12_t1_sh[3]), .B(
        prince_inst_sbox_inst12_xyyy_inst_n48), .S(
        prince_inst_sbox_inst12_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst12_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst12_xyyy_inst_U9 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sbox_inst12_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst12_xyyy_inst_U8 ( .A1(prince_inst_sin_x[48]), 
        .A2(prince_inst_sin_y[51]), .ZN(prince_inst_sbox_inst12_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst12_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst12_t1_sh[3]), .ZN(
        prince_inst_sbox_inst12_s1_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst12_xyyy_inst_U6 ( .A1(prince_inst_sin_y[51]), 
        .A2(prince_inst_sbox_inst12_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst12_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst12_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst12_xyyy_inst_U4 ( .A(prince_inst_sin_y[49]), 
        .ZN(prince_inst_sbox_inst12_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst12_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst12_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst12_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst12_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst12_xyyy_inst_U2 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_x[48]), .ZN(prince_inst_sbox_inst12_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst12_xyyy_inst_U1 ( .A(prince_inst_sin_y[50]), 
        .ZN(prince_inst_sbox_inst12_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst12_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U27 ( .A1(prince_inst_sin_y[48]), 
        .A2(prince_inst_sbox_inst12_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst12_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U24 ( .A1(prince_inst_sin_y[48]), 
        .A2(prince_inst_sbox_inst12_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst12_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U21 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst12_yxxx_inst_U19 ( .A(prince_inst_sin_x[51]), 
        .ZN(prince_inst_sbox_inst12_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst12_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst12_yxxx_inst_n52), .B(
        prince_inst_sbox_inst12_yxxx_inst_n51), .S(
        prince_inst_sbox_inst12_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst12_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n53), .A2(prince_inst_sin_x[51]), 
        .ZN(prince_inst_sbox_inst12_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst12_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n48), .A2(prince_inst_sin_y[48]), 
        .ZN(prince_inst_sbox_inst12_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n47), .A2(prince_inst_sin_x[51]), 
        .ZN(prince_inst_sbox_inst12_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U13 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sbox_inst12_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst12_yxxx_inst_n59), .B(
        prince_inst_sbox_inst12_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst12_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst12_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst12_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst12_yxxx_inst_U9 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sbox_inst12_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst12_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst12_yxxx_inst_U8 ( .A(
        prince_inst_sbox_inst12_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n51) );
  OR2_X1 prince_inst_sbox_inst12_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst12_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst12_yxxx_inst_U6 ( .A1(prince_inst_sin_x[49]), 
        .A2(prince_inst_sbox_inst12_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst12_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst12_yxxx_inst_U5 ( .A(prince_inst_sin_x[50]), 
        .ZN(prince_inst_sbox_inst12_yxxx_inst_n55) );
  INV_X1 prince_inst_sbox_inst12_yxxx_inst_U4 ( .A(prince_inst_sin_y[48]), 
        .ZN(prince_inst_sbox_inst12_yxxx_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst12_yxxx_inst_U3 ( .A1(
        prince_inst_sbox_inst12_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst12_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst12_yxxx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst12_yxxx_inst_U2 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_yxxx_inst_n45)
         );
  INV_X1 prince_inst_sbox_inst12_yxxx_inst_U1 ( .A(prince_inst_sin_x[49]), 
        .ZN(prince_inst_sbox_inst12_yxxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst12_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst12_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst12_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst12_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst12_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n64), .A3(prince_inst_sin_y[51]), 
        .ZN(prince_inst_sbox_inst12_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst12_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n63), .A2(prince_inst_sin_y[50]), 
        .A3(prince_inst_sin_y[51]), .ZN(prince_inst_sbox_inst12_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst12_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst12_yxyy_inst_n62), .B(
        prince_inst_sbox_inst12_yxyy_inst_n61), .S(prince_inst_sin_y[48]), .Z(
        prince_inst_sbox_inst12_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst12_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst12_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst12_yxyy_inst_n64), .B(
        prince_inst_sbox_inst12_yxyy_inst_n60), .S(
        prince_inst_sbox_inst12_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst12_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst12_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst12_yxyy_inst_n62), .B(
        prince_inst_sbox_inst12_yxyy_inst_n54), .S(
        prince_inst_sbox_inst12_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst12_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst12_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst12_yxyy_inst_n53), .B(
        prince_inst_sbox_inst12_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst12_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst12_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst12_yxyy_inst_n68), .B(
        prince_inst_sbox_inst12_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst12_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U15 ( .A1(prince_inst_sin_y[51]), 
        .A2(prince_inst_sin_y[48]), .ZN(prince_inst_sbox_inst12_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst12_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst12_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst12_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst12_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst12_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst12_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst12_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst12_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n64), .A2(prince_inst_sin_y[50]), 
        .A3(prince_inst_sin_y[48]), .ZN(prince_inst_sbox_inst12_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst12_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U9 ( .A1(prince_inst_sin_y[51]), 
        .A2(prince_inst_sbox_inst12_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst12_yxyy_inst_U8 ( .A1(prince_inst_sin_y[50]), 
        .A2(prince_inst_sbox_inst12_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst12_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst12_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst12_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst12_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst12_yxyy_inst_U5 ( .A(prince_inst_sin_y[48]), 
        .ZN(prince_inst_sbox_inst12_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst12_yxyy_inst_U4 ( .A(prince_inst_sin_x[49]), 
        .ZN(prince_inst_sbox_inst12_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst12_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst12_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst12_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst12_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst12_yxyy_inst_U2 ( .A(prince_inst_sin_y[51]), 
        .ZN(prince_inst_sbox_inst12_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst12_yxyy_inst_U1 ( .A(prince_inst_sin_y[50]), 
        .ZN(prince_inst_sbox_inst12_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst12_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U29 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sbox_inst12_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst12_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst12_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst12_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n75), .A2(prince_inst_sin_y[51]), 
        .A3(prince_inst_sbox_inst12_yyxy_inst_n70), .A4(prince_inst_sin_x[50]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst12_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n69), .A3(prince_inst_sin_y[49]), 
        .A4(prince_inst_sbox_inst12_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst12_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst12_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst12_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst12_yyxy_inst_U23 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_x[50]), .A3(prince_inst_sin_y[48]), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst12_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n69), .A2(prince_inst_sin_y[49]), 
        .A3(prince_inst_sin_y[51]), .ZN(prince_inst_sbox_inst12_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst12_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n75), .A2(prince_inst_sin_x[50]), 
        .A3(prince_inst_sin_y[51]), .ZN(prince_inst_sbox_inst12_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst12_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst12_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst12_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n61), .A2(prince_inst_sin_x[50]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst12_yyxy_inst_U18 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_y[51]), .A3(prince_inst_sbox_inst12_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst12_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst12_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst12_yyxy_inst_U16 ( .A1(prince_inst_sin_y[51]), 
        .A2(prince_inst_sbox_inst12_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst12_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst12_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst12_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n58), .A3(prince_inst_sin_y[48]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst12_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst12_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst12_yyxy_inst_U13 ( .A1(prince_inst_sin_y[48]), 
        .A2(prince_inst_sbox_inst12_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst12_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst12_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst12_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst12_yyxy_inst_n54), .B(
        prince_inst_sbox_inst12_yyxy_inst_n55), .S(
        prince_inst_sbox_inst12_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst12_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst12_yyxy_inst_U9 ( .A(prince_inst_sin_x[50]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n75), .A2(prince_inst_sin_y[51]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst12_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst12_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst12_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U5 ( .A1(prince_inst_sin_x[50]), 
        .A2(prince_inst_sbox_inst12_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst12_yyxy_inst_U4 ( .A(prince_inst_sin_y[49]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst12_yyxy_inst_U3 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sbox_inst12_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst12_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst12_yyxy_inst_U2 ( .A(prince_inst_sin_y[48]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst12_yyxy_inst_U1 ( .A(prince_inst_sin_y[51]), 
        .ZN(prince_inst_sbox_inst12_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst12_yyyx_inst_n58), .B(
        prince_inst_sbox_inst12_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst12_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst12_yyyx_inst_n56), .B(
        prince_inst_sbox_inst12_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst12_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst12_yyyx_inst_n54), .B(
        prince_inst_sbox_inst12_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst12_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst12_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst12_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst12_yyyx_inst_U21 ( .A1(prince_inst_sin_x[51]), 
        .A2(prince_inst_sbox_inst12_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst12_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst12_yyyx_inst_U20 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_y[50]), .A3(prince_inst_sbox_inst12_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst12_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst12_yyyx_inst_n50), .B(
        prince_inst_sbox_inst12_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst12_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst12_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n56), .A2(prince_inst_sin_y[50]), 
        .ZN(prince_inst_sbox_inst12_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst12_yyyx_inst_U17 ( .A1(prince_inst_sin_y[49]), 
        .A2(prince_inst_sin_y[48]), .A3(prince_inst_sin_y[50]), .ZN(
        prince_inst_sbox_inst12_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst12_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst12_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst12_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst12_yyyx_inst_U15 ( .A1(prince_inst_sin_x[51]), 
        .A2(prince_inst_sin_y[50]), .A3(prince_inst_sbox_inst12_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst12_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst12_yyyx_inst_U14 ( .A(prince_inst_sin_y[48]), 
        .ZN(prince_inst_sbox_inst12_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n58), .A2(prince_inst_sin_y[49]), 
        .ZN(prince_inst_sbox_inst12_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst12_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst12_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U11 ( .A1(prince_inst_sin_y[48]), 
        .A2(prince_inst_sbox_inst12_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst12_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst12_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst12_yyyx_inst_U9 ( .A1(prince_inst_sin_y[48]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst12_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst12_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst12_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst12_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n45), .A2(prince_inst_sin_y[48]), 
        .A3(prince_inst_sin_y[50]), .ZN(prince_inst_sbox_inst12_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst12_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst12_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst12_yyyx_inst_U4 ( .A1(prince_inst_sin_x[51]), 
        .A2(prince_inst_sin_y[50]), .ZN(prince_inst_sbox_inst12_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst12_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst12_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst12_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst12_yyyx_inst_U2 ( .A(prince_inst_sin_y[49]), 
        .ZN(prince_inst_sbox_inst12_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst12_yyyx_inst_U1 ( .A1(prince_inst_sin_y[48]), 
        .A2(prince_inst_sin_x[51]), .ZN(prince_inst_sbox_inst12_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst12_mux_s00_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[0]), .B(prince_inst_sbox_inst12_s0_sh[0]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh0_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s01_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[1]), .B(prince_inst_sbox_inst12_s0_sh[1]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh0_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s02_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[2]), .B(prince_inst_sbox_inst12_s0_sh[2]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh0_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s03_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[3]), .B(prince_inst_sbox_inst12_s0_sh[3]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh0_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s04_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[4]), .B(prince_inst_sbox_inst12_s0_sh[4]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh0_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s05_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[5]), .B(prince_inst_sbox_inst12_s0_sh[5]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh0_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s06_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[6]), .B(prince_inst_sbox_inst12_s0_sh[6]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh0_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s07_U1 ( .A(
        prince_inst_sbox_inst12_t0_sh[7]), .B(prince_inst_sbox_inst12_s0_sh[7]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh0_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s10_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[0]), .B(prince_inst_sbox_inst12_s1_sh[0]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh1_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s11_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[1]), .B(prince_inst_sbox_inst12_s1_sh[1]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh1_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s12_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[2]), .B(prince_inst_sbox_inst12_s1_sh[2]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh1_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s13_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[3]), .B(prince_inst_sbox_inst12_s1_sh[3]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh1_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s14_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[4]), .B(prince_inst_sbox_inst12_s1_sh[4]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh1_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s15_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[5]), .B(prince_inst_sbox_inst12_s1_sh[5]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh1_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s16_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[6]), .B(prince_inst_sbox_inst12_s1_sh[6]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh1_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s17_U1 ( .A(
        prince_inst_sbox_inst12_t1_sh[7]), .B(prince_inst_sbox_inst12_s1_sh[7]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh1_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s20_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[0]), .B(prince_inst_sbox_inst12_s2_sh[0]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh2_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s21_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[1]), .B(prince_inst_sbox_inst12_s2_sh[1]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh2_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s22_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[2]), .B(prince_inst_sbox_inst12_s2_sh[2]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh2_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s23_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[3]), .B(prince_inst_sbox_inst12_s2_sh[3]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh2_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s24_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[4]), .B(prince_inst_sbox_inst12_s2_sh[4]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh2_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s25_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[5]), .B(prince_inst_sbox_inst12_s2_sh[5]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh2_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s26_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[6]), .B(prince_inst_sbox_inst12_s2_sh[6]), .S(prince_inst_sbox_inst12_n9), .Z(prince_inst_sbox_inst12_sh2_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s27_U1 ( .A(
        prince_inst_sbox_inst12_t2_sh[7]), .B(prince_inst_sbox_inst12_s2_sh[7]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh2_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s30_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[0]), .B(prince_inst_sbox_inst12_s3_sh[0]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s31_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[1]), .B(prince_inst_sbox_inst12_s3_sh[1]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s32_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[2]), .B(prince_inst_sbox_inst12_s3_sh[2]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s33_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[3]), .B(prince_inst_sbox_inst12_s3_sh[3]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s34_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[4]), .B(prince_inst_sbox_inst12_s3_sh[4]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s35_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[5]), .B(prince_inst_sbox_inst12_s3_sh[5]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s36_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[6]), .B(prince_inst_sbox_inst12_s3_sh[6]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst12_mux_s37_U1 ( .A(
        prince_inst_sbox_inst12_t3_sh[7]), .B(prince_inst_sbox_inst12_s3_sh[7]), .S(prince_inst_sbox_inst12_n10), .Z(prince_inst_sbox_inst12_sh3_tmp[7]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk0_U1 ( .A(r[64]), .B(
        prince_inst_sbox_inst12_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[0]), .ZN(prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk1_U1 ( .A(r[65]), .B(
        prince_inst_sbox_inst12_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[1]), .ZN(prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk2_U1 ( .A(r[66]), .B(
        prince_inst_sbox_inst12_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[2]), .ZN(prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk3_U1 ( .A(r[67]), .B(
        prince_inst_sbox_inst12_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[3]), .ZN(prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk4_U1 ( .A(r[64]), .B(
        prince_inst_sbox_inst12_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[4]), .ZN(prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk5_U1 ( .A(r[65]), .B(
        prince_inst_sbox_inst12_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[5]), .ZN(prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk6_U1 ( .A(r[66]), .B(
        prince_inst_sbox_inst12_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[6]), .ZN(prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_msk7_U1 ( .A(r[67]), .B(
        prince_inst_sbox_inst12_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst12_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst0_y[7]), .ZN(prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst12_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst12_c_inst0_ax_n5), .ZN(prince_inst_sout_x[48]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst12_c_inst0_y[1]), .B(
        prince_inst_sbox_inst12_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst12_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst12_c_inst0_y[2]), .B(
        prince_inst_sbox_inst12_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst12_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst12_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst12_c_inst0_ay_n5), .ZN(final_y[32]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst12_c_inst0_y[5]), .B(
        prince_inst_sbox_inst12_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst12_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst12_c_inst0_y[6]), .B(
        prince_inst_sbox_inst12_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst12_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk0_U1 ( .A(r[68]), .B(
        prince_inst_sbox_inst12_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[0]), .ZN(prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk1_U1 ( .A(r[69]), .B(
        prince_inst_sbox_inst12_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[1]), .ZN(prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk2_U1 ( .A(r[70]), .B(
        prince_inst_sbox_inst12_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[2]), .ZN(prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk3_U1 ( .A(r[71]), .B(
        prince_inst_sbox_inst12_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[3]), .ZN(prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk4_U1 ( .A(r[68]), .B(
        prince_inst_sbox_inst12_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[4]), .ZN(prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk5_U1 ( .A(r[69]), .B(
        prince_inst_sbox_inst12_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[5]), .ZN(prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk6_U1 ( .A(r[70]), .B(
        prince_inst_sbox_inst12_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[6]), .ZN(prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_msk7_U1 ( .A(r[71]), .B(
        prince_inst_sbox_inst12_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst12_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst1_y[7]), .ZN(prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst12_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst12_c_inst1_ax_n5), .ZN(prince_inst_sout_x[49]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst12_c_inst1_y[1]), .B(
        prince_inst_sbox_inst12_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst12_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst12_c_inst1_y[2]), .B(
        prince_inst_sbox_inst12_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst12_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst12_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst12_c_inst1_ay_n5), .ZN(final_y[33]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst12_c_inst1_y[5]), .B(
        prince_inst_sbox_inst12_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst12_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst12_c_inst1_y[6]), .B(
        prince_inst_sbox_inst12_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst12_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk0_U1 ( .A(r[72]), .B(
        prince_inst_sbox_inst12_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[0]), .ZN(prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk1_U1 ( .A(r[73]), .B(
        prince_inst_sbox_inst12_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[1]), .ZN(prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk2_U1 ( .A(r[74]), .B(
        prince_inst_sbox_inst12_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[2]), .ZN(prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk3_U1 ( .A(r[75]), .B(
        prince_inst_sbox_inst12_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[3]), .ZN(prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk4_U1 ( .A(r[72]), .B(
        prince_inst_sbox_inst12_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[4]), .ZN(prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk5_U1 ( .A(r[73]), .B(
        prince_inst_sbox_inst12_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[5]), .ZN(prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk6_U1 ( .A(r[74]), .B(
        prince_inst_sbox_inst12_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[6]), .ZN(prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_msk7_U1 ( .A(r[75]), .B(
        prince_inst_sbox_inst12_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst12_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst2_y[7]), .ZN(prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst12_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst12_c_inst2_ax_n5), .ZN(prince_inst_sout_x[50]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst12_c_inst2_y[1]), .B(
        prince_inst_sbox_inst12_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst12_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst12_c_inst2_y[2]), .B(
        prince_inst_sbox_inst12_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst12_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst12_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst12_c_inst2_ay_n5), .ZN(final_y[34]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst12_c_inst2_y[5]), .B(
        prince_inst_sbox_inst12_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst12_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst12_c_inst2_y[6]), .B(
        prince_inst_sbox_inst12_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst12_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk0_U1 ( .A(r[76]), .B(
        prince_inst_sbox_inst12_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[0]), .ZN(prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk1_U1 ( .A(r[77]), .B(
        prince_inst_sbox_inst12_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[1]), .ZN(prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk2_U1 ( .A(r[78]), .B(
        prince_inst_sbox_inst12_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[2]), .ZN(prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk3_U1 ( .A(r[79]), .B(
        prince_inst_sbox_inst12_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[3]), .ZN(prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk4_U1 ( .A(r[76]), .B(
        prince_inst_sbox_inst12_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[4]), .ZN(prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk5_U1 ( .A(r[77]), .B(
        prince_inst_sbox_inst12_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[5]), .ZN(prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk6_U1 ( .A(r[78]), .B(
        prince_inst_sbox_inst12_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[6]), .ZN(prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_msk7_U1 ( .A(r[79]), .B(
        prince_inst_sbox_inst12_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst12_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst12_n7), .A3(
        prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst12_n12), .A2(prince_inst_sbox_inst12_c_inst3_y[7]), .ZN(prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst12_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst12_n12), .ZN(
        prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst12_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst12_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst12_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst12_c_inst3_ax_n5), .ZN(prince_inst_sout_x[51]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst12_c_inst3_y[1]), .B(
        prince_inst_sbox_inst12_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst12_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst12_c_inst3_y[2]), .B(
        prince_inst_sbox_inst12_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst12_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst12_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst12_c_inst3_ay_n5), .ZN(final_y[35]) );
  XNOR2_X1 prince_inst_sbox_inst12_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst12_c_inst3_y[5]), .B(
        prince_inst_sbox_inst12_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst12_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst12_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst12_c_inst3_y[6]), .B(
        prince_inst_sbox_inst12_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst12_c_inst3_ay_n6) );
  INV_X1 prince_inst_sbox_inst13_U7 ( .A(inv_sig), .ZN(
        prince_inst_sbox_inst13_n11) );
  INV_X4 prince_inst_sbox_inst13_U6 ( .A(prince_inst_sbox_inst13_n13), .ZN(
        prince_inst_sbox_inst13_n12) );
  INV_X1 prince_inst_sbox_inst13_U5 ( .A(prince_inst_sbox_inst13_n11), .ZN(
        prince_inst_sbox_inst13_n10) );
  INV_X1 prince_inst_sbox_inst13_U4 ( .A(prince_inst_sbox_inst13_n11), .ZN(
        prince_inst_sbox_inst13_n9) );
  INV_X1 prince_inst_sbox_inst13_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst13_n13) );
  INV_X1 prince_inst_sbox_inst13_U2 ( .A(rst), .ZN(prince_inst_sbox_inst13_n8)
         );
  INV_X2 prince_inst_sbox_inst13_U1 ( .A(prince_inst_sbox_inst13_n8), .ZN(
        prince_inst_sbox_inst13_n7) );
  NAND3_X1 prince_inst_sbox_inst13_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n68), .A3(prince_inst_sin_x[52]), 
        .ZN(prince_inst_sbox_inst13_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst13_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U25 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sbox_inst13_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst13_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst13_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst13_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst13_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst13_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n67), .A2(prince_inst_sin_x[54]), 
        .A3(prince_inst_sin_x[52]), .A4(prince_inst_sin_y[55]), .ZN(
        prince_inst_sbox_inst13_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst13_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n61), .A2(prince_inst_sin_x[53]), 
        .A3(prince_inst_sin_x[54]), .ZN(prince_inst_sbox_inst13_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst13_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n66), .A3(prince_inst_sin_x[53]), 
        .A4(prince_inst_sin_x[52]), .ZN(prince_inst_sbox_inst13_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst13_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst13_xxxy_inst_n59), .B(prince_inst_sin_y[55]), .Z(
        prince_inst_sbox_inst13_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst13_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U18 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sin_x[53]), .ZN(prince_inst_sbox_inst13_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst13_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst13_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n65), .A2(prince_inst_sin_x[54]), 
        .ZN(prince_inst_sbox_inst13_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst13_xxxy_inst_U15 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sin_y[55]), .A3(prince_inst_sbox_inst13_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst13_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst13_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst13_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst13_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst13_xxxy_inst_U13 ( .A(prince_inst_sin_x[52]), 
        .B(prince_inst_sin_x[53]), .S(prince_inst_sbox_inst13_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst13_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst13_xxxy_inst_U12 ( .A(prince_inst_sin_y[55]), 
        .ZN(prince_inst_sbox_inst13_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U11 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sin_x[52]), .ZN(prince_inst_sbox_inst13_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst13_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst13_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst13_xxxy_inst_n60), .B(
        prince_inst_sbox_inst13_xxxy_inst_n53), .S(
        prince_inst_sbox_inst13_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst13_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U8 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sbox_inst13_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst13_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U7 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sin_y[55]), .ZN(prince_inst_sbox_inst13_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst13_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst13_t1_sh[0]), .ZN(
        prince_inst_sbox_inst13_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst13_xxxy_inst_U5 ( .A(prince_inst_sin_x[54]), 
        .ZN(prince_inst_sbox_inst13_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U4 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sbox_inst13_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst13_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst13_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst13_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst13_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst13_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst13_xxxy_inst_U2 ( .A(prince_inst_sin_x[52]), 
        .ZN(prince_inst_sbox_inst13_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst13_xxxy_inst_U1 ( .A(prince_inst_sin_x[53]), 
        .ZN(prince_inst_sbox_inst13_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst13_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst13_t1_sh[1]), .B(
        prince_inst_sbox_inst13_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst13_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst13_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst13_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst13_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst13_xxyx_inst_n52), .B(
        prince_inst_sbox_inst13_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst13_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U23 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst13_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst13_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n48), .A2(prince_inst_sin_x[55]), 
        .A3(prince_inst_sin_x[52]), .ZN(prince_inst_sbox_inst13_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst13_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst13_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst13_xxyx_inst_U18 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sbox_inst13_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst13_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst13_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst13_xxyx_inst_U16 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sin_x[52]), .A3(prince_inst_sbox_inst13_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst13_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst13_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n46), .A2(prince_inst_sin_x[55]), 
        .A3(prince_inst_sin_x[53]), .ZN(prince_inst_sbox_inst13_xxyx_inst_n44)
         );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst13_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst13_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst13_xxyx_inst_n54), .B(
        prince_inst_sbox_inst13_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst13_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U12 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sin_y[54]), .ZN(prince_inst_sbox_inst13_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst13_xxyx_inst_U11 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sbox_inst13_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst13_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst13_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst13_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst13_xxyx_inst_U10 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst13_xxyx_inst_U9 ( .A1(prince_inst_sin_x[55]), 
        .A2(prince_inst_sbox_inst13_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst13_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst13_xxyx_inst_U8 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sbox_inst13_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst13_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst13_xxyx_inst_U7 ( .A(prince_inst_sin_y[54]), 
        .ZN(prince_inst_sbox_inst13_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst13_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst13_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst13_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n53), .A2(prince_inst_sin_x[53]), 
        .A3(prince_inst_sin_y[54]), .A4(prince_inst_sin_x[52]), .ZN(
        prince_inst_sbox_inst13_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst13_xxyx_inst_U4 ( .A(prince_inst_sin_x[55]), 
        .ZN(prince_inst_sbox_inst13_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst13_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst13_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst13_xxyx_inst_n43), .A3(prince_inst_sin_x[55]), 
        .A4(prince_inst_sin_y[54]), .ZN(prince_inst_sbox_inst13_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst13_xxyx_inst_U2 ( .A(prince_inst_sin_x[52]), 
        .ZN(prince_inst_sbox_inst13_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst13_xxyx_inst_U1 ( .A(prince_inst_sin_x[53]), 
        .ZN(prince_inst_sbox_inst13_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst13_xyxx_inst_n74), .B(
        prince_inst_sbox_inst13_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst13_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst13_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst13_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst13_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U26 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sbox_inst13_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U25 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst13_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst13_xyxx_inst_n72), .B(
        prince_inst_sbox_inst13_s0_sh[2]), .S(
        prince_inst_sbox_inst13_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst13_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst13_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n74), .A2(prince_inst_sin_x[55]), 
        .ZN(prince_inst_sbox_inst13_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst13_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U21 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sbox_inst13_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst13_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst13_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst13_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst13_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst13_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst13_xyxx_inst_U15 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_x[52]), .ZN(prince_inst_sbox_inst13_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst13_xyxx_inst_U13 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U12 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_x[54]), .ZN(prince_inst_sbox_inst13_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst13_xyxx_inst_n58), .B(
        prince_inst_sbox_inst13_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst13_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst13_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst13_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst13_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst13_xyxx_inst_U9 ( .A(prince_inst_sin_x[55]), 
        .ZN(prince_inst_sbox_inst13_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst13_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n54), .A2(prince_inst_sin_x[52]), 
        .ZN(prince_inst_sbox_inst13_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst13_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst13_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst13_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst13_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst13_xyxx_inst_U5 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sbox_inst13_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst13_xyxx_inst_U4 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst13_xyxx_inst_U3 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sbox_inst13_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst13_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst13_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst13_xyxx_inst_U2 ( .A(prince_inst_sin_y[53]), 
        .ZN(prince_inst_sbox_inst13_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst13_xyxx_inst_U1 ( .A(prince_inst_sin_x[54]), 
        .ZN(prince_inst_sbox_inst13_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst13_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst13_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst13_xyyy_inst_n59), .B(
        prince_inst_sbox_inst13_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst13_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst13_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst13_xyyy_inst_U25 ( .A1(prince_inst_sin_y[54]), 
        .A2(prince_inst_sin_y[55]), .A3(prince_inst_sbox_inst13_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst13_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U24 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sbox_inst13_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U23 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sbox_inst13_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst13_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst13_xyyy_inst_U19 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sin_y[54]), .A3(prince_inst_sbox_inst13_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst13_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst13_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst13_xyyy_inst_n49), .B(
        prince_inst_sbox_inst13_xyyy_inst_n48), .S(
        prince_inst_sbox_inst13_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst13_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst13_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst13_xyyy_inst_U16 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sbox_inst13_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst13_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst13_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst13_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst13_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst13_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst13_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst13_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst13_xyyy_inst_U12 ( .A(prince_inst_sin_y[55]), 
        .ZN(prince_inst_sbox_inst13_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst13_xyyy_inst_U11 ( .A1(prince_inst_sin_y[55]), 
        .A2(prince_inst_sbox_inst13_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst13_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst13_t1_sh[3]), .B(
        prince_inst_sbox_inst13_xyyy_inst_n48), .S(
        prince_inst_sbox_inst13_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst13_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst13_xyyy_inst_U9 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sbox_inst13_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst13_xyyy_inst_U8 ( .A1(prince_inst_sin_x[52]), 
        .A2(prince_inst_sin_y[55]), .ZN(prince_inst_sbox_inst13_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst13_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst13_t1_sh[3]), .ZN(
        prince_inst_sbox_inst13_s1_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst13_xyyy_inst_U6 ( .A1(prince_inst_sin_y[55]), 
        .A2(prince_inst_sbox_inst13_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst13_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst13_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst13_xyyy_inst_U4 ( .A(prince_inst_sin_y[53]), 
        .ZN(prince_inst_sbox_inst13_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst13_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst13_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst13_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst13_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst13_xyyy_inst_U2 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_x[52]), .ZN(prince_inst_sbox_inst13_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst13_xyyy_inst_U1 ( .A(prince_inst_sin_y[54]), 
        .ZN(prince_inst_sbox_inst13_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst13_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U27 ( .A1(prince_inst_sin_y[52]), 
        .A2(prince_inst_sbox_inst13_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst13_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U24 ( .A1(prince_inst_sin_y[52]), 
        .A2(prince_inst_sbox_inst13_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst13_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U21 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst13_yxxx_inst_U19 ( .A(prince_inst_sin_x[55]), 
        .ZN(prince_inst_sbox_inst13_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst13_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst13_yxxx_inst_n52), .B(
        prince_inst_sbox_inst13_yxxx_inst_n51), .S(
        prince_inst_sbox_inst13_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst13_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n53), .A2(prince_inst_sin_x[55]), 
        .ZN(prince_inst_sbox_inst13_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst13_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n48), .A2(prince_inst_sin_y[52]), 
        .ZN(prince_inst_sbox_inst13_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n47), .A2(prince_inst_sin_x[55]), 
        .ZN(prince_inst_sbox_inst13_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U13 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sbox_inst13_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst13_yxxx_inst_n59), .B(
        prince_inst_sbox_inst13_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst13_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst13_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst13_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst13_yxxx_inst_U9 ( .A1(prince_inst_sin_x[53]), 
        .A2(prince_inst_sbox_inst13_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst13_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst13_yxxx_inst_U8 ( .A(prince_inst_sin_x[54]), 
        .ZN(prince_inst_sbox_inst13_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst13_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst13_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst13_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst13_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst13_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst13_yxxx_inst_U5 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sbox_inst13_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst13_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst13_yxxx_inst_U4 ( .A(prince_inst_sin_y[52]), 
        .ZN(prince_inst_sbox_inst13_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst13_yxxx_inst_U3 ( .A(prince_inst_sin_x[53]), 
        .ZN(prince_inst_sbox_inst13_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst13_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst13_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst13_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst13_yxxx_inst_U1 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst13_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst13_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst13_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst13_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst13_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n64), .A3(prince_inst_sin_y[55]), 
        .ZN(prince_inst_sbox_inst13_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst13_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n63), .A2(prince_inst_sin_y[54]), 
        .A3(prince_inst_sin_y[55]), .ZN(prince_inst_sbox_inst13_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst13_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst13_yxyy_inst_n62), .B(
        prince_inst_sbox_inst13_yxyy_inst_n61), .S(prince_inst_sin_y[52]), .Z(
        prince_inst_sbox_inst13_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst13_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst13_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst13_yxyy_inst_n64), .B(
        prince_inst_sbox_inst13_yxyy_inst_n60), .S(
        prince_inst_sbox_inst13_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst13_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst13_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst13_yxyy_inst_n62), .B(
        prince_inst_sbox_inst13_yxyy_inst_n54), .S(
        prince_inst_sbox_inst13_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst13_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst13_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst13_yxyy_inst_n53), .B(
        prince_inst_sbox_inst13_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst13_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst13_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst13_yxyy_inst_n68), .B(
        prince_inst_sbox_inst13_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst13_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U15 ( .A1(prince_inst_sin_y[55]), 
        .A2(prince_inst_sin_y[52]), .ZN(prince_inst_sbox_inst13_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst13_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst13_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst13_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst13_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst13_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst13_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst13_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst13_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n64), .A2(prince_inst_sin_y[54]), 
        .A3(prince_inst_sin_y[52]), .ZN(prince_inst_sbox_inst13_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst13_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U9 ( .A1(prince_inst_sin_y[55]), 
        .A2(prince_inst_sbox_inst13_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst13_yxyy_inst_U8 ( .A1(prince_inst_sin_y[54]), 
        .A2(prince_inst_sbox_inst13_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst13_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst13_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst13_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst13_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst13_yxyy_inst_U5 ( .A(prince_inst_sin_y[52]), 
        .ZN(prince_inst_sbox_inst13_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst13_yxyy_inst_U4 ( .A(prince_inst_sin_x[53]), 
        .ZN(prince_inst_sbox_inst13_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst13_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst13_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst13_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst13_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst13_yxyy_inst_U2 ( .A(prince_inst_sin_y[55]), 
        .ZN(prince_inst_sbox_inst13_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst13_yxyy_inst_U1 ( .A(prince_inst_sin_y[54]), 
        .ZN(prince_inst_sbox_inst13_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst13_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U29 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sbox_inst13_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst13_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst13_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst13_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n75), .A2(prince_inst_sin_y[55]), 
        .A3(prince_inst_sbox_inst13_yyxy_inst_n70), .A4(prince_inst_sin_x[54]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst13_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n69), .A3(prince_inst_sin_y[53]), 
        .A4(prince_inst_sbox_inst13_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst13_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst13_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst13_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst13_yyxy_inst_U23 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_x[54]), .A3(prince_inst_sin_y[52]), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst13_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n69), .A2(prince_inst_sin_y[53]), 
        .A3(prince_inst_sin_y[55]), .ZN(prince_inst_sbox_inst13_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst13_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n75), .A2(prince_inst_sin_x[54]), 
        .A3(prince_inst_sin_y[55]), .ZN(prince_inst_sbox_inst13_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst13_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst13_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst13_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n61), .A2(prince_inst_sin_x[54]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst13_yyxy_inst_U18 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_y[55]), .A3(prince_inst_sbox_inst13_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst13_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst13_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst13_yyxy_inst_U16 ( .A1(prince_inst_sin_y[55]), 
        .A2(prince_inst_sbox_inst13_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst13_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst13_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst13_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n58), .A3(prince_inst_sin_y[52]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst13_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst13_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst13_yyxy_inst_U13 ( .A1(prince_inst_sin_y[52]), 
        .A2(prince_inst_sbox_inst13_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst13_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst13_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst13_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst13_yyxy_inst_n54), .B(
        prince_inst_sbox_inst13_yyxy_inst_n55), .S(
        prince_inst_sbox_inst13_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst13_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst13_yyxy_inst_U9 ( .A(prince_inst_sin_x[54]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n75), .A2(prince_inst_sin_y[55]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst13_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst13_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst13_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U5 ( .A1(prince_inst_sin_x[54]), 
        .A2(prince_inst_sbox_inst13_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst13_yyxy_inst_U4 ( .A(prince_inst_sin_y[53]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst13_yyxy_inst_U3 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sbox_inst13_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst13_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst13_yyxy_inst_U2 ( .A(prince_inst_sin_y[52]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst13_yyxy_inst_U1 ( .A(prince_inst_sin_y[55]), 
        .ZN(prince_inst_sbox_inst13_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst13_yyyx_inst_n58), .B(
        prince_inst_sbox_inst13_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst13_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst13_yyyx_inst_n56), .B(
        prince_inst_sbox_inst13_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst13_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst13_yyyx_inst_n54), .B(
        prince_inst_sbox_inst13_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst13_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst13_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst13_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst13_yyyx_inst_U21 ( .A1(prince_inst_sin_x[55]), 
        .A2(prince_inst_sbox_inst13_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst13_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst13_yyyx_inst_U20 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_y[54]), .A3(prince_inst_sbox_inst13_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst13_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst13_yyyx_inst_n50), .B(
        prince_inst_sbox_inst13_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst13_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst13_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n56), .A2(prince_inst_sin_y[54]), 
        .ZN(prince_inst_sbox_inst13_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst13_yyyx_inst_U17 ( .A1(prince_inst_sin_y[53]), 
        .A2(prince_inst_sin_y[52]), .A3(prince_inst_sin_y[54]), .ZN(
        prince_inst_sbox_inst13_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst13_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst13_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst13_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst13_yyyx_inst_U15 ( .A1(prince_inst_sin_x[55]), 
        .A2(prince_inst_sin_y[54]), .A3(prince_inst_sbox_inst13_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst13_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst13_yyyx_inst_U14 ( .A(prince_inst_sin_y[52]), 
        .ZN(prince_inst_sbox_inst13_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n58), .A2(prince_inst_sin_y[53]), 
        .ZN(prince_inst_sbox_inst13_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst13_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst13_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U11 ( .A1(prince_inst_sin_y[52]), 
        .A2(prince_inst_sbox_inst13_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst13_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst13_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst13_yyyx_inst_U9 ( .A1(prince_inst_sin_y[52]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst13_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst13_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst13_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst13_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n45), .A2(prince_inst_sin_y[52]), 
        .A3(prince_inst_sin_y[54]), .ZN(prince_inst_sbox_inst13_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst13_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst13_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst13_yyyx_inst_U4 ( .A1(prince_inst_sin_x[55]), 
        .A2(prince_inst_sin_y[54]), .ZN(prince_inst_sbox_inst13_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst13_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst13_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst13_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst13_yyyx_inst_U2 ( .A(prince_inst_sin_y[53]), 
        .ZN(prince_inst_sbox_inst13_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst13_yyyx_inst_U1 ( .A1(prince_inst_sin_y[52]), 
        .A2(prince_inst_sin_x[55]), .ZN(prince_inst_sbox_inst13_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst13_mux_s00_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[0]), .B(prince_inst_sbox_inst13_s0_sh[0]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh0_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s01_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[1]), .B(prince_inst_sbox_inst13_s0_sh[1]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh0_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s02_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[2]), .B(prince_inst_sbox_inst13_s0_sh[2]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh0_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s03_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[3]), .B(prince_inst_sbox_inst13_s0_sh[3]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh0_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s04_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[4]), .B(prince_inst_sbox_inst13_s0_sh[4]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh0_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s05_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[5]), .B(prince_inst_sbox_inst13_s0_sh[5]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh0_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s06_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[6]), .B(prince_inst_sbox_inst13_s0_sh[6]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh0_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s07_U1 ( .A(
        prince_inst_sbox_inst13_t0_sh[7]), .B(prince_inst_sbox_inst13_s0_sh[7]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh0_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s10_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[0]), .B(prince_inst_sbox_inst13_s1_sh[0]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh1_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s11_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[1]), .B(prince_inst_sbox_inst13_s1_sh[1]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh1_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s12_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[2]), .B(prince_inst_sbox_inst13_s1_sh[2]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh1_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s13_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[3]), .B(prince_inst_sbox_inst13_s1_sh[3]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh1_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s14_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[4]), .B(prince_inst_sbox_inst13_s1_sh[4]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh1_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s15_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[5]), .B(prince_inst_sbox_inst13_s1_sh[5]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh1_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s16_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[6]), .B(prince_inst_sbox_inst13_s1_sh[6]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh1_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s17_U1 ( .A(
        prince_inst_sbox_inst13_t1_sh[7]), .B(prince_inst_sbox_inst13_s1_sh[7]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh1_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s20_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[0]), .B(prince_inst_sbox_inst13_s2_sh[0]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh2_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s21_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[1]), .B(prince_inst_sbox_inst13_s2_sh[1]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh2_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s22_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[2]), .B(prince_inst_sbox_inst13_s2_sh[2]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh2_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s23_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[3]), .B(prince_inst_sbox_inst13_s2_sh[3]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh2_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s24_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[4]), .B(prince_inst_sbox_inst13_s2_sh[4]), .S(inv_sig), .Z(prince_inst_sbox_inst13_sh2_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s25_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[5]), .B(prince_inst_sbox_inst13_s2_sh[5]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh2_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s26_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[6]), .B(prince_inst_sbox_inst13_s2_sh[6]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh2_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s27_U1 ( .A(
        prince_inst_sbox_inst13_t2_sh[7]), .B(prince_inst_sbox_inst13_s2_sh[7]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh2_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s30_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[0]), .B(prince_inst_sbox_inst13_s3_sh[0]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh3_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s31_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[1]), .B(prince_inst_sbox_inst13_s3_sh[1]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh3_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s32_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[2]), .B(prince_inst_sbox_inst13_s3_sh[2]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh3_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s33_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[3]), .B(prince_inst_sbox_inst13_s3_sh[3]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh3_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s34_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[4]), .B(prince_inst_sbox_inst13_s3_sh[4]), .S(prince_inst_sbox_inst13_n9), .Z(prince_inst_sbox_inst13_sh3_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s35_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[5]), .B(prince_inst_sbox_inst13_s3_sh[5]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh3_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s36_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[6]), .B(prince_inst_sbox_inst13_s3_sh[6]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh3_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst13_mux_s37_U1 ( .A(
        prince_inst_sbox_inst13_t3_sh[7]), .B(prince_inst_sbox_inst13_s3_sh[7]), .S(prince_inst_sbox_inst13_n10), .Z(prince_inst_sbox_inst13_sh3_tmp[7]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk0_U1 ( .A(r[80]), .B(
        prince_inst_sbox_inst13_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[0]), .ZN(prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk1_U1 ( .A(r[81]), .B(
        prince_inst_sbox_inst13_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[1]), .ZN(prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk2_U1 ( .A(r[82]), .B(
        prince_inst_sbox_inst13_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[2]), .ZN(prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk3_U1 ( .A(r[83]), .B(
        prince_inst_sbox_inst13_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[3]), .ZN(prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk4_U1 ( .A(r[80]), .B(
        prince_inst_sbox_inst13_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[4]), .ZN(prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk5_U1 ( .A(r[81]), .B(
        prince_inst_sbox_inst13_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[5]), .ZN(prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk6_U1 ( .A(r[82]), .B(
        prince_inst_sbox_inst13_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[6]), .ZN(prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_msk7_U1 ( .A(r[83]), .B(
        prince_inst_sbox_inst13_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst13_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst0_y[7]), .ZN(prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst13_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst13_c_inst0_ax_n5), .ZN(prince_inst_sout_x[52]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst13_c_inst0_y[1]), .B(
        prince_inst_sbox_inst13_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst13_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst13_c_inst0_y[2]), .B(
        prince_inst_sbox_inst13_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst13_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst13_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst13_c_inst0_ay_n5), .ZN(final_y[20]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst13_c_inst0_y[5]), .B(
        prince_inst_sbox_inst13_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst13_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst13_c_inst0_y[6]), .B(
        prince_inst_sbox_inst13_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst13_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk0_U1 ( .A(r[84]), .B(
        prince_inst_sbox_inst13_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[0]), .ZN(prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk1_U1 ( .A(r[85]), .B(
        prince_inst_sbox_inst13_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[1]), .ZN(prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk2_U1 ( .A(r[86]), .B(
        prince_inst_sbox_inst13_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[2]), .ZN(prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk3_U1 ( .A(r[87]), .B(
        prince_inst_sbox_inst13_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[3]), .ZN(prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk4_U1 ( .A(r[84]), .B(
        prince_inst_sbox_inst13_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[4]), .ZN(prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk5_U1 ( .A(r[85]), .B(
        prince_inst_sbox_inst13_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[5]), .ZN(prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk6_U1 ( .A(r[86]), .B(
        prince_inst_sbox_inst13_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[6]), .ZN(prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_msk7_U1 ( .A(r[87]), .B(
        prince_inst_sbox_inst13_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst13_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst1_y[7]), .ZN(prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst13_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst13_c_inst1_ax_n5), .ZN(prince_inst_sout_x[53]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst13_c_inst1_y[1]), .B(
        prince_inst_sbox_inst13_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst13_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst13_c_inst1_y[2]), .B(
        prince_inst_sbox_inst13_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst13_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst13_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst13_c_inst1_ay_n5), .ZN(final_y[21]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst13_c_inst1_y[5]), .B(
        prince_inst_sbox_inst13_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst13_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst13_c_inst1_y[6]), .B(
        prince_inst_sbox_inst13_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst13_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk0_U1 ( .A(r[88]), .B(
        prince_inst_sbox_inst13_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[0]), .ZN(prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk1_U1 ( .A(r[89]), .B(
        prince_inst_sbox_inst13_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[1]), .ZN(prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk2_U1 ( .A(r[90]), .B(
        prince_inst_sbox_inst13_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[2]), .ZN(prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk3_U1 ( .A(r[91]), .B(
        prince_inst_sbox_inst13_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[3]), .ZN(prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk4_U1 ( .A(r[88]), .B(
        prince_inst_sbox_inst13_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[4]), .ZN(prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk5_U1 ( .A(r[89]), .B(
        prince_inst_sbox_inst13_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[5]), .ZN(prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk6_U1 ( .A(r[90]), .B(
        prince_inst_sbox_inst13_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[6]), .ZN(prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_msk7_U1 ( .A(r[91]), .B(
        prince_inst_sbox_inst13_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst13_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst2_y[7]), .ZN(prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst13_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst13_c_inst2_ax_n5), .ZN(prince_inst_sout_x[54]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst13_c_inst2_y[1]), .B(
        prince_inst_sbox_inst13_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst13_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst13_c_inst2_y[2]), .B(
        prince_inst_sbox_inst13_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst13_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst13_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst13_c_inst2_ay_n5), .ZN(final_y[22]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst13_c_inst2_y[5]), .B(
        prince_inst_sbox_inst13_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst13_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst13_c_inst2_y[6]), .B(
        prince_inst_sbox_inst13_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst13_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk0_U1 ( .A(r[92]), .B(
        prince_inst_sbox_inst13_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[0]), .ZN(prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk1_U1 ( .A(r[93]), .B(
        prince_inst_sbox_inst13_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[1]), .ZN(prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk2_U1 ( .A(r[94]), .B(
        prince_inst_sbox_inst13_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[2]), .ZN(prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk3_U1 ( .A(r[95]), .B(
        prince_inst_sbox_inst13_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[3]), .ZN(prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk4_U1 ( .A(r[92]), .B(
        prince_inst_sbox_inst13_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[4]), .ZN(prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk5_U1 ( .A(r[93]), .B(
        prince_inst_sbox_inst13_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[5]), .ZN(prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk6_U1 ( .A(r[94]), .B(
        prince_inst_sbox_inst13_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[6]), .ZN(prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_msk7_U1 ( .A(r[95]), .B(
        prince_inst_sbox_inst13_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst13_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst13_n7), .A3(
        prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst13_n12), .A2(prince_inst_sbox_inst13_c_inst3_y[7]), .ZN(prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst13_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst13_n12), .ZN(
        prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst13_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst13_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst13_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst13_c_inst3_ax_n5), .ZN(prince_inst_sout_x[55]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst13_c_inst3_y[1]), .B(
        prince_inst_sbox_inst13_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst13_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst13_c_inst3_y[2]), .B(
        prince_inst_sbox_inst13_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst13_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst13_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst13_c_inst3_ay_n5), .ZN(final_y[23]) );
  XNOR2_X1 prince_inst_sbox_inst13_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst13_c_inst3_y[5]), .B(
        prince_inst_sbox_inst13_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst13_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst13_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst13_c_inst3_y[6]), .B(
        prince_inst_sbox_inst13_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst13_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst14_U7 ( .A(prince_inst_sbox_inst14_n13), .ZN(
        prince_inst_sbox_inst14_n12) );
  INV_X1 prince_inst_sbox_inst14_U6 ( .A(prince_inst_n33), .ZN(
        prince_inst_sbox_inst14_n11) );
  INV_X1 prince_inst_sbox_inst14_U5 ( .A(prince_inst_sbox_inst14_n11), .ZN(
        prince_inst_sbox_inst14_n9) );
  INV_X1 prince_inst_sbox_inst14_U4 ( .A(prince_inst_sbox_inst14_n11), .ZN(
        prince_inst_sbox_inst14_n10) );
  INV_X1 prince_inst_sbox_inst14_U3 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst14_n13) );
  INV_X1 prince_inst_sbox_inst14_U2 ( .A(rst), .ZN(prince_inst_sbox_inst14_n8)
         );
  INV_X2 prince_inst_sbox_inst14_U1 ( .A(prince_inst_sbox_inst14_n8), .ZN(
        prince_inst_sbox_inst14_n7) );
  NAND3_X1 prince_inst_sbox_inst14_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n68), .A3(prince_inst_sin_x[56]), 
        .ZN(prince_inst_sbox_inst14_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst14_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U25 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sbox_inst14_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst14_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst14_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst14_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst14_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst14_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n67), .A2(prince_inst_sin_x[58]), 
        .A3(prince_inst_sin_x[56]), .A4(prince_inst_sin_y[59]), .ZN(
        prince_inst_sbox_inst14_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst14_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n61), .A2(prince_inst_sin_x[57]), 
        .A3(prince_inst_sin_x[58]), .ZN(prince_inst_sbox_inst14_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst14_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n66), .A3(prince_inst_sin_x[57]), 
        .A4(prince_inst_sin_x[56]), .ZN(prince_inst_sbox_inst14_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst14_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst14_xxxy_inst_n59), .B(prince_inst_sin_y[59]), .Z(
        prince_inst_sbox_inst14_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst14_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U18 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sin_x[57]), .ZN(prince_inst_sbox_inst14_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst14_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst14_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n65), .A2(prince_inst_sin_x[58]), 
        .ZN(prince_inst_sbox_inst14_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst14_xxxy_inst_U15 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sin_y[59]), .A3(prince_inst_sbox_inst14_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst14_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst14_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst14_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst14_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst14_xxxy_inst_U13 ( .A(prince_inst_sin_x[56]), 
        .B(prince_inst_sin_x[57]), .S(prince_inst_sbox_inst14_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst14_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst14_xxxy_inst_U12 ( .A(prince_inst_sin_y[59]), 
        .ZN(prince_inst_sbox_inst14_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U11 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sin_x[56]), .ZN(prince_inst_sbox_inst14_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst14_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst14_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst14_xxxy_inst_n60), .B(
        prince_inst_sbox_inst14_xxxy_inst_n53), .S(
        prince_inst_sbox_inst14_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst14_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U8 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sbox_inst14_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst14_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U7 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sin_y[59]), .ZN(prince_inst_sbox_inst14_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst14_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst14_t1_sh[0]), .ZN(
        prince_inst_sbox_inst14_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst14_xxxy_inst_U5 ( .A(prince_inst_sin_x[58]), 
        .ZN(prince_inst_sbox_inst14_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U4 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sbox_inst14_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst14_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst14_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst14_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst14_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst14_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst14_xxxy_inst_U2 ( .A(prince_inst_sin_x[56]), 
        .ZN(prince_inst_sbox_inst14_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst14_xxxy_inst_U1 ( .A(prince_inst_sin_x[57]), 
        .ZN(prince_inst_sbox_inst14_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst14_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst14_t1_sh[1]), .B(
        prince_inst_sbox_inst14_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst14_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst14_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst14_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst14_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst14_xxyx_inst_n52), .B(
        prince_inst_sbox_inst14_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst14_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U23 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst14_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst14_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n48), .A2(prince_inst_sin_x[59]), 
        .A3(prince_inst_sin_x[56]), .ZN(prince_inst_sbox_inst14_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst14_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst14_t2_sh[1]) );
  OR2_X1 prince_inst_sbox_inst14_xxyx_inst_U18 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sbox_inst14_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst14_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n44), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n45), .ZN(
        prince_inst_sbox_inst14_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst14_xxyx_inst_U16 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sin_x[56]), .A3(prince_inst_sbox_inst14_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst14_xxyx_inst_n45) );
  NAND3_X1 prince_inst_sbox_inst14_xxyx_inst_U15 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n46), .A2(prince_inst_sin_x[59]), 
        .A3(prince_inst_sin_x[57]), .ZN(prince_inst_sbox_inst14_xxyx_inst_n44)
         );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst14_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst14_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst14_xxyx_inst_n54), .B(
        prince_inst_sbox_inst14_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst14_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U12 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sin_y[58]), .ZN(prince_inst_sbox_inst14_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst14_xxyx_inst_U11 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sbox_inst14_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst14_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst14_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst14_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst14_xxyx_inst_U10 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst14_xxyx_inst_U9 ( .A1(prince_inst_sin_x[59]), 
        .A2(prince_inst_sbox_inst14_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst14_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst14_xxyx_inst_U8 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sbox_inst14_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst14_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst14_xxyx_inst_U7 ( .A(prince_inst_sin_y[58]), 
        .ZN(prince_inst_sbox_inst14_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst14_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst14_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst14_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n53), .A2(prince_inst_sin_x[57]), 
        .A3(prince_inst_sin_y[58]), .A4(prince_inst_sin_x[56]), .ZN(
        prince_inst_sbox_inst14_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst14_xxyx_inst_U4 ( .A(prince_inst_sin_x[59]), 
        .ZN(prince_inst_sbox_inst14_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst14_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst14_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst14_xxyx_inst_n43), .A3(prince_inst_sin_x[59]), 
        .A4(prince_inst_sin_y[58]), .ZN(prince_inst_sbox_inst14_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst14_xxyx_inst_U2 ( .A(prince_inst_sin_x[56]), 
        .ZN(prince_inst_sbox_inst14_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst14_xxyx_inst_U1 ( .A(prince_inst_sin_x[57]), 
        .ZN(prince_inst_sbox_inst14_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst14_xyxx_inst_n74), .B(
        prince_inst_sbox_inst14_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst14_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst14_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst14_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst14_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U26 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sbox_inst14_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U25 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst14_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst14_xyxx_inst_n72), .B(
        prince_inst_sbox_inst14_s0_sh[2]), .S(
        prince_inst_sbox_inst14_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst14_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst14_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n74), .A2(prince_inst_sin_x[59]), 
        .ZN(prince_inst_sbox_inst14_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst14_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U21 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sbox_inst14_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst14_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst14_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n74) );
  XNOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U19 ( .A(
        prince_inst_sbox_inst14_xyxx_inst_n61), .B(
        prince_inst_sbox_inst14_xyxx_inst_n60), .ZN(
        prince_inst_sbox_inst14_t1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst14_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U17 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst14_xyxx_inst_U16 ( .A(
        prince_inst_sbox_inst14_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U15 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n58) );
  NAND2_X1 prince_inst_sbox_inst14_xyxx_inst_U14 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_x[56]), .ZN(prince_inst_sbox_inst14_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U13 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst14_xyxx_inst_U12 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_xyxx_inst_n57)
         );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U11 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_x[58]), .ZN(prince_inst_sbox_inst14_xyxx_inst_n70)
         );
  NOR3_X1 prince_inst_sbox_inst14_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst14_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst14_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst14_xyxx_inst_U9 ( .A(prince_inst_sin_x[59]), 
        .ZN(prince_inst_sbox_inst14_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst14_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n54), .A2(prince_inst_sin_x[56]), 
        .ZN(prince_inst_sbox_inst14_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst14_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst14_xyxx_inst_n61), .A2(
        prince_inst_sbox_inst14_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst14_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst14_xyxx_inst_U5 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sbox_inst14_xyxx_inst_n60), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst14_xyxx_inst_U4 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_xyxx_inst_n60)
         );
  NOR3_X1 prince_inst_sbox_inst14_xyxx_inst_U3 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sbox_inst14_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst14_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst14_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst14_xyxx_inst_U2 ( .A(prince_inst_sin_y[57]), 
        .ZN(prince_inst_sbox_inst14_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst14_xyxx_inst_U1 ( .A(prince_inst_sin_x[58]), 
        .ZN(prince_inst_sbox_inst14_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst14_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst14_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst14_xyyy_inst_n59), .B(
        prince_inst_sbox_inst14_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst14_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst14_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst14_xyyy_inst_U25 ( .A1(prince_inst_sin_y[58]), 
        .A2(prince_inst_sin_y[59]), .A3(prince_inst_sbox_inst14_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst14_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U24 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sbox_inst14_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U23 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sbox_inst14_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst14_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst14_xyyy_inst_U19 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sin_y[58]), .A3(prince_inst_sbox_inst14_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst14_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst14_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst14_xyyy_inst_n49), .B(
        prince_inst_sbox_inst14_xyyy_inst_n48), .S(
        prince_inst_sbox_inst14_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst14_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst14_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst14_xyyy_inst_U16 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sbox_inst14_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst14_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst14_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst14_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst14_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst14_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst14_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst14_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst14_xyyy_inst_U12 ( .A(prince_inst_sin_y[59]), 
        .ZN(prince_inst_sbox_inst14_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst14_xyyy_inst_U11 ( .A1(prince_inst_sin_y[59]), 
        .A2(prince_inst_sbox_inst14_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst14_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst14_t1_sh[3]), .B(
        prince_inst_sbox_inst14_xyyy_inst_n48), .S(
        prince_inst_sbox_inst14_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst14_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst14_xyyy_inst_U9 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sbox_inst14_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst14_xyyy_inst_U8 ( .A1(prince_inst_sin_x[56]), 
        .A2(prince_inst_sin_y[59]), .ZN(prince_inst_sbox_inst14_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst14_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst14_t1_sh[3]), .ZN(
        prince_inst_sbox_inst14_s1_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst14_xyyy_inst_U6 ( .A1(prince_inst_sin_y[59]), 
        .A2(prince_inst_sbox_inst14_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst14_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst14_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst14_xyyy_inst_U4 ( .A(prince_inst_sin_y[57]), 
        .ZN(prince_inst_sbox_inst14_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst14_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst14_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst14_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst14_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst14_xyyy_inst_U2 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_x[56]), .ZN(prince_inst_sbox_inst14_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst14_xyyy_inst_U1 ( .A(prince_inst_sin_y[58]), 
        .ZN(prince_inst_sbox_inst14_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst14_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U27 ( .A1(prince_inst_sin_y[56]), 
        .A2(prince_inst_sbox_inst14_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U26 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst14_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U24 ( .A1(prince_inst_sin_y[56]), 
        .A2(prince_inst_sbox_inst14_yxxx_inst_n57), .ZN(
        prince_inst_sbox_inst14_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U23 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n57) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U21 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_yxxx_inst_n54)
         );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n62) );
  INV_X1 prince_inst_sbox_inst14_yxxx_inst_U19 ( .A(prince_inst_sin_x[59]), 
        .ZN(prince_inst_sbox_inst14_yxxx_inst_n58) );
  MUX2_X1 prince_inst_sbox_inst14_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst14_yxxx_inst_n52), .B(
        prince_inst_sbox_inst14_yxxx_inst_n51), .S(
        prince_inst_sbox_inst14_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst14_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n53), .A2(prince_inst_sin_x[59]), 
        .ZN(prince_inst_sbox_inst14_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n61), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst14_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n48), .A2(prince_inst_sin_y[56]), 
        .ZN(prince_inst_sbox_inst14_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n47), .A2(prince_inst_sin_x[59]), 
        .ZN(prince_inst_sbox_inst14_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U13 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sbox_inst14_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n61) );
  XNOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst14_yxxx_inst_n59), .B(
        prince_inst_sbox_inst14_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst14_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst14_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst14_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst14_yxxx_inst_U9 ( .A1(prince_inst_sin_x[57]), 
        .A2(prince_inst_sbox_inst14_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst14_yxxx_inst_n55), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n59) );
  INV_X1 prince_inst_sbox_inst14_yxxx_inst_U8 ( .A(prince_inst_sin_x[58]), 
        .ZN(prince_inst_sbox_inst14_yxxx_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst14_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst14_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst14_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst14_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst14_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst14_yxxx_inst_U5 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sbox_inst14_yxxx_inst_n53), .A3(
        prince_inst_sbox_inst14_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst14_yxxx_inst_U4 ( .A(prince_inst_sin_y[56]), 
        .ZN(prince_inst_sbox_inst14_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst14_yxxx_inst_U3 ( .A(prince_inst_sin_x[57]), 
        .ZN(prince_inst_sbox_inst14_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst14_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst14_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst14_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst14_yxxx_inst_U1 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst14_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst14_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst14_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst14_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst14_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n64), .A3(prince_inst_sin_y[59]), 
        .ZN(prince_inst_sbox_inst14_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst14_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n63), .A2(prince_inst_sin_y[58]), 
        .A3(prince_inst_sin_y[59]), .ZN(prince_inst_sbox_inst14_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst14_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst14_yxyy_inst_n62), .B(
        prince_inst_sbox_inst14_yxyy_inst_n61), .S(prince_inst_sin_y[56]), .Z(
        prince_inst_sbox_inst14_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst14_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst14_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst14_yxyy_inst_n64), .B(
        prince_inst_sbox_inst14_yxyy_inst_n60), .S(
        prince_inst_sbox_inst14_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst14_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst14_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst14_yxyy_inst_n62), .B(
        prince_inst_sbox_inst14_yxyy_inst_n54), .S(
        prince_inst_sbox_inst14_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst14_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst14_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst14_yxyy_inst_n53), .B(
        prince_inst_sbox_inst14_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst14_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst14_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst14_yxyy_inst_n68), .B(
        prince_inst_sbox_inst14_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst14_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U15 ( .A1(prince_inst_sin_y[59]), 
        .A2(prince_inst_sin_y[56]), .ZN(prince_inst_sbox_inst14_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst14_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst14_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst14_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst14_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst14_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst14_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst14_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst14_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n64), .A2(prince_inst_sin_y[58]), 
        .A3(prince_inst_sin_y[56]), .ZN(prince_inst_sbox_inst14_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst14_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U9 ( .A1(prince_inst_sin_y[59]), 
        .A2(prince_inst_sbox_inst14_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst14_yxyy_inst_U8 ( .A1(prince_inst_sin_y[58]), 
        .A2(prince_inst_sbox_inst14_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst14_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst14_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst14_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst14_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst14_yxyy_inst_U5 ( .A(prince_inst_sin_y[56]), 
        .ZN(prince_inst_sbox_inst14_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst14_yxyy_inst_U4 ( .A(prince_inst_sin_x[57]), 
        .ZN(prince_inst_sbox_inst14_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst14_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst14_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst14_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst14_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst14_yxyy_inst_U2 ( .A(prince_inst_sin_y[59]), 
        .ZN(prince_inst_sbox_inst14_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst14_yxyy_inst_U1 ( .A(prince_inst_sin_y[58]), 
        .ZN(prince_inst_sbox_inst14_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst14_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U29 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sbox_inst14_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst14_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst14_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst14_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n75), .A2(prince_inst_sin_y[59]), 
        .A3(prince_inst_sbox_inst14_yyxy_inst_n70), .A4(prince_inst_sin_x[58]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst14_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n69), .A3(prince_inst_sin_y[57]), 
        .A4(prince_inst_sbox_inst14_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst14_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst14_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst14_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst14_yyxy_inst_U23 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_x[58]), .A3(prince_inst_sin_y[56]), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst14_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n69), .A2(prince_inst_sin_y[57]), 
        .A3(prince_inst_sin_y[59]), .ZN(prince_inst_sbox_inst14_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst14_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n75), .A2(prince_inst_sin_x[58]), 
        .A3(prince_inst_sin_y[59]), .ZN(prince_inst_sbox_inst14_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst14_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst14_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst14_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n61), .A2(prince_inst_sin_x[58]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst14_yyxy_inst_U18 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_y[59]), .A3(prince_inst_sbox_inst14_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst14_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst14_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst14_yyxy_inst_U16 ( .A1(prince_inst_sin_y[59]), 
        .A2(prince_inst_sbox_inst14_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst14_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst14_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst14_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n58), .A3(prince_inst_sin_y[56]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst14_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst14_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst14_yyxy_inst_U13 ( .A1(prince_inst_sin_y[56]), 
        .A2(prince_inst_sbox_inst14_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst14_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst14_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst14_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst14_yyxy_inst_n54), .B(
        prince_inst_sbox_inst14_yyxy_inst_n55), .S(
        prince_inst_sbox_inst14_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst14_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst14_yyxy_inst_U9 ( .A(prince_inst_sin_x[58]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n75), .A2(prince_inst_sin_y[59]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst14_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst14_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst14_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U5 ( .A1(prince_inst_sin_x[58]), 
        .A2(prince_inst_sbox_inst14_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst14_yyxy_inst_U4 ( .A(prince_inst_sin_y[57]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst14_yyxy_inst_U3 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sbox_inst14_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst14_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst14_yyxy_inst_U2 ( .A(prince_inst_sin_y[56]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst14_yyxy_inst_U1 ( .A(prince_inst_sin_y[59]), 
        .ZN(prince_inst_sbox_inst14_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst14_yyyx_inst_n58), .B(
        prince_inst_sbox_inst14_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst14_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst14_yyyx_inst_n56), .B(
        prince_inst_sbox_inst14_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst14_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst14_yyyx_inst_n54), .B(
        prince_inst_sbox_inst14_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst14_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst14_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst14_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst14_yyyx_inst_U21 ( .A1(prince_inst_sin_x[59]), 
        .A2(prince_inst_sbox_inst14_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst14_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst14_yyyx_inst_U20 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_y[58]), .A3(prince_inst_sbox_inst14_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst14_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst14_yyyx_inst_n50), .B(
        prince_inst_sbox_inst14_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst14_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst14_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n56), .A2(prince_inst_sin_y[58]), 
        .ZN(prince_inst_sbox_inst14_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst14_yyyx_inst_U17 ( .A1(prince_inst_sin_y[57]), 
        .A2(prince_inst_sin_y[56]), .A3(prince_inst_sin_y[58]), .ZN(
        prince_inst_sbox_inst14_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst14_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst14_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst14_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst14_yyyx_inst_U15 ( .A1(prince_inst_sin_x[59]), 
        .A2(prince_inst_sin_y[58]), .A3(prince_inst_sbox_inst14_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst14_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst14_yyyx_inst_U14 ( .A(prince_inst_sin_y[56]), 
        .ZN(prince_inst_sbox_inst14_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n58), .A2(prince_inst_sin_y[57]), 
        .ZN(prince_inst_sbox_inst14_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst14_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst14_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U11 ( .A1(prince_inst_sin_y[56]), 
        .A2(prince_inst_sbox_inst14_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst14_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst14_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst14_yyyx_inst_U9 ( .A1(prince_inst_sin_y[56]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst14_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst14_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst14_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst14_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n45), .A2(prince_inst_sin_y[56]), 
        .A3(prince_inst_sin_y[58]), .ZN(prince_inst_sbox_inst14_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst14_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst14_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst14_yyyx_inst_U4 ( .A1(prince_inst_sin_x[59]), 
        .A2(prince_inst_sin_y[58]), .ZN(prince_inst_sbox_inst14_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst14_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst14_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst14_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst14_yyyx_inst_U2 ( .A(prince_inst_sin_y[57]), 
        .ZN(prince_inst_sbox_inst14_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst14_yyyx_inst_U1 ( .A1(prince_inst_sin_y[56]), 
        .A2(prince_inst_sin_x[59]), .ZN(prince_inst_sbox_inst14_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst14_mux_s00_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[0]), .B(prince_inst_sbox_inst14_s0_sh[0]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh0_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s01_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[1]), .B(prince_inst_sbox_inst14_s0_sh[1]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh0_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s02_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[2]), .B(prince_inst_sbox_inst14_s0_sh[2]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh0_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s03_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[3]), .B(prince_inst_sbox_inst14_s0_sh[3]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh0_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s04_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[4]), .B(prince_inst_sbox_inst14_s0_sh[4]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh0_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s05_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[5]), .B(prince_inst_sbox_inst14_s0_sh[5]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh0_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s06_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[6]), .B(prince_inst_sbox_inst14_s0_sh[6]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh0_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s07_U1 ( .A(
        prince_inst_sbox_inst14_t0_sh[7]), .B(prince_inst_sbox_inst14_s0_sh[7]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh0_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s10_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[0]), .B(prince_inst_sbox_inst14_s1_sh[0]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh1_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s11_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[1]), .B(prince_inst_sbox_inst14_s1_sh[1]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh1_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s12_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[2]), .B(prince_inst_sbox_inst14_s1_sh[2]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh1_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s13_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[3]), .B(prince_inst_sbox_inst14_s1_sh[3]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh1_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s14_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[4]), .B(prince_inst_sbox_inst14_s1_sh[4]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh1_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s15_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[5]), .B(prince_inst_sbox_inst14_s1_sh[5]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh1_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s16_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[6]), .B(prince_inst_sbox_inst14_s1_sh[6]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh1_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s17_U1 ( .A(
        prince_inst_sbox_inst14_t1_sh[7]), .B(prince_inst_sbox_inst14_s1_sh[7]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh1_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s20_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[0]), .B(prince_inst_sbox_inst14_s2_sh[0]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh2_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s21_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[1]), .B(prince_inst_sbox_inst14_s2_sh[1]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh2_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s22_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[2]), .B(prince_inst_sbox_inst14_s2_sh[2]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh2_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s23_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[3]), .B(prince_inst_sbox_inst14_s2_sh[3]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh2_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s24_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[4]), .B(prince_inst_sbox_inst14_s2_sh[4]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh2_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s25_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[5]), .B(prince_inst_sbox_inst14_s2_sh[5]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh2_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s26_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[6]), .B(prince_inst_sbox_inst14_s2_sh[6]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh2_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s27_U1 ( .A(
        prince_inst_sbox_inst14_t2_sh[7]), .B(prince_inst_sbox_inst14_s2_sh[7]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh2_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s30_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[0]), .B(prince_inst_sbox_inst14_s3_sh[0]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh3_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s31_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[1]), .B(prince_inst_sbox_inst14_s3_sh[1]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh3_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s32_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[2]), .B(prince_inst_sbox_inst14_s3_sh[2]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh3_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s33_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[3]), .B(prince_inst_sbox_inst14_s3_sh[3]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh3_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s34_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[4]), .B(prince_inst_sbox_inst14_s3_sh[4]), .S(prince_inst_sbox_inst14_n9), .Z(prince_inst_sbox_inst14_sh3_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s35_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[5]), .B(prince_inst_sbox_inst14_s3_sh[5]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh3_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s36_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[6]), .B(prince_inst_sbox_inst14_s3_sh[6]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh3_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst14_mux_s37_U1 ( .A(
        prince_inst_sbox_inst14_t3_sh[7]), .B(prince_inst_sbox_inst14_s3_sh[7]), .S(prince_inst_sbox_inst14_n10), .Z(prince_inst_sbox_inst14_sh3_tmp[7]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk0_U1 ( .A(r[96]), .B(
        prince_inst_sbox_inst14_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[0]), .ZN(prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk1_U1 ( .A(r[97]), .B(
        prince_inst_sbox_inst14_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[1]), .ZN(prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk2_U1 ( .A(r[98]), .B(
        prince_inst_sbox_inst14_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[2]), .ZN(prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk3_U1 ( .A(r[99]), .B(
        prince_inst_sbox_inst14_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[3]), .ZN(prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk4_U1 ( .A(r[96]), .B(
        prince_inst_sbox_inst14_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[4]), .ZN(prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk5_U1 ( .A(r[97]), .B(
        prince_inst_sbox_inst14_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[5]), .ZN(prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk6_U1 ( .A(r[98]), .B(
        prince_inst_sbox_inst14_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[6]), .ZN(prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_msk7_U1 ( .A(r[99]), .B(
        prince_inst_sbox_inst14_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst14_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst0_y[7]), .ZN(prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst14_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst14_c_inst0_ax_n5), .ZN(prince_inst_sout_x[56]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst14_c_inst0_y[1]), .B(
        prince_inst_sbox_inst14_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst14_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst14_c_inst0_y[2]), .B(
        prince_inst_sbox_inst14_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst14_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst14_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst14_c_inst0_ay_n5), .ZN(final_y[8]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst14_c_inst0_y[5]), .B(
        prince_inst_sbox_inst14_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst14_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst14_c_inst0_y[6]), .B(
        prince_inst_sbox_inst14_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst14_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk0_U1 ( .A(r[100]), .B(
        prince_inst_sbox_inst14_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[0]), .ZN(prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk1_U1 ( .A(r[101]), .B(
        prince_inst_sbox_inst14_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[1]), .ZN(prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk2_U1 ( .A(r[102]), .B(
        prince_inst_sbox_inst14_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[2]), .ZN(prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk3_U1 ( .A(r[103]), .B(
        prince_inst_sbox_inst14_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[3]), .ZN(prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk4_U1 ( .A(r[100]), .B(
        prince_inst_sbox_inst14_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[4]), .ZN(prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk5_U1 ( .A(r[101]), .B(
        prince_inst_sbox_inst14_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[5]), .ZN(prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk6_U1 ( .A(r[102]), .B(
        prince_inst_sbox_inst14_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[6]), .ZN(prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_msk7_U1 ( .A(r[103]), .B(
        prince_inst_sbox_inst14_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst14_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst1_y[7]), .ZN(prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst14_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst14_c_inst1_ax_n5), .ZN(prince_inst_sout_x[57]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst14_c_inst1_y[1]), .B(
        prince_inst_sbox_inst14_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst14_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst14_c_inst1_y[2]), .B(
        prince_inst_sbox_inst14_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst14_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst14_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst14_c_inst1_ay_n5), .ZN(final_y[9]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst14_c_inst1_y[5]), .B(
        prince_inst_sbox_inst14_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst14_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst14_c_inst1_y[6]), .B(
        prince_inst_sbox_inst14_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst14_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk0_U1 ( .A(r[104]), .B(
        prince_inst_sbox_inst14_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[0]), .ZN(prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk1_U1 ( .A(r[105]), .B(
        prince_inst_sbox_inst14_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[1]), .ZN(prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk2_U1 ( .A(r[106]), .B(
        prince_inst_sbox_inst14_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[2]), .ZN(prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk3_U1 ( .A(r[107]), .B(
        prince_inst_sbox_inst14_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[3]), .ZN(prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk4_U1 ( .A(r[104]), .B(
        prince_inst_sbox_inst14_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[4]), .ZN(prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk5_U1 ( .A(r[105]), .B(
        prince_inst_sbox_inst14_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[5]), .ZN(prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk6_U1 ( .A(r[106]), .B(
        prince_inst_sbox_inst14_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[6]), .ZN(prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_msk7_U1 ( .A(r[107]), .B(
        prince_inst_sbox_inst14_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst14_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst2_y[7]), .ZN(prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst14_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst14_c_inst2_ax_n5), .ZN(prince_inst_sout_x[58]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst14_c_inst2_y[1]), .B(
        prince_inst_sbox_inst14_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst14_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst14_c_inst2_y[2]), .B(
        prince_inst_sbox_inst14_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst14_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst14_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst14_c_inst2_ay_n5), .ZN(final_y[10]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst14_c_inst2_y[5]), .B(
        prince_inst_sbox_inst14_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst14_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst14_c_inst2_y[6]), .B(
        prince_inst_sbox_inst14_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst14_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk0_U1 ( .A(r[108]), .B(
        prince_inst_sbox_inst14_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[0]), .ZN(prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk1_U1 ( .A(r[109]), .B(
        prince_inst_sbox_inst14_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[1]), .ZN(prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk2_U1 ( .A(r[110]), .B(
        prince_inst_sbox_inst14_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[2]), .ZN(prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk3_U1 ( .A(r[111]), .B(
        prince_inst_sbox_inst14_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[3]), .ZN(prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk4_U1 ( .A(r[108]), .B(
        prince_inst_sbox_inst14_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[4]), .ZN(prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk5_U1 ( .A(r[109]), .B(
        prince_inst_sbox_inst14_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[5]), .ZN(prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk6_U1 ( .A(r[110]), .B(
        prince_inst_sbox_inst14_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[6]), .ZN(prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_msk7_U1 ( .A(r[111]), .B(
        prince_inst_sbox_inst14_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst14_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n12), .A2(
        prince_inst_sbox_inst14_n7), .A3(
        prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst14_n12), .A2(prince_inst_sbox_inst14_c_inst3_y[7]), .ZN(prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst14_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst14_n12), .ZN(
        prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst14_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst14_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst14_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst14_c_inst3_ax_n5), .ZN(prince_inst_sout_x[59]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst14_c_inst3_y[1]), .B(
        prince_inst_sbox_inst14_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst14_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst14_c_inst3_y[2]), .B(
        prince_inst_sbox_inst14_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst14_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst14_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst14_c_inst3_ay_n5), .ZN(final_y[11]) );
  XNOR2_X1 prince_inst_sbox_inst14_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst14_c_inst3_y[5]), .B(
        prince_inst_sbox_inst14_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst14_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst14_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst14_c_inst3_y[6]), .B(
        prince_inst_sbox_inst14_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst14_c_inst3_ay_n6) );
  INV_X4 prince_inst_sbox_inst15_U5 ( .A(prince_inst_sbox_inst15_n10), .ZN(
        prince_inst_sbox_inst15_n9) );
  INV_X1 prince_inst_sbox_inst15_U4 ( .A(prince_inst_n33), .ZN(
        prince_inst_sbox_inst15_n8) );
  INV_X1 prince_inst_sbox_inst15_U3 ( .A(prince_inst_sbox_inst15_n8), .ZN(
        prince_inst_sbox_inst15_n6) );
  INV_X1 prince_inst_sbox_inst15_U2 ( .A(prince_inst_sbox_inst15_n8), .ZN(
        prince_inst_sbox_inst15_n7) );
  INV_X1 prince_inst_sbox_inst15_U1 ( .A(en_sig), .ZN(
        prince_inst_sbox_inst15_n10) );
  NAND3_X1 prince_inst_sbox_inst15_xxxy_inst_U27 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n69), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n68), .A3(prince_inst_sin_x[60]), 
        .ZN(prince_inst_sbox_inst15_s3_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U26 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n66), .ZN(
        prince_inst_sbox_inst15_xxxy_inst_n68) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U25 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sbox_inst15_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst15_xxxy_inst_n69) );
  NAND3_X1 prince_inst_sbox_inst15_xxxy_inst_U24 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n64), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n63), .A3(
        prince_inst_sbox_inst15_xxxy_inst_n62), .ZN(
        prince_inst_sbox_inst15_t0_sh[0]) );
  NAND4_X1 prince_inst_sbox_inst15_xxxy_inst_U23 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n67), .A2(prince_inst_sin_x[62]), 
        .A3(prince_inst_sin_x[60]), .A4(prince_inst_sin_y[63]), .ZN(
        prince_inst_sbox_inst15_xxxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst15_xxxy_inst_U22 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n61), .A2(prince_inst_sin_x[61]), 
        .A3(prince_inst_sin_x[62]), .ZN(prince_inst_sbox_inst15_xxxy_inst_n63)
         );
  NAND4_X1 prince_inst_sbox_inst15_xxxy_inst_U21 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n66), .A3(prince_inst_sin_x[61]), 
        .A4(prince_inst_sin_x[60]), .ZN(prince_inst_sbox_inst15_xxxy_inst_n64)
         );
  XOR2_X1 prince_inst_sbox_inst15_xxxy_inst_U20 ( .A(
        prince_inst_sbox_inst15_xxxy_inst_n59), .B(prince_inst_sin_y[63]), .Z(
        prince_inst_sbox_inst15_s0_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U19 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n58), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n57), .ZN(
        prince_inst_sbox_inst15_xxxy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U18 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sin_x[61]), .ZN(prince_inst_sbox_inst15_xxxy_inst_n58)
         );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U17 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n56), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n55), .ZN(
        prince_inst_sbox_inst15_s2_sh[0]) );
  OR2_X1 prince_inst_sbox_inst15_xxxy_inst_U16 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n65), .A2(prince_inst_sin_x[62]), 
        .ZN(prince_inst_sbox_inst15_xxxy_inst_n55) );
  NAND3_X1 prince_inst_sbox_inst15_xxxy_inst_U15 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sin_y[63]), .A3(prince_inst_sbox_inst15_xxxy_inst_n67), 
        .ZN(prince_inst_sbox_inst15_xxxy_inst_n56) );
  NAND3_X1 prince_inst_sbox_inst15_xxxy_inst_U14 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n60), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n57), .A3(
        prince_inst_sbox_inst15_xxxy_inst_n54), .ZN(
        prince_inst_sbox_inst15_t3_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst15_xxxy_inst_U13 ( .A(prince_inst_sin_x[60]), 
        .B(prince_inst_sin_x[61]), .S(prince_inst_sbox_inst15_xxxy_inst_n66), 
        .Z(prince_inst_sbox_inst15_xxxy_inst_n54) );
  INV_X1 prince_inst_sbox_inst15_xxxy_inst_U12 ( .A(prince_inst_sin_y[63]), 
        .ZN(prince_inst_sbox_inst15_xxxy_inst_n66) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U11 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sin_x[60]), .ZN(prince_inst_sbox_inst15_xxxy_inst_n57)
         );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U10 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n53), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst15_s1_sh[0]) );
  MUX2_X1 prince_inst_sbox_inst15_xxxy_inst_U9 ( .A(
        prince_inst_sbox_inst15_xxxy_inst_n60), .B(
        prince_inst_sbox_inst15_xxxy_inst_n53), .S(
        prince_inst_sbox_inst15_xxxy_inst_n52), .Z(
        prince_inst_sbox_inst15_t2_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U8 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sbox_inst15_xxxy_inst_n65), .ZN(
        prince_inst_sbox_inst15_xxxy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U7 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sin_y[63]), .ZN(prince_inst_sbox_inst15_xxxy_inst_n65)
         );
  INV_X1 prince_inst_sbox_inst15_xxxy_inst_U6 ( .A(
        prince_inst_sbox_inst15_t1_sh[0]), .ZN(
        prince_inst_sbox_inst15_xxxy_inst_n53) );
  INV_X1 prince_inst_sbox_inst15_xxxy_inst_U5 ( .A(prince_inst_sin_x[62]), 
        .ZN(prince_inst_sbox_inst15_xxxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U4 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sbox_inst15_xxxy_inst_n51), .ZN(
        prince_inst_sbox_inst15_t1_sh[0]) );
  NAND2_X1 prince_inst_sbox_inst15_xxxy_inst_U3 ( .A1(
        prince_inst_sbox_inst15_xxxy_inst_n67), .A2(
        prince_inst_sbox_inst15_xxxy_inst_n61), .ZN(
        prince_inst_sbox_inst15_xxxy_inst_n51) );
  INV_X1 prince_inst_sbox_inst15_xxxy_inst_U2 ( .A(prince_inst_sin_x[60]), 
        .ZN(prince_inst_sbox_inst15_xxxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst15_xxxy_inst_U1 ( .A(prince_inst_sin_x[61]), 
        .ZN(prince_inst_sbox_inst15_xxxy_inst_n67) );
  XOR2_X1 prince_inst_sbox_inst15_xxyx_inst_U26 ( .A(
        prince_inst_sbox_inst15_t1_sh[1]), .B(
        prince_inst_sbox_inst15_xxyx_inst_n55), .Z(
        prince_inst_sbox_inst15_s1_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst15_xxyx_inst_U25 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n54), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n53), .ZN(
        prince_inst_sbox_inst15_xxyx_inst_n55) );
  XOR2_X1 prince_inst_sbox_inst15_xxyx_inst_U24 ( .A(
        prince_inst_sbox_inst15_xxyx_inst_n52), .B(
        prince_inst_sbox_inst15_xxyx_inst_n51), .Z(
        prince_inst_sbox_inst15_t1_sh[1]) );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U23 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_xxyx_inst_n51)
         );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U22 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n50), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n49), .ZN(
        prince_inst_sbox_inst15_t0_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst15_xxyx_inst_U21 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n48), .A2(prince_inst_sin_x[63]), 
        .A3(prince_inst_sin_x[60]), .ZN(prince_inst_sbox_inst15_xxyx_inst_n49)
         );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U20 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst15_xxyx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U19 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n45), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst15_s2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst15_xxyx_inst_U18 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n46), .A2(prince_inst_sin_x[63]), 
        .A3(prince_inst_sin_x[61]), .ZN(prince_inst_sbox_inst15_xxyx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U17 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n52), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n44), .ZN(
        prince_inst_sbox_inst15_t2_sh[1]) );
  NAND3_X1 prince_inst_sbox_inst15_xxyx_inst_U16 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sin_x[60]), .A3(prince_inst_sbox_inst15_xxyx_inst_n53), 
        .ZN(prince_inst_sbox_inst15_xxyx_inst_n44) );
  OR2_X1 prince_inst_sbox_inst15_xxyx_inst_U15 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sbox_inst15_xxyx_inst_n54), .ZN(
        prince_inst_sbox_inst15_xxyx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U14 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n43), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n50), .ZN(
        prince_inst_sbox_inst15_s0_sh[1]) );
  XOR2_X1 prince_inst_sbox_inst15_xxyx_inst_U13 ( .A(
        prince_inst_sbox_inst15_xxyx_inst_n54), .B(
        prince_inst_sbox_inst15_xxyx_inst_n53), .Z(
        prince_inst_sbox_inst15_xxyx_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U12 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sin_y[62]), .ZN(prince_inst_sbox_inst15_xxyx_inst_n54)
         );
  NOR4_X1 prince_inst_sbox_inst15_xxyx_inst_U11 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sbox_inst15_xxyx_inst_n42), .A3(
        prince_inst_sbox_inst15_xxyx_inst_n41), .A4(
        prince_inst_sbox_inst15_xxyx_inst_n40), .ZN(
        prince_inst_sbox_inst15_s3_sh[1]) );
  NOR2_X1 prince_inst_sbox_inst15_xxyx_inst_U10 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_xxyx_inst_n40)
         );
  NOR2_X1 prince_inst_sbox_inst15_xxyx_inst_U9 ( .A1(prince_inst_sin_x[63]), 
        .A2(prince_inst_sbox_inst15_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst15_xxyx_inst_n41) );
  NOR2_X1 prince_inst_sbox_inst15_xxyx_inst_U8 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sbox_inst15_xxyx_inst_n46), .ZN(
        prince_inst_sbox_inst15_xxyx_inst_n42) );
  INV_X1 prince_inst_sbox_inst15_xxyx_inst_U7 ( .A(prince_inst_sin_y[62]), 
        .ZN(prince_inst_sbox_inst15_xxyx_inst_n46) );
  NAND2_X1 prince_inst_sbox_inst15_xxyx_inst_U6 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n39), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n38), .ZN(
        prince_inst_sbox_inst15_t3_sh[1]) );
  NAND4_X1 prince_inst_sbox_inst15_xxyx_inst_U5 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n53), .A2(prince_inst_sin_x[61]), 
        .A3(prince_inst_sin_y[62]), .A4(prince_inst_sin_x[60]), .ZN(
        prince_inst_sbox_inst15_xxyx_inst_n38) );
  INV_X1 prince_inst_sbox_inst15_xxyx_inst_U4 ( .A(prince_inst_sin_x[63]), 
        .ZN(prince_inst_sbox_inst15_xxyx_inst_n53) );
  NAND4_X1 prince_inst_sbox_inst15_xxyx_inst_U3 ( .A1(
        prince_inst_sbox_inst15_xxyx_inst_n47), .A2(
        prince_inst_sbox_inst15_xxyx_inst_n43), .A3(prince_inst_sin_x[63]), 
        .A4(prince_inst_sin_y[62]), .ZN(prince_inst_sbox_inst15_xxyx_inst_n39)
         );
  INV_X1 prince_inst_sbox_inst15_xxyx_inst_U2 ( .A(prince_inst_sin_x[60]), 
        .ZN(prince_inst_sbox_inst15_xxyx_inst_n43) );
  INV_X1 prince_inst_sbox_inst15_xxyx_inst_U1 ( .A(prince_inst_sin_x[61]), 
        .ZN(prince_inst_sbox_inst15_xxyx_inst_n47) );
  XNOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U30 ( .A(
        prince_inst_sbox_inst15_xyxx_inst_n74), .B(
        prince_inst_sbox_inst15_xyxx_inst_n73), .ZN(
        prince_inst_sbox_inst15_t0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U29 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n71), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n73) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U28 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n69), .ZN(
        prince_inst_sbox_inst15_t3_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst15_xyxx_inst_U27 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n68), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst15_xyxx_inst_n66), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U26 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sbox_inst15_xyxx_inst_n65), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n66) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U25 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_xyxx_inst_n65)
         );
  MUX2_X1 prince_inst_sbox_inst15_xyxx_inst_U24 ( .A(
        prince_inst_sbox_inst15_xyxx_inst_n72), .B(
        prince_inst_sbox_inst15_s0_sh[2]), .S(
        prince_inst_sbox_inst15_xyxx_inst_n64), .Z(
        prince_inst_sbox_inst15_t2_sh[2]) );
  NAND2_X1 prince_inst_sbox_inst15_xyxx_inst_U23 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n74), .A2(prince_inst_sin_x[63]), 
        .ZN(prince_inst_sbox_inst15_xyxx_inst_n64) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U22 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n63), .ZN(
        prince_inst_sbox_inst15_s0_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U21 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sbox_inst15_xyxx_inst_n74), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n63) );
  INV_X1 prince_inst_sbox_inst15_xyxx_inst_U20 ( .A(
        prince_inst_sbox_inst15_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U19 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n71), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n61), .ZN(
        prince_inst_sbox_inst15_s3_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U18 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n60), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n68), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n61) );
  INV_X1 prince_inst_sbox_inst15_xyxx_inst_U17 ( .A(
        prince_inst_sbox_inst15_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n68) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U16 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n67), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n62), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst15_xyxx_inst_U15 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_x[60]), .ZN(prince_inst_sbox_inst15_xyxx_inst_n62)
         );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U14 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n70), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n59), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n71) );
  NAND2_X1 prince_inst_sbox_inst15_xyxx_inst_U13 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_xyxx_inst_n59)
         );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U12 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_x[62]), .ZN(prince_inst_sbox_inst15_xyxx_inst_n70)
         );
  XNOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U11 ( .A(
        prince_inst_sbox_inst15_xyxx_inst_n58), .B(
        prince_inst_sbox_inst15_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst15_t1_sh[2]) );
  NOR3_X1 prince_inst_sbox_inst15_xyxx_inst_U10 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n72), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n56), .A3(
        prince_inst_sbox_inst15_xyxx_inst_n55), .ZN(
        prince_inst_sbox_inst15_s2_sh[2]) );
  INV_X1 prince_inst_sbox_inst15_xyxx_inst_U9 ( .A(prince_inst_sin_x[63]), 
        .ZN(prince_inst_sbox_inst15_xyxx_inst_n55) );
  AND2_X1 prince_inst_sbox_inst15_xyxx_inst_U8 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n54), .A2(prince_inst_sin_x[60]), 
        .ZN(prince_inst_sbox_inst15_xyxx_inst_n56) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U7 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n54), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n67), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n72) );
  OR2_X1 prince_inst_sbox_inst15_xyxx_inst_U6 ( .A1(
        prince_inst_sbox_inst15_xyxx_inst_n58), .A2(
        prince_inst_sbox_inst15_xyxx_inst_n53), .ZN(
        prince_inst_sbox_inst15_s1_sh[2]) );
  NOR2_X1 prince_inst_sbox_inst15_xyxx_inst_U5 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sbox_inst15_xyxx_inst_n57), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst15_xyxx_inst_U4 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_xyxx_inst_n57)
         );
  NOR3_X1 prince_inst_sbox_inst15_xyxx_inst_U3 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sbox_inst15_xyxx_inst_n67), .A3(
        prince_inst_sbox_inst15_xyxx_inst_n54), .ZN(
        prince_inst_sbox_inst15_xyxx_inst_n58) );
  INV_X1 prince_inst_sbox_inst15_xyxx_inst_U2 ( .A(prince_inst_sin_y[61]), 
        .ZN(prince_inst_sbox_inst15_xyxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst15_xyxx_inst_U1 ( .A(prince_inst_sin_x[62]), 
        .ZN(prince_inst_sbox_inst15_xyxx_inst_n67) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U28 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n61), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n60), .ZN(
        prince_inst_sbox_inst15_s2_sh[3]) );
  XOR2_X1 prince_inst_sbox_inst15_xyyy_inst_U27 ( .A(
        prince_inst_sbox_inst15_xyyy_inst_n59), .B(
        prince_inst_sbox_inst15_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst15_xyyy_inst_n61) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U26 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n57), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n56), .ZN(
        prince_inst_sbox_inst15_t3_sh[3]) );
  OR3_X1 prince_inst_sbox_inst15_xyyy_inst_U25 ( .A1(prince_inst_sin_y[62]), 
        .A2(prince_inst_sin_y[63]), .A3(prince_inst_sbox_inst15_xyyy_inst_n60), 
        .ZN(prince_inst_sbox_inst15_xyyy_inst_n56) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U24 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sbox_inst15_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U23 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sbox_inst15_xyyy_inst_n54), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n57) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U22 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n53), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n52), .ZN(
        prince_inst_sbox_inst15_s3_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U21 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n51), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U20 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n54), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n55), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n53) );
  NOR3_X1 prince_inst_sbox_inst15_xyyy_inst_U19 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sin_y[62]), .A3(prince_inst_sbox_inst15_xyyy_inst_n50), 
        .ZN(prince_inst_sbox_inst15_xyyy_inst_n54) );
  MUX2_X1 prince_inst_sbox_inst15_xyyy_inst_U18 ( .A(
        prince_inst_sbox_inst15_xyyy_inst_n49), .B(
        prince_inst_sbox_inst15_xyyy_inst_n48), .S(
        prince_inst_sbox_inst15_xyyy_inst_n47), .Z(
        prince_inst_sbox_inst15_s0_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst15_xyyy_inst_U17 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n51), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n49) );
  NOR2_X1 prince_inst_sbox_inst15_xyyy_inst_U16 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sbox_inst15_xyyy_inst_n46), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst15_xyyy_inst_U15 ( .A(
        prince_inst_sbox_inst15_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n46) );
  NOR3_X1 prince_inst_sbox_inst15_xyyy_inst_U14 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n44), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n43), .A3(
        prince_inst_sbox_inst15_xyyy_inst_n58), .ZN(
        prince_inst_sbox_inst15_t0_sh[3]) );
  NOR3_X1 prince_inst_sbox_inst15_xyyy_inst_U13 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n42), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n48), .A3(
        prince_inst_sbox_inst15_xyyy_inst_n50), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n43) );
  INV_X1 prince_inst_sbox_inst15_xyyy_inst_U12 ( .A(prince_inst_sin_y[63]), 
        .ZN(prince_inst_sbox_inst15_xyyy_inst_n50) );
  NOR2_X1 prince_inst_sbox_inst15_xyyy_inst_U11 ( .A1(prince_inst_sin_y[63]), 
        .A2(prince_inst_sbox_inst15_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n44) );
  MUX2_X1 prince_inst_sbox_inst15_xyyy_inst_U10 ( .A(
        prince_inst_sbox_inst15_t1_sh[3]), .B(
        prince_inst_sbox_inst15_xyyy_inst_n48), .S(
        prince_inst_sbox_inst15_xyyy_inst_n58), .Z(
        prince_inst_sbox_inst15_t2_sh[3]) );
  AND2_X1 prince_inst_sbox_inst15_xyyy_inst_U9 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sbox_inst15_xyyy_inst_n47), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n58) );
  AND2_X1 prince_inst_sbox_inst15_xyyy_inst_U8 ( .A1(prince_inst_sin_x[60]), 
        .A2(prince_inst_sin_y[63]), .ZN(prince_inst_sbox_inst15_xyyy_inst_n47)
         );
  AND2_X1 prince_inst_sbox_inst15_xyyy_inst_U7 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n59), .A2(
        prince_inst_sbox_inst15_t1_sh[3]), .ZN(
        prince_inst_sbox_inst15_s1_sh[3]) );
  NAND2_X1 prince_inst_sbox_inst15_xyyy_inst_U6 ( .A1(prince_inst_sin_y[63]), 
        .A2(prince_inst_sbox_inst15_xyyy_inst_n45), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst15_xyyy_inst_U5 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n55), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n48), .ZN(
        prince_inst_sbox_inst15_xyyy_inst_n45) );
  INV_X1 prince_inst_sbox_inst15_xyyy_inst_U4 ( .A(prince_inst_sin_y[61]), 
        .ZN(prince_inst_sbox_inst15_xyyy_inst_n55) );
  NOR2_X1 prince_inst_sbox_inst15_xyyy_inst_U3 ( .A1(
        prince_inst_sbox_inst15_xyyy_inst_n48), .A2(
        prince_inst_sbox_inst15_xyyy_inst_n42), .ZN(
        prince_inst_sbox_inst15_t1_sh[3]) );
  NOR2_X1 prince_inst_sbox_inst15_xyyy_inst_U2 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_x[60]), .ZN(prince_inst_sbox_inst15_xyyy_inst_n42)
         );
  INV_X1 prince_inst_sbox_inst15_xyyy_inst_U1 ( .A(prince_inst_sin_y[62]), 
        .ZN(prince_inst_sbox_inst15_xyyy_inst_n48) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U28 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n64), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n63), .ZN(
        prince_inst_sbox_inst15_t2_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U27 ( .A1(prince_inst_sin_y[60]), 
        .A2(prince_inst_sbox_inst15_yxxx_inst_n62), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U26 ( .A1(prince_inst_sin_y[60]), 
        .A2(prince_inst_sbox_inst15_yxxx_inst_n61), .ZN(
        prince_inst_sbox_inst15_s3_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U25 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n62), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n60), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n61) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U24 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n59), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n58), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n60) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U23 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_yxxx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U22 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n57), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n62) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U21 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n54), .ZN(
        prince_inst_sbox_inst15_t3_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U20 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n53), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n56), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n54) );
  INV_X1 prince_inst_sbox_inst15_yxxx_inst_U19 ( .A(prince_inst_sin_x[63]), 
        .ZN(prince_inst_sbox_inst15_yxxx_inst_n56) );
  MUX2_X1 prince_inst_sbox_inst15_yxxx_inst_U18 ( .A(
        prince_inst_sbox_inst15_yxxx_inst_n52), .B(
        prince_inst_sbox_inst15_yxxx_inst_n51), .S(
        prince_inst_sbox_inst15_yxxx_inst_n50), .Z(
        prince_inst_sbox_inst15_t0_sh[4]) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U17 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n57), .A2(prince_inst_sin_x[63]), 
        .ZN(prince_inst_sbox_inst15_yxxx_inst_n52) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U16 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n55), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n49), .ZN(
        prince_inst_sbox_inst15_s2_sh[4]) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U15 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n48), .A2(prince_inst_sin_y[60]), 
        .ZN(prince_inst_sbox_inst15_yxxx_inst_n49) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U14 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n47), .A2(prince_inst_sin_x[63]), 
        .ZN(prince_inst_sbox_inst15_yxxx_inst_n48) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U13 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sbox_inst15_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n47) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U12 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n55) );
  XNOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U11 ( .A(
        prince_inst_sbox_inst15_yxxx_inst_n53), .B(
        prince_inst_sbox_inst15_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst15_t1_sh[4]) );
  OR2_X1 prince_inst_sbox_inst15_yxxx_inst_U10 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n46), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n53), .ZN(
        prince_inst_sbox_inst15_s1_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst15_yxxx_inst_U9 ( .A1(prince_inst_sin_x[61]), 
        .A2(prince_inst_sbox_inst15_yxxx_inst_n50), .A3(
        prince_inst_sbox_inst15_yxxx_inst_n59), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n53) );
  INV_X1 prince_inst_sbox_inst15_yxxx_inst_U8 ( .A(prince_inst_sin_x[62]), 
        .ZN(prince_inst_sbox_inst15_yxxx_inst_n59) );
  NOR2_X1 prince_inst_sbox_inst15_yxxx_inst_U7 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n57), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n46) );
  OR2_X1 prince_inst_sbox_inst15_yxxx_inst_U6 ( .A1(
        prince_inst_sbox_inst15_yxxx_inst_n51), .A2(
        prince_inst_sbox_inst15_yxxx_inst_n64), .ZN(
        prince_inst_sbox_inst15_s0_sh[4]) );
  NOR3_X1 prince_inst_sbox_inst15_yxxx_inst_U5 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sbox_inst15_yxxx_inst_n57), .A3(
        prince_inst_sbox_inst15_yxxx_inst_n50), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n64) );
  INV_X1 prince_inst_sbox_inst15_yxxx_inst_U4 ( .A(prince_inst_sin_y[60]), 
        .ZN(prince_inst_sbox_inst15_yxxx_inst_n50) );
  INV_X1 prince_inst_sbox_inst15_yxxx_inst_U3 ( .A(prince_inst_sin_x[61]), 
        .ZN(prince_inst_sbox_inst15_yxxx_inst_n57) );
  INV_X1 prince_inst_sbox_inst15_yxxx_inst_U2 ( .A(
        prince_inst_sbox_inst15_yxxx_inst_n45), .ZN(
        prince_inst_sbox_inst15_yxxx_inst_n51) );
  NAND2_X1 prince_inst_sbox_inst15_yxxx_inst_U1 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_yxxx_inst_n45)
         );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U28 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n68), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n67), .ZN(
        prince_inst_sbox_inst15_s1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst15_yxyy_inst_U27 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n66), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n67), .A3(
        prince_inst_sbox_inst15_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst15_t1_sh[5]) );
  NAND3_X1 prince_inst_sbox_inst15_yxyy_inst_U26 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n64), .A3(prince_inst_sin_y[63]), 
        .ZN(prince_inst_sbox_inst15_yxyy_inst_n67) );
  NAND3_X1 prince_inst_sbox_inst15_yxyy_inst_U25 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n63), .A2(prince_inst_sin_y[62]), 
        .A3(prince_inst_sin_y[63]), .ZN(prince_inst_sbox_inst15_yxyy_inst_n66)
         );
  MUX2_X1 prince_inst_sbox_inst15_yxyy_inst_U24 ( .A(
        prince_inst_sbox_inst15_yxyy_inst_n62), .B(
        prince_inst_sbox_inst15_yxyy_inst_n61), .S(prince_inst_sin_y[60]), .Z(
        prince_inst_sbox_inst15_t2_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst15_yxyy_inst_U23 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n61) );
  MUX2_X1 prince_inst_sbox_inst15_yxyy_inst_U22 ( .A(
        prince_inst_sbox_inst15_yxyy_inst_n64), .B(
        prince_inst_sbox_inst15_yxyy_inst_n60), .S(
        prince_inst_sbox_inst15_yxyy_inst_n65), .Z(
        prince_inst_sbox_inst15_t3_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U21 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n59), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n58), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U20 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n57), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n59) );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U19 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n56), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst15_yxyy_inst_U18 ( .A(
        prince_inst_sbox_inst15_yxyy_inst_n62), .B(
        prince_inst_sbox_inst15_yxyy_inst_n54), .S(
        prince_inst_sbox_inst15_yxyy_inst_n55), .Z(
        prince_inst_sbox_inst15_t0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst15_yxyy_inst_U17 ( .A(
        prince_inst_sbox_inst15_yxyy_inst_n53), .B(
        prince_inst_sbox_inst15_yxyy_inst_n54), .Z(
        prince_inst_sbox_inst15_s0_sh[5]) );
  XOR2_X1 prince_inst_sbox_inst15_yxyy_inst_U16 ( .A(
        prince_inst_sbox_inst15_yxyy_inst_n68), .B(
        prince_inst_sbox_inst15_yxyy_inst_n58), .Z(
        prince_inst_sbox_inst15_yxyy_inst_n53) );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U15 ( .A1(prince_inst_sin_y[63]), 
        .A2(prince_inst_sin_y[60]), .ZN(prince_inst_sbox_inst15_yxyy_inst_n58)
         );
  NOR4_X1 prince_inst_sbox_inst15_yxyy_inst_U14 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n52), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n54), .A3(
        prince_inst_sbox_inst15_yxyy_inst_n62), .A4(
        prince_inst_sbox_inst15_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst15_s3_sh[5]) );
  NOR2_X1 prince_inst_sbox_inst15_yxyy_inst_U13 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n63), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n62) );
  INV_X1 prince_inst_sbox_inst15_yxyy_inst_U12 ( .A(
        prince_inst_sbox_inst15_yxyy_inst_n68), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst15_yxyy_inst_U11 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n64), .A2(prince_inst_sin_y[62]), 
        .A3(prince_inst_sin_y[60]), .ZN(prince_inst_sbox_inst15_yxyy_inst_n68)
         );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U10 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n51), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n50), .ZN(
        prince_inst_sbox_inst15_s2_sh[5]) );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U9 ( .A1(prince_inst_sin_y[63]), 
        .A2(prince_inst_sbox_inst15_yxyy_inst_n49), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n50) );
  NAND2_X1 prince_inst_sbox_inst15_yxyy_inst_U8 ( .A1(prince_inst_sin_y[62]), 
        .A2(prince_inst_sbox_inst15_yxyy_inst_n64), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n49) );
  INV_X1 prince_inst_sbox_inst15_yxyy_inst_U7 ( .A(
        prince_inst_sbox_inst15_yxyy_inst_n63), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n64) );
  OR3_X1 prince_inst_sbox_inst15_yxyy_inst_U6 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n54), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n63), .A3(
        prince_inst_sbox_inst15_yxyy_inst_n55), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n51) );
  INV_X1 prince_inst_sbox_inst15_yxyy_inst_U5 ( .A(prince_inst_sin_y[60]), 
        .ZN(prince_inst_sbox_inst15_yxyy_inst_n55) );
  INV_X1 prince_inst_sbox_inst15_yxyy_inst_U4 ( .A(prince_inst_sin_x[61]), 
        .ZN(prince_inst_sbox_inst15_yxyy_inst_n63) );
  NOR2_X1 prince_inst_sbox_inst15_yxyy_inst_U3 ( .A1(
        prince_inst_sbox_inst15_yxyy_inst_n65), .A2(
        prince_inst_sbox_inst15_yxyy_inst_n56), .ZN(
        prince_inst_sbox_inst15_yxyy_inst_n54) );
  INV_X1 prince_inst_sbox_inst15_yxyy_inst_U2 ( .A(prince_inst_sin_y[63]), 
        .ZN(prince_inst_sbox_inst15_yxyy_inst_n56) );
  INV_X1 prince_inst_sbox_inst15_yxyy_inst_U1 ( .A(prince_inst_sin_y[62]), 
        .ZN(prince_inst_sbox_inst15_yxyy_inst_n65) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U31 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n75), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n74), .ZN(
        prince_inst_sbox_inst15_s1_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U30 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n73), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n72), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n74) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U29 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sbox_inst15_yyxy_inst_n71), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n72) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U28 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n70), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n73) );
  NAND2_X1 prince_inst_sbox_inst15_yyxy_inst_U27 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n68), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n67), .ZN(
        prince_inst_sbox_inst15_s3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst15_yyxy_inst_U26 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n75), .A2(prince_inst_sin_y[63]), 
        .A3(prince_inst_sbox_inst15_yyxy_inst_n70), .A4(prince_inst_sin_x[62]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n67) );
  NAND4_X1 prince_inst_sbox_inst15_yyxy_inst_U25 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n69), .A3(prince_inst_sin_y[61]), 
        .A4(prince_inst_sbox_inst15_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n68) );
  NAND3_X1 prince_inst_sbox_inst15_yyxy_inst_U24 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n66), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n65), .A3(
        prince_inst_sbox_inst15_yyxy_inst_n64), .ZN(
        prince_inst_sbox_inst15_t1_sh[6]) );
  NAND3_X1 prince_inst_sbox_inst15_yyxy_inst_U23 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_x[62]), .A3(prince_inst_sin_y[60]), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n64) );
  NAND3_X1 prince_inst_sbox_inst15_yyxy_inst_U22 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n69), .A2(prince_inst_sin_y[61]), 
        .A3(prince_inst_sin_y[63]), .ZN(prince_inst_sbox_inst15_yyxy_inst_n65)
         );
  NAND3_X1 prince_inst_sbox_inst15_yyxy_inst_U21 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n75), .A2(prince_inst_sin_x[62]), 
        .A3(prince_inst_sin_y[63]), .ZN(prince_inst_sbox_inst15_yyxy_inst_n66)
         );
  NAND2_X1 prince_inst_sbox_inst15_yyxy_inst_U20 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n63), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n62), .ZN(
        prince_inst_sbox_inst15_t2_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst15_yyxy_inst_U19 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n61), .A2(prince_inst_sin_x[62]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n62) );
  NAND3_X1 prince_inst_sbox_inst15_yyxy_inst_U18 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_y[63]), .A3(prince_inst_sbox_inst15_yyxy_inst_n70), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n63) );
  NAND2_X1 prince_inst_sbox_inst15_yyxy_inst_U17 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n60), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n59), .ZN(
        prince_inst_sbox_inst15_t3_sh[6]) );
  NAND4_X1 prince_inst_sbox_inst15_yyxy_inst_U16 ( .A1(prince_inst_sin_y[63]), 
        .A2(prince_inst_sbox_inst15_yyxy_inst_n70), .A3(
        prince_inst_sbox_inst15_yyxy_inst_n75), .A4(
        prince_inst_sbox_inst15_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n59) );
  NAND3_X1 prince_inst_sbox_inst15_yyxy_inst_U15 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n58), .A3(prince_inst_sin_y[60]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n60) );
  NAND2_X1 prince_inst_sbox_inst15_yyxy_inst_U14 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n57), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n56), .ZN(
        prince_inst_sbox_inst15_s0_sh[6]) );
  NAND2_X1 prince_inst_sbox_inst15_yyxy_inst_U13 ( .A1(prince_inst_sin_y[60]), 
        .A2(prince_inst_sbox_inst15_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n56) );
  INV_X1 prince_inst_sbox_inst15_yyxy_inst_U12 ( .A(
        prince_inst_sbox_inst15_yyxy_inst_n55), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n57) );
  MUX2_X1 prince_inst_sbox_inst15_yyxy_inst_U11 ( .A(
        prince_inst_sbox_inst15_yyxy_inst_n54), .B(
        prince_inst_sbox_inst15_yyxy_inst_n55), .S(
        prince_inst_sbox_inst15_yyxy_inst_n70), .Z(
        prince_inst_sbox_inst15_t0_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U10 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n69), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n55) );
  INV_X1 prince_inst_sbox_inst15_yyxy_inst_U9 ( .A(prince_inst_sin_x[62]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n69) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U8 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n75), .A2(prince_inst_sin_y[63]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n54) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U7 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n71), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n53), .ZN(
        prince_inst_sbox_inst15_s2_sh[6]) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U6 ( .A1(
        prince_inst_sbox_inst15_yyxy_inst_n61), .A2(
        prince_inst_sbox_inst15_yyxy_inst_n58), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n53) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U5 ( .A1(prince_inst_sin_x[62]), 
        .A2(prince_inst_sbox_inst15_yyxy_inst_n75), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n58) );
  INV_X1 prince_inst_sbox_inst15_yyxy_inst_U4 ( .A(prince_inst_sin_y[61]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n75) );
  NOR2_X1 prince_inst_sbox_inst15_yyxy_inst_U3 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sbox_inst15_yyxy_inst_n70), .ZN(
        prince_inst_sbox_inst15_yyxy_inst_n61) );
  INV_X1 prince_inst_sbox_inst15_yyxy_inst_U2 ( .A(prince_inst_sin_y[60]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n70) );
  INV_X1 prince_inst_sbox_inst15_yyxy_inst_U1 ( .A(prince_inst_sin_y[63]), 
        .ZN(prince_inst_sbox_inst15_yyxy_inst_n71) );
  XNOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U25 ( .A(
        prince_inst_sbox_inst15_yyyx_inst_n58), .B(
        prince_inst_sbox_inst15_yyyx_inst_n57), .ZN(
        prince_inst_sbox_inst15_s0_sh[7]) );
  XOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U24 ( .A(
        prince_inst_sbox_inst15_yyyx_inst_n56), .B(
        prince_inst_sbox_inst15_yyyx_inst_n55), .Z(
        prince_inst_sbox_inst15_yyyx_inst_n57) );
  XNOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U23 ( .A(
        prince_inst_sbox_inst15_yyyx_inst_n54), .B(
        prince_inst_sbox_inst15_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst15_t1_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst15_yyyx_inst_U22 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n53), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n52), .ZN(
        prince_inst_sbox_inst15_t3_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst15_yyyx_inst_U21 ( .A1(prince_inst_sin_x[63]), 
        .A2(prince_inst_sbox_inst15_yyyx_inst_n54), .ZN(
        prince_inst_sbox_inst15_yyyx_inst_n52) );
  NAND3_X1 prince_inst_sbox_inst15_yyyx_inst_U20 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_y[62]), .A3(prince_inst_sbox_inst15_yyyx_inst_n51), 
        .ZN(prince_inst_sbox_inst15_yyyx_inst_n53) );
  XNOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U19 ( .A(
        prince_inst_sbox_inst15_yyyx_inst_n50), .B(
        prince_inst_sbox_inst15_yyyx_inst_n49), .ZN(
        prince_inst_sbox_inst15_t2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst15_yyyx_inst_U18 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n56), .A2(prince_inst_sin_y[62]), 
        .ZN(prince_inst_sbox_inst15_yyyx_inst_n50) );
  NAND3_X1 prince_inst_sbox_inst15_yyyx_inst_U17 ( .A1(prince_inst_sin_y[61]), 
        .A2(prince_inst_sin_y[60]), .A3(prince_inst_sin_y[62]), .ZN(
        prince_inst_sbox_inst15_yyyx_inst_n56) );
  NOR3_X1 prince_inst_sbox_inst15_yyyx_inst_U16 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n48), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n47), .A3(
        prince_inst_sbox_inst15_yyyx_inst_n46), .ZN(
        prince_inst_sbox_inst15_s3_sh[7]) );
  NOR3_X1 prince_inst_sbox_inst15_yyyx_inst_U15 ( .A1(prince_inst_sin_x[63]), 
        .A2(prince_inst_sin_y[62]), .A3(prince_inst_sbox_inst15_yyyx_inst_n45), 
        .ZN(prince_inst_sbox_inst15_yyyx_inst_n46) );
  INV_X1 prince_inst_sbox_inst15_yyyx_inst_U14 ( .A(prince_inst_sin_y[60]), 
        .ZN(prince_inst_sbox_inst15_yyyx_inst_n47) );
  NOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U13 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n58), .A2(prince_inst_sin_y[61]), 
        .ZN(prince_inst_sbox_inst15_yyyx_inst_n48) );
  OR2_X1 prince_inst_sbox_inst15_yyyx_inst_U12 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n44), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n43), .ZN(
        prince_inst_sbox_inst15_t0_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U11 ( .A1(prince_inst_sin_y[60]), 
        .A2(prince_inst_sbox_inst15_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst15_yyyx_inst_n43) );
  NOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U10 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n55), .ZN(
        prince_inst_sbox_inst15_yyyx_inst_n44) );
  NAND2_X1 prince_inst_sbox_inst15_yyyx_inst_U9 ( .A1(prince_inst_sin_y[60]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_yyyx_inst_n55)
         );
  OR2_X1 prince_inst_sbox_inst15_yyyx_inst_U8 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n54), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n42), .ZN(
        prince_inst_sbox_inst15_s1_sh[7]) );
  NOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U7 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n45), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst15_yyyx_inst_n42) );
  AND3_X1 prince_inst_sbox_inst15_yyyx_inst_U6 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n45), .A2(prince_inst_sin_y[60]), 
        .A3(prince_inst_sin_y[62]), .ZN(prince_inst_sbox_inst15_yyyx_inst_n54)
         );
  AND2_X1 prince_inst_sbox_inst15_yyyx_inst_U5 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n49), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n58), .ZN(
        prince_inst_sbox_inst15_s2_sh[7]) );
  NAND2_X1 prince_inst_sbox_inst15_yyyx_inst_U4 ( .A1(prince_inst_sin_x[63]), 
        .A2(prince_inst_sin_y[62]), .ZN(prince_inst_sbox_inst15_yyyx_inst_n58)
         );
  NOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U3 ( .A1(
        prince_inst_sbox_inst15_yyyx_inst_n51), .A2(
        prince_inst_sbox_inst15_yyyx_inst_n45), .ZN(
        prince_inst_sbox_inst15_yyyx_inst_n49) );
  INV_X1 prince_inst_sbox_inst15_yyyx_inst_U2 ( .A(prince_inst_sin_y[61]), 
        .ZN(prince_inst_sbox_inst15_yyyx_inst_n45) );
  NOR2_X1 prince_inst_sbox_inst15_yyyx_inst_U1 ( .A1(prince_inst_sin_y[60]), 
        .A2(prince_inst_sin_x[63]), .ZN(prince_inst_sbox_inst15_yyyx_inst_n51)
         );
  MUX2_X1 prince_inst_sbox_inst15_mux_s00_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[0]), .B(prince_inst_sbox_inst15_s0_sh[0]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh0_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s01_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[1]), .B(prince_inst_sbox_inst15_s0_sh[1]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh0_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s02_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[2]), .B(prince_inst_sbox_inst15_s0_sh[2]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh0_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s03_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[3]), .B(prince_inst_sbox_inst15_s0_sh[3]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh0_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s04_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[4]), .B(prince_inst_sbox_inst15_s0_sh[4]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh0_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s05_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[5]), .B(prince_inst_sbox_inst15_s0_sh[5]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh0_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s06_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[6]), .B(prince_inst_sbox_inst15_s0_sh[6]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh0_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s07_U1 ( .A(
        prince_inst_sbox_inst15_t0_sh[7]), .B(prince_inst_sbox_inst15_s0_sh[7]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh0_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s10_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[0]), .B(prince_inst_sbox_inst15_s1_sh[0]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh1_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s11_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[1]), .B(prince_inst_sbox_inst15_s1_sh[1]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh1_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s12_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[2]), .B(prince_inst_sbox_inst15_s1_sh[2]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh1_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s13_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[3]), .B(prince_inst_sbox_inst15_s1_sh[3]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh1_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s14_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[4]), .B(prince_inst_sbox_inst15_s1_sh[4]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh1_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s15_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[5]), .B(prince_inst_sbox_inst15_s1_sh[5]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh1_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s16_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[6]), .B(prince_inst_sbox_inst15_s1_sh[6]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh1_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s17_U1 ( .A(
        prince_inst_sbox_inst15_t1_sh[7]), .B(prince_inst_sbox_inst15_s1_sh[7]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh1_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s20_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[0]), .B(prince_inst_sbox_inst15_s2_sh[0]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh2_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s21_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[1]), .B(prince_inst_sbox_inst15_s2_sh[1]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh2_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s22_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[2]), .B(prince_inst_sbox_inst15_s2_sh[2]), .S(prince_inst_n33), .Z(prince_inst_sbox_inst15_sh2_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s23_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[3]), .B(prince_inst_sbox_inst15_s2_sh[3]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh2_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s24_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[4]), .B(prince_inst_sbox_inst15_s2_sh[4]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh2_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s25_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[5]), .B(prince_inst_sbox_inst15_s2_sh[5]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh2_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s26_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[6]), .B(prince_inst_sbox_inst15_s2_sh[6]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh2_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s27_U1 ( .A(
        prince_inst_sbox_inst15_t2_sh[7]), .B(prince_inst_sbox_inst15_s2_sh[7]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh2_tmp[7]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s30_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[0]), .B(prince_inst_sbox_inst15_s3_sh[0]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh3_tmp[0]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s31_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[1]), .B(prince_inst_sbox_inst15_s3_sh[1]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh3_tmp[1]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s32_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[2]), .B(prince_inst_sbox_inst15_s3_sh[2]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh3_tmp[2]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s33_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[3]), .B(prince_inst_sbox_inst15_s3_sh[3]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh3_tmp[3]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s34_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[4]), .B(prince_inst_sbox_inst15_s3_sh[4]), .S(prince_inst_sbox_inst15_n6), .Z(prince_inst_sbox_inst15_sh3_tmp[4]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s35_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[5]), .B(prince_inst_sbox_inst15_s3_sh[5]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh3_tmp[5]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s36_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[6]), .B(prince_inst_sbox_inst15_s3_sh[6]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh3_tmp[6]) );
  MUX2_X1 prince_inst_sbox_inst15_mux_s37_U1 ( .A(
        prince_inst_sbox_inst15_t3_sh[7]), .B(prince_inst_sbox_inst15_s3_sh[7]), .S(prince_inst_sbox_inst15_n7), .Z(prince_inst_sbox_inst15_sh3_tmp[7]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk0_U1 ( .A(r[112]), .B(
        prince_inst_sbox_inst15_sh0_tmp[0]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[0]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk0_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[0]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk1_U1 ( .A(r[113]), .B(
        prince_inst_sbox_inst15_sh0_tmp[1]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[1]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk1_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[1]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk2_U1 ( .A(r[114]), .B(
        prince_inst_sbox_inst15_sh0_tmp[2]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[2]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk2_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[2]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk3_U1 ( .A(r[115]), .B(
        prince_inst_sbox_inst15_sh0_tmp[3]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[3]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk3_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[3]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk4_U1 ( .A(r[112]), .B(
        prince_inst_sbox_inst15_sh0_tmp[4]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[4]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk4_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[4]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk5_U1 ( .A(r[113]), .B(
        prince_inst_sbox_inst15_sh0_tmp[5]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[5]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk5_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[5]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk6_U1 ( .A(r[114]), .B(
        prince_inst_sbox_inst15_sh0_tmp[6]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[6]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk6_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[6]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_msk7_U1 ( .A(r[115]), .B(
        prince_inst_sbox_inst15_sh0_tmp[7]), .Z(
        prince_inst_sbox_inst15_c_inst0_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst0_y[7]), 
        .ZN(prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst0_msk7_xr), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst0_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst0_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst0_ax_U3 ( .A(
        prince_inst_sbox_inst15_c_inst0_ax_n6), .B(
        prince_inst_sbox_inst15_c_inst0_ax_n5), .ZN(prince_inst_sout_x[60]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst0_ax_U2 ( .A(
        prince_inst_sbox_inst15_c_inst0_y[1]), .B(
        prince_inst_sbox_inst15_c_inst0_y[0]), .ZN(
        prince_inst_sbox_inst15_c_inst0_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_ax_U1 ( .A(
        prince_inst_sbox_inst15_c_inst0_y[2]), .B(
        prince_inst_sbox_inst15_c_inst0_y[3]), .Z(
        prince_inst_sbox_inst15_c_inst0_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst0_ay_U3 ( .A(
        prince_inst_sbox_inst15_c_inst0_ay_n6), .B(
        prince_inst_sbox_inst15_c_inst0_ay_n5), .ZN(final_y[60]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst0_ay_U2 ( .A(
        prince_inst_sbox_inst15_c_inst0_y[5]), .B(
        prince_inst_sbox_inst15_c_inst0_y[4]), .ZN(
        prince_inst_sbox_inst15_c_inst0_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst0_ay_U1 ( .A(
        prince_inst_sbox_inst15_c_inst0_y[6]), .B(
        prince_inst_sbox_inst15_c_inst0_y[7]), .Z(
        prince_inst_sbox_inst15_c_inst0_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk0_U1 ( .A(r[116]), .B(
        prince_inst_sbox_inst15_sh1_tmp[0]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[0]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk0_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[0]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk1_U1 ( .A(r[117]), .B(
        prince_inst_sbox_inst15_sh1_tmp[1]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[1]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk1_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[1]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk2_U1 ( .A(r[118]), .B(
        prince_inst_sbox_inst15_sh1_tmp[2]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[2]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk2_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[2]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk3_U1 ( .A(r[119]), .B(
        prince_inst_sbox_inst15_sh1_tmp[3]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[3]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk3_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[3]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk4_U1 ( .A(r[116]), .B(
        prince_inst_sbox_inst15_sh1_tmp[4]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[4]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk4_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[4]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk5_U1 ( .A(r[117]), .B(
        prince_inst_sbox_inst15_sh1_tmp[5]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[5]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk5_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[5]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk6_U1 ( .A(r[118]), .B(
        prince_inst_sbox_inst15_sh1_tmp[6]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[6]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk6_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[6]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_msk7_U1 ( .A(r[119]), .B(
        prince_inst_sbox_inst15_sh1_tmp[7]), .Z(
        prince_inst_sbox_inst15_c_inst1_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst1_y[7]), 
        .ZN(prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst1_msk7_xr), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst1_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst1_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst1_ax_U3 ( .A(
        prince_inst_sbox_inst15_c_inst1_ax_n6), .B(
        prince_inst_sbox_inst15_c_inst1_ax_n5), .ZN(prince_inst_sout_x[61]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst1_ax_U2 ( .A(
        prince_inst_sbox_inst15_c_inst1_y[1]), .B(
        prince_inst_sbox_inst15_c_inst1_y[0]), .ZN(
        prince_inst_sbox_inst15_c_inst1_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_ax_U1 ( .A(
        prince_inst_sbox_inst15_c_inst1_y[2]), .B(
        prince_inst_sbox_inst15_c_inst1_y[3]), .Z(
        prince_inst_sbox_inst15_c_inst1_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst1_ay_U3 ( .A(
        prince_inst_sbox_inst15_c_inst1_ay_n6), .B(
        prince_inst_sbox_inst15_c_inst1_ay_n5), .ZN(final_y[61]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst1_ay_U2 ( .A(
        prince_inst_sbox_inst15_c_inst1_y[5]), .B(
        prince_inst_sbox_inst15_c_inst1_y[4]), .ZN(
        prince_inst_sbox_inst15_c_inst1_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst1_ay_U1 ( .A(
        prince_inst_sbox_inst15_c_inst1_y[6]), .B(
        prince_inst_sbox_inst15_c_inst1_y[7]), .Z(
        prince_inst_sbox_inst15_c_inst1_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk0_U1 ( .A(r[120]), .B(
        prince_inst_sbox_inst15_sh2_tmp[0]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[0]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk0_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[0]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk1_U1 ( .A(r[121]), .B(
        prince_inst_sbox_inst15_sh2_tmp[1]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[1]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk1_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[1]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk2_U1 ( .A(r[122]), .B(
        prince_inst_sbox_inst15_sh2_tmp[2]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[2]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk2_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[2]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk3_U1 ( .A(r[123]), .B(
        prince_inst_sbox_inst15_sh2_tmp[3]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[3]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk3_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[3]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk4_U1 ( .A(r[120]), .B(
        prince_inst_sbox_inst15_sh2_tmp[4]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[4]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk4_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[4]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk5_U1 ( .A(r[121]), .B(
        prince_inst_sbox_inst15_sh2_tmp[5]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[5]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk5_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[5]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk6_U1 ( .A(r[122]), .B(
        prince_inst_sbox_inst15_sh2_tmp[6]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[6]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk6_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[6]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_msk7_U1 ( .A(r[123]), .B(
        prince_inst_sbox_inst15_sh2_tmp[7]), .Z(
        prince_inst_sbox_inst15_c_inst2_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst2_y[7]), 
        .ZN(prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst2_msk7_xr), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst2_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst2_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst2_ax_U3 ( .A(
        prince_inst_sbox_inst15_c_inst2_ax_n6), .B(
        prince_inst_sbox_inst15_c_inst2_ax_n5), .ZN(prince_inst_sout_x[62]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst2_ax_U2 ( .A(
        prince_inst_sbox_inst15_c_inst2_y[1]), .B(
        prince_inst_sbox_inst15_c_inst2_y[0]), .ZN(
        prince_inst_sbox_inst15_c_inst2_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_ax_U1 ( .A(
        prince_inst_sbox_inst15_c_inst2_y[2]), .B(
        prince_inst_sbox_inst15_c_inst2_y[3]), .Z(
        prince_inst_sbox_inst15_c_inst2_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst2_ay_U3 ( .A(
        prince_inst_sbox_inst15_c_inst2_ay_n6), .B(
        prince_inst_sbox_inst15_c_inst2_ay_n5), .ZN(final_y[62]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst2_ay_U2 ( .A(
        prince_inst_sbox_inst15_c_inst2_y[5]), .B(
        prince_inst_sbox_inst15_c_inst2_y[4]), .ZN(
        prince_inst_sbox_inst15_c_inst2_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst2_ay_U1 ( .A(
        prince_inst_sbox_inst15_c_inst2_y[6]), .B(
        prince_inst_sbox_inst15_c_inst2_y[7]), .Z(
        prince_inst_sbox_inst15_c_inst2_ay_n6) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk0_U1 ( .A(r[124]), .B(
        prince_inst_sbox_inst15_sh3_tmp[0]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk0_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[0]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk0_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk0_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[0]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk1_U1 ( .A(r[125]), .B(
        prince_inst_sbox_inst15_sh3_tmp[1]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk1_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[1]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk1_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk1_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[1]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk2_U1 ( .A(r[126]), .B(
        prince_inst_sbox_inst15_sh3_tmp[2]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk2_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[2]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk2_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk2_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[2]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk3_U1 ( .A(r[127]), .B(
        prince_inst_sbox_inst15_sh3_tmp[3]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk3_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[3]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk3_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk3_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[3]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk4_U1 ( .A(r[124]), .B(
        prince_inst_sbox_inst15_sh3_tmp[4]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk4_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[4]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk4_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk4_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[4]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk5_U1 ( .A(r[125]), .B(
        prince_inst_sbox_inst15_sh3_tmp[5]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk5_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[5]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk5_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk5_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[5]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk6_U1 ( .A(r[126]), .B(
        prince_inst_sbox_inst15_sh3_tmp[6]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk6_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[6]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk6_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk6_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[6]) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_msk7_U1 ( .A(r[127]), .B(
        prince_inst_sbox_inst15_sh3_tmp[7]), .Z(
        prince_inst_sbox_inst15_c_inst3_msk7_xr) );
  NOR3_X1 prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_U6 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n12), .A2(rst), .A3(
        prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n11), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n6) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_U5 ( .A1(
        prince_inst_sbox_inst15_n9), .A2(prince_inst_sbox_inst15_c_inst3_y[7]), 
        .ZN(prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n11) );
  NOR2_X1 prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_U4 ( .A1(
        prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n10), .A2(
        prince_inst_sbox_inst15_c_inst3_msk7_xr), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n12) );
  INV_X1 prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_U3 ( .A(
        prince_inst_sbox_inst15_n9), .ZN(
        prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n10) );
  DFF_X1 prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_s_current_state_reg ( .D(
        prince_inst_sbox_inst15_c_inst3_msk7_reg_xr_n6), .CK(clk), .Q(
        prince_inst_sbox_inst15_c_inst3_y[7]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst3_ax_U3 ( .A(
        prince_inst_sbox_inst15_c_inst3_ax_n6), .B(
        prince_inst_sbox_inst15_c_inst3_ax_n5), .ZN(prince_inst_sout_x[63]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst3_ax_U2 ( .A(
        prince_inst_sbox_inst15_c_inst3_y[1]), .B(
        prince_inst_sbox_inst15_c_inst3_y[0]), .ZN(
        prince_inst_sbox_inst15_c_inst3_ax_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_ax_U1 ( .A(
        prince_inst_sbox_inst15_c_inst3_y[2]), .B(
        prince_inst_sbox_inst15_c_inst3_y[3]), .Z(
        prince_inst_sbox_inst15_c_inst3_ax_n6) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst3_ay_U3 ( .A(
        prince_inst_sbox_inst15_c_inst3_ay_n6), .B(
        prince_inst_sbox_inst15_c_inst3_ay_n5), .ZN(final_y[63]) );
  XNOR2_X1 prince_inst_sbox_inst15_c_inst3_ay_U2 ( .A(
        prince_inst_sbox_inst15_c_inst3_y[5]), .B(
        prince_inst_sbox_inst15_c_inst3_y[4]), .ZN(
        prince_inst_sbox_inst15_c_inst3_ay_n5) );
  XOR2_X1 prince_inst_sbox_inst15_c_inst3_ay_U1 ( .A(
        prince_inst_sbox_inst15_c_inst3_y[6]), .B(
        prince_inst_sbox_inst15_c_inst3_y[7]), .Z(
        prince_inst_sbox_inst15_c_inst3_ay_n6) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a0_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a0_n1), .B(prince_inst_min_x[4]), .ZN(
        rout_x[0]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a0_U1 ( .A(prince_inst_min_x[0]), .B(
        prince_inst_min_x[8]), .ZN(prince_inst_mx_inst_m1_inst1_a0_n1) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a1_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a1_n3), .B(prince_inst_min_x[9]), .ZN(
        rout_x[1]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a1_U1 ( .A(prince_inst_min_x[5]), .B(
        prince_inst_min_x[13]), .ZN(prince_inst_mx_inst_m1_inst1_a1_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a2_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a2_n3), .B(prince_inst_min_x[10]), .ZN(
        rout_x[2]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a2_U1 ( .A(prince_inst_min_x[2]), .B(
        prince_inst_min_x[14]), .ZN(prince_inst_mx_inst_m1_inst1_a2_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a3_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a3_n3), .B(prince_inst_min_x[7]), .ZN(
        rout_x[3]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a3_U1 ( .A(prince_inst_min_x[3]), .B(
        prince_inst_min_x[15]), .ZN(prince_inst_mx_inst_m1_inst1_a3_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a4_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a4_n3), .B(prince_inst_min_x[4]), .ZN(
        rout_x[4]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a4_U1 ( .A(prince_inst_min_x[0]), .B(
        prince_inst_min_x[12]), .ZN(prince_inst_mx_inst_m1_inst1_a4_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a5_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a5_n3), .B(prince_inst_min_x[5]), .ZN(
        rout_x[5]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a5_U1 ( .A(prince_inst_min_x[1]), .B(
        prince_inst_min_x[9]), .ZN(prince_inst_mx_inst_m1_inst1_a5_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a6_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a6_n3), .B(prince_inst_min_x[10]), .ZN(
        rout_x[6]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a6_U1 ( .A(prince_inst_min_x[6]), .B(
        prince_inst_min_x[14]), .ZN(prince_inst_mx_inst_m1_inst1_a6_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a7_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a7_n3), .B(prince_inst_min_x[11]), .ZN(
        rout_x[7]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a7_U1 ( .A(prince_inst_min_x[3]), .B(
        prince_inst_min_x[15]), .ZN(prince_inst_mx_inst_m1_inst1_a7_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a8_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a8_n3), .B(prince_inst_min_x[8]), .ZN(
        rout_x[8]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a8_U1 ( .A(prince_inst_min_x[0]), .B(
        prince_inst_min_x[12]), .ZN(prince_inst_mx_inst_m1_inst1_a8_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a9_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a9_n3), .B(prince_inst_min_x[5]), .ZN(
        rout_x[9]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a9_U1 ( .A(prince_inst_min_x[1]), .B(
        prince_inst_min_x[13]), .ZN(prince_inst_mx_inst_m1_inst1_a9_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a10_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a10_n3), .B(prince_inst_min_x[6]), .ZN(
        rout_x[10]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a10_U1 ( .A(prince_inst_min_x[2]), .B(
        prince_inst_min_x[10]), .ZN(prince_inst_mx_inst_m1_inst1_a10_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a11_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a11_n3), .B(prince_inst_min_x[11]), .ZN(
        rout_x[11]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a11_U1 ( .A(prince_inst_min_x[7]), .B(
        prince_inst_min_x[15]), .ZN(prince_inst_mx_inst_m1_inst1_a11_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a12_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a12_n3), .B(prince_inst_min_x[8]), .ZN(
        rout_x[12]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a12_U1 ( .A(prince_inst_min_x[4]), .B(
        prince_inst_min_x[12]), .ZN(prince_inst_mx_inst_m1_inst1_a12_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a13_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a13_n3), .B(prince_inst_min_x[9]), .ZN(
        rout_x[13]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a13_U1 ( .A(prince_inst_min_x[1]), .B(
        prince_inst_min_x[13]), .ZN(prince_inst_mx_inst_m1_inst1_a13_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a14_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a14_n3), .B(prince_inst_min_x[6]), .ZN(
        rout_x[14]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a14_U1 ( .A(prince_inst_min_x[2]), .B(
        prince_inst_min_x[14]), .ZN(prince_inst_mx_inst_m1_inst1_a14_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a15_U2 ( .A(
        prince_inst_mx_inst_m1_inst1_a15_n3), .B(prince_inst_min_x[7]), .ZN(
        rout_x[15]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst1_a15_U1 ( .A(prince_inst_min_x[3]), .B(
        prince_inst_min_x[11]), .ZN(prince_inst_mx_inst_m1_inst1_a15_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a0_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a0_n3), .B(prince_inst_min_x[24]), .ZN(
        rout_x[16]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a0_U1 ( .A(prince_inst_min_x[20]), .B(
        prince_inst_min_x[28]), .ZN(prince_inst_mx_inst_m2_inst1_a0_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a1_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a1_n3), .B(prince_inst_min_x[25]), .ZN(
        rout_x[17]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a1_U1 ( .A(prince_inst_min_x[17]), .B(
        prince_inst_min_x[29]), .ZN(prince_inst_mx_inst_m2_inst1_a1_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a2_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a2_n3), .B(prince_inst_min_x[22]), .ZN(
        rout_x[18]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a2_U1 ( .A(prince_inst_min_x[18]), .B(
        prince_inst_min_x[30]), .ZN(prince_inst_mx_inst_m2_inst1_a2_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a3_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a3_n3), .B(prince_inst_min_x[23]), .ZN(
        rout_x[19]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a3_U1 ( .A(prince_inst_min_x[19]), .B(
        prince_inst_min_x[27]), .ZN(prince_inst_mx_inst_m2_inst1_a3_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a4_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a4_n3), .B(prince_inst_min_x[20]), .ZN(
        rout_x[20]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a4_U1 ( .A(prince_inst_min_x[16]), .B(
        prince_inst_min_x[24]), .ZN(prince_inst_mx_inst_m2_inst1_a4_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a5_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a5_n3), .B(prince_inst_min_x[25]), .ZN(
        rout_x[21]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a5_U1 ( .A(prince_inst_min_x[21]), .B(
        prince_inst_min_x[29]), .ZN(prince_inst_mx_inst_m2_inst1_a5_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a6_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a6_n3), .B(prince_inst_min_x[26]), .ZN(
        rout_x[22]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a6_U1 ( .A(prince_inst_min_x[18]), .B(
        prince_inst_min_x[30]), .ZN(prince_inst_mx_inst_m2_inst1_a6_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a7_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a7_n3), .B(prince_inst_min_x[23]), .ZN(
        rout_x[23]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a7_U1 ( .A(prince_inst_min_x[19]), .B(
        prince_inst_min_x[31]), .ZN(prince_inst_mx_inst_m2_inst1_a7_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a8_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a8_n3), .B(prince_inst_min_x[20]), .ZN(
        rout_x[24]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a8_U1 ( .A(prince_inst_min_x[16]), .B(
        prince_inst_min_x[28]), .ZN(prince_inst_mx_inst_m2_inst1_a8_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a9_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a9_n3), .B(prince_inst_min_x[21]), .ZN(
        rout_x[25]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a9_U1 ( .A(prince_inst_min_x[17]), .B(
        prince_inst_min_x[25]), .ZN(prince_inst_mx_inst_m2_inst1_a9_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a10_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a10_n3), .B(prince_inst_min_x[26]), .ZN(
        rout_x[26]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a10_U1 ( .A(prince_inst_min_x[22]), 
        .B(prince_inst_min_x[30]), .ZN(prince_inst_mx_inst_m2_inst1_a10_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a11_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a11_n3), .B(prince_inst_min_x[27]), .ZN(
        rout_x[27]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a11_U1 ( .A(prince_inst_min_x[19]), 
        .B(prince_inst_min_x[31]), .ZN(prince_inst_mx_inst_m2_inst1_a11_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a12_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a12_n3), .B(prince_inst_min_x[24]), .ZN(
        rout_x[28]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a12_U1 ( .A(prince_inst_min_x[16]), 
        .B(prince_inst_min_x[28]), .ZN(prince_inst_mx_inst_m2_inst1_a12_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a13_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a13_n3), .B(prince_inst_min_x[21]), .ZN(
        rout_x[29]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a13_U1 ( .A(prince_inst_min_x[17]), 
        .B(prince_inst_min_x[29]), .ZN(prince_inst_mx_inst_m2_inst1_a13_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a14_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a14_n3), .B(prince_inst_min_x[22]), .ZN(
        rout_x[30]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a14_U1 ( .A(prince_inst_min_x[18]), 
        .B(prince_inst_min_x[26]), .ZN(prince_inst_mx_inst_m2_inst1_a14_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a15_U2 ( .A(
        prince_inst_mx_inst_m2_inst1_a15_n3), .B(prince_inst_min_x[27]), .ZN(
        rout_x[31]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst1_a15_U1 ( .A(prince_inst_min_x[23]), 
        .B(prince_inst_min_x[31]), .ZN(prince_inst_mx_inst_m2_inst1_a15_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a0_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a0_n3), .B(prince_inst_min_x[40]), .ZN(
        rout_x[32]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a0_U1 ( .A(prince_inst_min_x[36]), .B(
        prince_inst_min_x[44]), .ZN(prince_inst_mx_inst_m2_inst2_a0_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a1_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a1_n3), .B(prince_inst_min_x[41]), .ZN(
        rout_x[33]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a1_U1 ( .A(prince_inst_min_x[33]), .B(
        prince_inst_min_x[45]), .ZN(prince_inst_mx_inst_m2_inst2_a1_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a2_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a2_n3), .B(prince_inst_min_x[38]), .ZN(
        rout_x[34]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a2_U1 ( .A(prince_inst_min_x[34]), .B(
        prince_inst_min_x[46]), .ZN(prince_inst_mx_inst_m2_inst2_a2_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a3_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a3_n3), .B(prince_inst_min_x[39]), .ZN(
        rout_x[35]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a3_U1 ( .A(prince_inst_min_x[35]), .B(
        prince_inst_min_x[43]), .ZN(prince_inst_mx_inst_m2_inst2_a3_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a4_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a4_n3), .B(prince_inst_min_x[36]), .ZN(
        rout_x[36]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a4_U1 ( .A(prince_inst_min_x[32]), .B(
        prince_inst_min_x[40]), .ZN(prince_inst_mx_inst_m2_inst2_a4_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a5_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a5_n3), .B(prince_inst_min_x[41]), .ZN(
        rout_x[37]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a5_U1 ( .A(prince_inst_min_x[37]), .B(
        prince_inst_min_x[45]), .ZN(prince_inst_mx_inst_m2_inst2_a5_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a6_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a6_n3), .B(prince_inst_min_x[42]), .ZN(
        rout_x[38]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a6_U1 ( .A(prince_inst_min_x[34]), .B(
        prince_inst_min_x[46]), .ZN(prince_inst_mx_inst_m2_inst2_a6_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a7_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a7_n3), .B(prince_inst_min_x[39]), .ZN(
        rout_x[39]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a7_U1 ( .A(prince_inst_min_x[35]), .B(
        prince_inst_min_x[47]), .ZN(prince_inst_mx_inst_m2_inst2_a7_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a8_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a8_n3), .B(prince_inst_min_x[36]), .ZN(
        rout_x[40]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a8_U1 ( .A(prince_inst_min_x[32]), .B(
        prince_inst_min_x[44]), .ZN(prince_inst_mx_inst_m2_inst2_a8_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a9_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a9_n3), .B(prince_inst_min_x[37]), .ZN(
        rout_x[41]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a9_U1 ( .A(prince_inst_min_x[33]), .B(
        prince_inst_min_x[41]), .ZN(prince_inst_mx_inst_m2_inst2_a9_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a10_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a10_n3), .B(prince_inst_min_x[42]), .ZN(
        rout_x[42]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a10_U1 ( .A(prince_inst_min_x[38]), 
        .B(prince_inst_min_x[46]), .ZN(prince_inst_mx_inst_m2_inst2_a10_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a11_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a11_n3), .B(prince_inst_min_x[43]), .ZN(
        rout_x[43]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a11_U1 ( .A(prince_inst_min_x[35]), 
        .B(prince_inst_min_x[47]), .ZN(prince_inst_mx_inst_m2_inst2_a11_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a12_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a12_n3), .B(prince_inst_min_x[40]), .ZN(
        rout_x[44]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a12_U1 ( .A(prince_inst_min_x[32]), 
        .B(prince_inst_min_x[44]), .ZN(prince_inst_mx_inst_m2_inst2_a12_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a13_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a13_n3), .B(prince_inst_min_x[37]), .ZN(
        rout_x[45]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a13_U1 ( .A(prince_inst_min_x[33]), 
        .B(prince_inst_min_x[45]), .ZN(prince_inst_mx_inst_m2_inst2_a13_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a14_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a14_n3), .B(prince_inst_min_x[38]), .ZN(
        rout_x[46]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a14_U1 ( .A(prince_inst_min_x[34]), 
        .B(prince_inst_min_x[42]), .ZN(prince_inst_mx_inst_m2_inst2_a14_n3) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a15_U2 ( .A(
        prince_inst_mx_inst_m2_inst2_a15_n3), .B(prince_inst_min_x[43]), .ZN(
        rout_x[47]) );
  XNOR2_X1 prince_inst_mx_inst_m2_inst2_a15_U1 ( .A(prince_inst_min_x[39]), 
        .B(prince_inst_min_x[47]), .ZN(prince_inst_mx_inst_m2_inst2_a15_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a0_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a0_n3), .B(prince_inst_min_x[52]), .ZN(
        rout_x[48]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a0_U1 ( .A(prince_inst_min_x[48]), .B(
        prince_inst_min_x[56]), .ZN(prince_inst_mx_inst_m1_inst2_a0_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a1_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a1_n3), .B(prince_inst_min_x[57]), .ZN(
        rout_x[49]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a1_U1 ( .A(prince_inst_min_x[53]), .B(
        prince_inst_min_x[61]), .ZN(prince_inst_mx_inst_m1_inst2_a1_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a2_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a2_n3), .B(prince_inst_min_x[58]), .ZN(
        rout_x[50]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a2_U1 ( .A(prince_inst_min_x[50]), .B(
        prince_inst_min_x[62]), .ZN(prince_inst_mx_inst_m1_inst2_a2_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a3_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a3_n3), .B(prince_inst_min_x[55]), .ZN(
        rout_x[51]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a3_U1 ( .A(prince_inst_min_x[51]), .B(
        prince_inst_min_x[63]), .ZN(prince_inst_mx_inst_m1_inst2_a3_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a4_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a4_n3), .B(prince_inst_min_x[52]), .ZN(
        rout_x[52]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a4_U1 ( .A(prince_inst_min_x[48]), .B(
        prince_inst_min_x[60]), .ZN(prince_inst_mx_inst_m1_inst2_a4_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a5_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a5_n3), .B(prince_inst_min_x[53]), .ZN(
        rout_x[53]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a5_U1 ( .A(prince_inst_min_x[49]), .B(
        prince_inst_min_x[57]), .ZN(prince_inst_mx_inst_m1_inst2_a5_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a6_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a6_n3), .B(prince_inst_min_x[58]), .ZN(
        rout_x[54]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a6_U1 ( .A(prince_inst_min_x[54]), .B(
        prince_inst_min_x[62]), .ZN(prince_inst_mx_inst_m1_inst2_a6_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a7_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a7_n3), .B(prince_inst_min_x[59]), .ZN(
        rout_x[55]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a7_U1 ( .A(prince_inst_min_x[51]), .B(
        prince_inst_min_x[63]), .ZN(prince_inst_mx_inst_m1_inst2_a7_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a8_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a8_n3), .B(prince_inst_min_x[56]), .ZN(
        rout_x[56]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a8_U1 ( .A(prince_inst_min_x[48]), .B(
        prince_inst_min_x[60]), .ZN(prince_inst_mx_inst_m1_inst2_a8_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a9_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a9_n3), .B(prince_inst_min_x[53]), .ZN(
        rout_x[57]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a9_U1 ( .A(prince_inst_min_x[49]), .B(
        prince_inst_min_x[61]), .ZN(prince_inst_mx_inst_m1_inst2_a9_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a10_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a10_n3), .B(prince_inst_min_x[54]), .ZN(
        rout_x[58]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a10_U1 ( .A(prince_inst_min_x[50]), 
        .B(prince_inst_min_x[58]), .ZN(prince_inst_mx_inst_m1_inst2_a10_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a11_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a11_n3), .B(prince_inst_min_x[59]), .ZN(
        rout_x[59]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a11_U1 ( .A(prince_inst_min_x[55]), 
        .B(prince_inst_min_x[63]), .ZN(prince_inst_mx_inst_m1_inst2_a11_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a12_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a12_n3), .B(prince_inst_min_x[56]), .ZN(
        rout_x[60]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a12_U1 ( .A(prince_inst_min_x[52]), 
        .B(prince_inst_min_x[60]), .ZN(prince_inst_mx_inst_m1_inst2_a12_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a13_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a13_n3), .B(prince_inst_min_x[57]), .ZN(
        rout_x[61]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a13_U1 ( .A(prince_inst_min_x[49]), 
        .B(prince_inst_min_x[61]), .ZN(prince_inst_mx_inst_m1_inst2_a13_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a14_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a14_n3), .B(prince_inst_min_x[54]), .ZN(
        rout_x[62]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a14_U1 ( .A(prince_inst_min_x[50]), 
        .B(prince_inst_min_x[62]), .ZN(prince_inst_mx_inst_m1_inst2_a14_n3) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a15_U2 ( .A(
        prince_inst_mx_inst_m1_inst2_a15_n3), .B(prince_inst_min_x[55]), .ZN(
        rout_x[63]) );
  XNOR2_X1 prince_inst_mx_inst_m1_inst2_a15_U1 ( .A(prince_inst_min_x[51]), 
        .B(prince_inst_min_x[59]), .ZN(prince_inst_mx_inst_m1_inst2_a15_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a0_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a0_n3), .B(prince_inst_min_y[4]), .ZN(
        rout_y[0]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a0_U1 ( .A(prince_inst_min_y[0]), .B(
        prince_inst_min_y[8]), .ZN(prince_inst_my_inst_m1_inst1_a0_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a1_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a1_n3), .B(prince_inst_min_y[9]), .ZN(
        rout_y[1]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a1_U1 ( .A(prince_inst_min_y[5]), .B(
        prince_inst_min_y[13]), .ZN(prince_inst_my_inst_m1_inst1_a1_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a2_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a2_n3), .B(prince_inst_min_y[10]), .ZN(
        rout_y[2]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a2_U1 ( .A(prince_inst_min_y[2]), .B(
        prince_inst_min_y[14]), .ZN(prince_inst_my_inst_m1_inst1_a2_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a3_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a3_n3), .B(prince_inst_min_y[7]), .ZN(
        rout_y[3]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a3_U1 ( .A(prince_inst_min_y[3]), .B(
        prince_inst_min_y[15]), .ZN(prince_inst_my_inst_m1_inst1_a3_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a4_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a4_n3), .B(prince_inst_min_y[4]), .ZN(
        rout_y[4]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a4_U1 ( .A(prince_inst_min_y[0]), .B(
        prince_inst_min_y[12]), .ZN(prince_inst_my_inst_m1_inst1_a4_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a5_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a5_n3), .B(prince_inst_min_y[5]), .ZN(
        rout_y[5]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a5_U1 ( .A(prince_inst_min_y[1]), .B(
        prince_inst_min_y[9]), .ZN(prince_inst_my_inst_m1_inst1_a5_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a6_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a6_n3), .B(prince_inst_min_y[10]), .ZN(
        rout_y[6]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a6_U1 ( .A(prince_inst_min_y[6]), .B(
        prince_inst_min_y[14]), .ZN(prince_inst_my_inst_m1_inst1_a6_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a7_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a7_n3), .B(prince_inst_min_y[11]), .ZN(
        rout_y[7]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a7_U1 ( .A(prince_inst_min_y[3]), .B(
        prince_inst_min_y[15]), .ZN(prince_inst_my_inst_m1_inst1_a7_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a8_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a8_n3), .B(prince_inst_min_y[8]), .ZN(
        rout_y[8]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a8_U1 ( .A(prince_inst_min_y[0]), .B(
        prince_inst_min_y[12]), .ZN(prince_inst_my_inst_m1_inst1_a8_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a9_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a9_n3), .B(prince_inst_min_y[5]), .ZN(
        rout_y[9]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a9_U1 ( .A(prince_inst_min_y[1]), .B(
        prince_inst_min_y[13]), .ZN(prince_inst_my_inst_m1_inst1_a9_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a10_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a10_n3), .B(prince_inst_min_y[6]), .ZN(
        rout_y[10]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a10_U1 ( .A(prince_inst_min_y[2]), .B(
        prince_inst_min_y[10]), .ZN(prince_inst_my_inst_m1_inst1_a10_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a11_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a11_n3), .B(prince_inst_min_y[11]), .ZN(
        rout_y[11]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a11_U1 ( .A(prince_inst_min_y[7]), .B(
        prince_inst_min_y[15]), .ZN(prince_inst_my_inst_m1_inst1_a11_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a12_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a12_n3), .B(prince_inst_min_y[8]), .ZN(
        rout_y[12]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a12_U1 ( .A(prince_inst_min_y[4]), .B(
        prince_inst_min_y[12]), .ZN(prince_inst_my_inst_m1_inst1_a12_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a13_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a13_n3), .B(prince_inst_min_y[9]), .ZN(
        rout_y[13]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a13_U1 ( .A(prince_inst_min_y[1]), .B(
        prince_inst_min_y[13]), .ZN(prince_inst_my_inst_m1_inst1_a13_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a14_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a14_n3), .B(prince_inst_min_y[6]), .ZN(
        rout_y[14]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a14_U1 ( .A(prince_inst_min_y[2]), .B(
        prince_inst_min_y[14]), .ZN(prince_inst_my_inst_m1_inst1_a14_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a15_U2 ( .A(
        prince_inst_my_inst_m1_inst1_a15_n3), .B(prince_inst_min_y[7]), .ZN(
        rout_y[15]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst1_a15_U1 ( .A(prince_inst_min_y[3]), .B(
        prince_inst_min_y[11]), .ZN(prince_inst_my_inst_m1_inst1_a15_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a0_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a0_n3), .B(prince_inst_min_y[24]), .ZN(
        rout_y[16]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a0_U1 ( .A(prince_inst_min_y[20]), .B(
        prince_inst_min_y[28]), .ZN(prince_inst_my_inst_m2_inst1_a0_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a1_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a1_n3), .B(prince_inst_min_y[25]), .ZN(
        rout_y[17]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a1_U1 ( .A(prince_inst_min_y[17]), .B(
        prince_inst_min_y[29]), .ZN(prince_inst_my_inst_m2_inst1_a1_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a2_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a2_n3), .B(prince_inst_min_y[22]), .ZN(
        rout_y[18]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a2_U1 ( .A(prince_inst_min_y[18]), .B(
        prince_inst_min_y[30]), .ZN(prince_inst_my_inst_m2_inst1_a2_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a3_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a3_n3), .B(prince_inst_min_y[23]), .ZN(
        rout_y[19]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a3_U1 ( .A(prince_inst_min_y[19]), .B(
        prince_inst_min_y[27]), .ZN(prince_inst_my_inst_m2_inst1_a3_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a4_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a4_n3), .B(prince_inst_min_y[20]), .ZN(
        rout_y[20]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a4_U1 ( .A(prince_inst_min_y[16]), .B(
        prince_inst_min_y[24]), .ZN(prince_inst_my_inst_m2_inst1_a4_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a5_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a5_n3), .B(prince_inst_min_y[25]), .ZN(
        rout_y[21]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a5_U1 ( .A(prince_inst_min_y[21]), .B(
        prince_inst_min_y[29]), .ZN(prince_inst_my_inst_m2_inst1_a5_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a6_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a6_n3), .B(prince_inst_min_y[26]), .ZN(
        rout_y[22]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a6_U1 ( .A(prince_inst_min_y[18]), .B(
        prince_inst_min_y[30]), .ZN(prince_inst_my_inst_m2_inst1_a6_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a7_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a7_n3), .B(prince_inst_min_y[23]), .ZN(
        rout_y[23]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a7_U1 ( .A(prince_inst_min_y[19]), .B(
        prince_inst_min_y[31]), .ZN(prince_inst_my_inst_m2_inst1_a7_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a8_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a8_n3), .B(prince_inst_min_y[20]), .ZN(
        rout_y[24]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a8_U1 ( .A(prince_inst_min_y[16]), .B(
        prince_inst_min_y[28]), .ZN(prince_inst_my_inst_m2_inst1_a8_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a9_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a9_n3), .B(prince_inst_min_y[21]), .ZN(
        rout_y[25]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a9_U1 ( .A(prince_inst_min_y[17]), .B(
        prince_inst_min_y[25]), .ZN(prince_inst_my_inst_m2_inst1_a9_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a10_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a10_n3), .B(prince_inst_min_y[26]), .ZN(
        rout_y[26]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a10_U1 ( .A(prince_inst_min_y[22]), 
        .B(prince_inst_min_y[30]), .ZN(prince_inst_my_inst_m2_inst1_a10_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a11_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a11_n3), .B(prince_inst_min_y[27]), .ZN(
        rout_y[27]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a11_U1 ( .A(prince_inst_min_y[19]), 
        .B(prince_inst_min_y[31]), .ZN(prince_inst_my_inst_m2_inst1_a11_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a12_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a12_n3), .B(prince_inst_min_y[24]), .ZN(
        rout_y[28]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a12_U1 ( .A(prince_inst_min_y[16]), 
        .B(prince_inst_min_y[28]), .ZN(prince_inst_my_inst_m2_inst1_a12_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a13_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a13_n3), .B(prince_inst_min_y[21]), .ZN(
        rout_y[29]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a13_U1 ( .A(prince_inst_min_y[17]), 
        .B(prince_inst_min_y[29]), .ZN(prince_inst_my_inst_m2_inst1_a13_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a14_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a14_n3), .B(prince_inst_min_y[22]), .ZN(
        rout_y[30]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a14_U1 ( .A(prince_inst_min_y[18]), 
        .B(prince_inst_min_y[26]), .ZN(prince_inst_my_inst_m2_inst1_a14_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a15_U2 ( .A(
        prince_inst_my_inst_m2_inst1_a15_n3), .B(prince_inst_min_y[27]), .ZN(
        rout_y[31]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst1_a15_U1 ( .A(prince_inst_min_y[23]), 
        .B(prince_inst_min_y[31]), .ZN(prince_inst_my_inst_m2_inst1_a15_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a0_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a0_n3), .B(prince_inst_min_y[40]), .ZN(
        rout_y[32]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a0_U1 ( .A(prince_inst_min_y[36]), .B(
        prince_inst_min_y[44]), .ZN(prince_inst_my_inst_m2_inst2_a0_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a1_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a1_n3), .B(prince_inst_min_y[41]), .ZN(
        rout_y[33]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a1_U1 ( .A(prince_inst_min_y[33]), .B(
        prince_inst_min_y[45]), .ZN(prince_inst_my_inst_m2_inst2_a1_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a2_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a2_n3), .B(prince_inst_min_y[38]), .ZN(
        rout_y[34]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a2_U1 ( .A(prince_inst_min_y[34]), .B(
        prince_inst_min_y[46]), .ZN(prince_inst_my_inst_m2_inst2_a2_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a3_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a3_n3), .B(prince_inst_min_y[39]), .ZN(
        rout_y[35]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a3_U1 ( .A(prince_inst_min_y[35]), .B(
        prince_inst_min_y[43]), .ZN(prince_inst_my_inst_m2_inst2_a3_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a4_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a4_n3), .B(prince_inst_min_y[36]), .ZN(
        rout_y[36]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a4_U1 ( .A(prince_inst_min_y[32]), .B(
        prince_inst_min_y[40]), .ZN(prince_inst_my_inst_m2_inst2_a4_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a5_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a5_n3), .B(prince_inst_min_y[41]), .ZN(
        rout_y[37]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a5_U1 ( .A(prince_inst_min_y[37]), .B(
        prince_inst_min_y[45]), .ZN(prince_inst_my_inst_m2_inst2_a5_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a6_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a6_n3), .B(prince_inst_min_y[42]), .ZN(
        rout_y[38]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a6_U1 ( .A(prince_inst_min_y[34]), .B(
        prince_inst_min_y[46]), .ZN(prince_inst_my_inst_m2_inst2_a6_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a7_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a7_n3), .B(prince_inst_min_y[39]), .ZN(
        rout_y[39]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a7_U1 ( .A(prince_inst_min_y[35]), .B(
        prince_inst_min_y[47]), .ZN(prince_inst_my_inst_m2_inst2_a7_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a8_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a8_n3), .B(prince_inst_min_y[36]), .ZN(
        rout_y[40]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a8_U1 ( .A(prince_inst_min_y[32]), .B(
        prince_inst_min_y[44]), .ZN(prince_inst_my_inst_m2_inst2_a8_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a9_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a9_n3), .B(prince_inst_min_y[37]), .ZN(
        rout_y[41]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a9_U1 ( .A(prince_inst_min_y[33]), .B(
        prince_inst_min_y[41]), .ZN(prince_inst_my_inst_m2_inst2_a9_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a10_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a10_n3), .B(prince_inst_min_y[42]), .ZN(
        rout_y[42]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a10_U1 ( .A(prince_inst_min_y[38]), 
        .B(prince_inst_min_y[46]), .ZN(prince_inst_my_inst_m2_inst2_a10_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a11_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a11_n3), .B(prince_inst_min_y[43]), .ZN(
        rout_y[43]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a11_U1 ( .A(prince_inst_min_y[35]), 
        .B(prince_inst_min_y[47]), .ZN(prince_inst_my_inst_m2_inst2_a11_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a12_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a12_n3), .B(prince_inst_min_y[40]), .ZN(
        rout_y[44]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a12_U1 ( .A(prince_inst_min_y[32]), 
        .B(prince_inst_min_y[44]), .ZN(prince_inst_my_inst_m2_inst2_a12_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a13_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a13_n3), .B(prince_inst_min_y[37]), .ZN(
        rout_y[45]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a13_U1 ( .A(prince_inst_min_y[33]), 
        .B(prince_inst_min_y[45]), .ZN(prince_inst_my_inst_m2_inst2_a13_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a14_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a14_n3), .B(prince_inst_min_y[38]), .ZN(
        rout_y[46]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a14_U1 ( .A(prince_inst_min_y[34]), 
        .B(prince_inst_min_y[42]), .ZN(prince_inst_my_inst_m2_inst2_a14_n3) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a15_U2 ( .A(
        prince_inst_my_inst_m2_inst2_a15_n3), .B(prince_inst_min_y[43]), .ZN(
        rout_y[47]) );
  XNOR2_X1 prince_inst_my_inst_m2_inst2_a15_U1 ( .A(prince_inst_min_y[39]), 
        .B(prince_inst_min_y[47]), .ZN(prince_inst_my_inst_m2_inst2_a15_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a0_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a0_n3), .B(prince_inst_min_y[52]), .ZN(
        rout_y[48]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a0_U1 ( .A(prince_inst_min_y[48]), .B(
        prince_inst_min_y[56]), .ZN(prince_inst_my_inst_m1_inst2_a0_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a1_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a1_n3), .B(prince_inst_min_y[57]), .ZN(
        rout_y[49]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a1_U1 ( .A(prince_inst_min_y[53]), .B(
        prince_inst_min_y[61]), .ZN(prince_inst_my_inst_m1_inst2_a1_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a2_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a2_n3), .B(prince_inst_min_y[58]), .ZN(
        rout_y[50]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a2_U1 ( .A(prince_inst_min_y[50]), .B(
        prince_inst_min_y[62]), .ZN(prince_inst_my_inst_m1_inst2_a2_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a3_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a3_n3), .B(prince_inst_min_y[55]), .ZN(
        rout_y[51]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a3_U1 ( .A(prince_inst_min_y[51]), .B(
        prince_inst_min_y[63]), .ZN(prince_inst_my_inst_m1_inst2_a3_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a4_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a4_n3), .B(prince_inst_min_y[52]), .ZN(
        rout_y[52]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a4_U1 ( .A(prince_inst_min_y[48]), .B(
        prince_inst_min_y[60]), .ZN(prince_inst_my_inst_m1_inst2_a4_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a5_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a5_n3), .B(prince_inst_min_y[53]), .ZN(
        rout_y[53]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a5_U1 ( .A(prince_inst_min_y[49]), .B(
        prince_inst_min_y[57]), .ZN(prince_inst_my_inst_m1_inst2_a5_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a6_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a6_n3), .B(prince_inst_min_y[58]), .ZN(
        rout_y[54]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a6_U1 ( .A(prince_inst_min_y[54]), .B(
        prince_inst_min_y[62]), .ZN(prince_inst_my_inst_m1_inst2_a6_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a7_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a7_n3), .B(prince_inst_min_y[59]), .ZN(
        rout_y[55]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a7_U1 ( .A(prince_inst_min_y[51]), .B(
        prince_inst_min_y[63]), .ZN(prince_inst_my_inst_m1_inst2_a7_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a8_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a8_n3), .B(prince_inst_min_y[56]), .ZN(
        rout_y[56]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a8_U1 ( .A(prince_inst_min_y[48]), .B(
        prince_inst_min_y[60]), .ZN(prince_inst_my_inst_m1_inst2_a8_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a9_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a9_n3), .B(prince_inst_min_y[53]), .ZN(
        rout_y[57]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a9_U1 ( .A(prince_inst_min_y[49]), .B(
        prince_inst_min_y[61]), .ZN(prince_inst_my_inst_m1_inst2_a9_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a10_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a10_n3), .B(prince_inst_min_y[54]), .ZN(
        rout_y[58]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a10_U1 ( .A(prince_inst_min_y[50]), 
        .B(prince_inst_min_y[58]), .ZN(prince_inst_my_inst_m1_inst2_a10_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a11_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a11_n3), .B(prince_inst_min_y[59]), .ZN(
        rout_y[59]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a11_U1 ( .A(prince_inst_min_y[55]), 
        .B(prince_inst_min_y[63]), .ZN(prince_inst_my_inst_m1_inst2_a11_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a12_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a12_n3), .B(prince_inst_min_y[56]), .ZN(
        rout_y[60]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a12_U1 ( .A(prince_inst_min_y[52]), 
        .B(prince_inst_min_y[60]), .ZN(prince_inst_my_inst_m1_inst2_a12_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a13_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a13_n3), .B(prince_inst_min_y[57]), .ZN(
        rout_y[61]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a13_U1 ( .A(prince_inst_min_y[49]), 
        .B(prince_inst_min_y[61]), .ZN(prince_inst_my_inst_m1_inst2_a13_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a14_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a14_n3), .B(prince_inst_min_y[54]), .ZN(
        rout_y[62]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a14_U1 ( .A(prince_inst_min_y[50]), 
        .B(prince_inst_min_y[62]), .ZN(prince_inst_my_inst_m1_inst2_a14_n3) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a15_U2 ( .A(
        prince_inst_my_inst_m1_inst2_a15_n3), .B(prince_inst_min_y[55]), .ZN(
        rout_y[63]) );
  XNOR2_X1 prince_inst_my_inst_m1_inst2_a15_U1 ( .A(prince_inst_min_y[51]), 
        .B(prince_inst_min_y[59]), .ZN(prince_inst_my_inst_m1_inst2_a15_n3) );
  AND2_X1 mux_c0_U67 ( .A1(mux_c0_n265), .A2(final_x_k[59]), .ZN(c0[59]) );
  AND2_X1 mux_c0_U66 ( .A1(done), .A2(final_x_k[49]), .ZN(c0[49]) );
  AND2_X1 mux_c0_U65 ( .A1(mux_c0_n265), .A2(final_x_k[57]), .ZN(c0[57]) );
  AND2_X1 mux_c0_U64 ( .A1(done), .A2(final_x_k[41]), .ZN(c0[41]) );
  AND2_X1 mux_c0_U63 ( .A1(mux_c0_n265), .A2(final_x_k[55]), .ZN(c0[55]) );
  AND2_X1 mux_c0_U62 ( .A1(mux_c0_n265), .A2(final_x_k[60]), .ZN(c0[60]) );
  AND2_X1 mux_c0_U61 ( .A1(done), .A2(final_x_k[52]), .ZN(c0[52]) );
  AND2_X1 mux_c0_U60 ( .A1(mux_c0_n265), .A2(final_x_k[58]), .ZN(c0[58]) );
  AND2_X1 mux_c0_U59 ( .A1(mux_c0_n264), .A2(final_x_k[44]), .ZN(c0[44]) );
  AND2_X1 mux_c0_U58 ( .A1(done), .A2(final_x_k[36]), .ZN(c0[36]) );
  AND2_X1 mux_c0_U57 ( .A1(mux_c0_n265), .A2(final_x_k[45]), .ZN(c0[45]) );
  AND2_X1 mux_c0_U56 ( .A1(mux_c0_n264), .A2(final_x_k[34]), .ZN(c0[34]) );
  AND2_X1 mux_c0_U55 ( .A1(mux_c0_n265), .A2(final_x_k[48]), .ZN(c0[48]) );
  AND2_X1 mux_c0_U54 ( .A1(mux_c0_n265), .A2(final_x_k[61]), .ZN(c0[61]) );
  AND2_X1 mux_c0_U53 ( .A1(mux_c0_n264), .A2(final_x_k[32]), .ZN(c0[32]) );
  AND2_X1 mux_c0_U52 ( .A1(done), .A2(final_x_k[42]), .ZN(c0[42]) );
  AND2_X1 mux_c0_U51 ( .A1(mux_c0_n265), .A2(final_x_k[29]), .ZN(c0[29]) );
  AND2_X1 mux_c0_U50 ( .A1(mux_c0_n264), .A2(final_x_k[31]), .ZN(c0[31]) );
  AND2_X1 mux_c0_U49 ( .A1(done), .A2(final_x_k[53]), .ZN(c0[53]) );
  AND2_X1 mux_c0_U48 ( .A1(mux_c0_n265), .A2(final_x_k[26]), .ZN(c0[26]) );
  AND2_X1 mux_c0_U47 ( .A1(mux_c0_n265), .A2(final_x_k[43]), .ZN(c0[43]) );
  AND2_X1 mux_c0_U46 ( .A1(mux_c0_n265), .A2(final_x_k[56]), .ZN(c0[56]) );
  AND2_X1 mux_c0_U45 ( .A1(mux_c0_n264), .A2(final_x_k[25]), .ZN(c0[25]) );
  AND2_X1 mux_c0_U44 ( .A1(mux_c0_n265), .A2(final_x_k[35]), .ZN(c0[35]) );
  AND2_X1 mux_c0_U43 ( .A1(mux_c0_n265), .A2(final_x_k[37]), .ZN(c0[37]) );
  AND2_X1 mux_c0_U42 ( .A1(done), .A2(final_x_k[54]), .ZN(c0[54]) );
  AND2_X1 mux_c0_U41 ( .A1(mux_c0_n265), .A2(final_x_k[27]), .ZN(c0[27]) );
  AND2_X1 mux_c0_U40 ( .A1(mux_c0_n265), .A2(final_x_k[23]), .ZN(c0[23]) );
  AND2_X1 mux_c0_U39 ( .A1(mux_c0_n265), .A2(final_x_k[33]), .ZN(c0[33]) );
  AND2_X1 mux_c0_U38 ( .A1(done), .A2(final_x_k[51]), .ZN(c0[51]) );
  AND2_X1 mux_c0_U37 ( .A1(mux_c0_n265), .A2(final_x_k[50]), .ZN(c0[50]) );
  AND2_X1 mux_c0_U36 ( .A1(mux_c0_n264), .A2(final_x_k[22]), .ZN(c0[22]) );
  AND2_X1 mux_c0_U35 ( .A1(mux_c0_n265), .A2(final_x_k[21]), .ZN(c0[21]) );
  AND2_X1 mux_c0_U34 ( .A1(mux_c0_n264), .A2(final_x_k[20]), .ZN(c0[20]) );
  AND2_X1 mux_c0_U33 ( .A1(mux_c0_n264), .A2(final_x_k[24]), .ZN(c0[24]) );
  AND2_X1 mux_c0_U32 ( .A1(done), .A2(final_x_k[47]), .ZN(c0[47]) );
  AND2_X1 mux_c0_U31 ( .A1(mux_c0_n264), .A2(final_x_k[28]), .ZN(c0[28]) );
  AND2_X1 mux_c0_U30 ( .A1(mux_c0_n265), .A2(final_x_k[19]), .ZN(c0[19]) );
  AND2_X1 mux_c0_U29 ( .A1(mux_c0_n264), .A2(final_x_k[18]), .ZN(c0[18]) );
  AND2_X1 mux_c0_U28 ( .A1(mux_c0_n265), .A2(final_x_k[17]), .ZN(c0[17]) );
  AND2_X1 mux_c0_U27 ( .A1(mux_c0_n264), .A2(final_x_k[16]), .ZN(c0[16]) );
  AND2_X1 mux_c0_U26 ( .A1(mux_c0_n265), .A2(final_x_k[15]), .ZN(c0[15]) );
  AND2_X1 mux_c0_U25 ( .A1(mux_c0_n264), .A2(final_x_k[14]), .ZN(c0[14]) );
  AND2_X1 mux_c0_U24 ( .A1(mux_c0_n265), .A2(final_x_k[13]), .ZN(c0[13]) );
  AND2_X1 mux_c0_U23 ( .A1(mux_c0_n265), .A2(final_x_k[40]), .ZN(c0[40]) );
  AND2_X1 mux_c0_U22 ( .A1(mux_c0_n264), .A2(final_x_k[39]), .ZN(c0[39]) );
  AND2_X1 mux_c0_U21 ( .A1(mux_c0_n264), .A2(final_x_k[38]), .ZN(c0[38]) );
  AND2_X1 mux_c0_U20 ( .A1(mux_c0_n264), .A2(final_x_k[12]), .ZN(c0[12]) );
  AND2_X1 mux_c0_U19 ( .A1(mux_c0_n265), .A2(final_x_k[11]), .ZN(c0[11]) );
  AND2_X1 mux_c0_U18 ( .A1(mux_c0_n264), .A2(final_x_k[10]), .ZN(c0[10]) );
  AND2_X1 mux_c0_U17 ( .A1(mux_c0_n264), .A2(final_x_k[9]), .ZN(c0[9]) );
  AND2_X1 mux_c0_U16 ( .A1(mux_c0_n264), .A2(final_x_k[8]), .ZN(c0[8]) );
  AND2_X1 mux_c0_U15 ( .A1(mux_c0_n264), .A2(final_x_k[7]), .ZN(c0[7]) );
  AND2_X1 mux_c0_U14 ( .A1(done), .A2(final_x_k[30]), .ZN(c0[30]) );
  AND2_X1 mux_c0_U13 ( .A1(mux_c0_n264), .A2(final_x_k[6]), .ZN(c0[6]) );
  AND2_X1 mux_c0_U12 ( .A1(done), .A2(final_x_k[46]), .ZN(c0[46]) );
  AND2_X1 mux_c0_U11 ( .A1(mux_c0_n264), .A2(final_x_k[5]), .ZN(c0[5]) );
  AND2_X1 mux_c0_U10 ( .A1(mux_c0_n264), .A2(final_x_k[4]), .ZN(c0[4]) );
  AND2_X1 mux_c0_U9 ( .A1(mux_c0_n265), .A2(final_x_k[62]), .ZN(c0[62]) );
  AND2_X1 mux_c0_U8 ( .A1(mux_c0_n264), .A2(final_x_k[3]), .ZN(c0[3]) );
  AND2_X1 mux_c0_U7 ( .A1(mux_c0_n264), .A2(final_x_k[2]), .ZN(c0[2]) );
  AND2_X1 mux_c0_U6 ( .A1(mux_c0_n264), .A2(final_x_k[1]), .ZN(c0[1]) );
  AND2_X1 mux_c0_U5 ( .A1(mux_c0_n264), .A2(final_x_k[0]), .ZN(c0[0]) );
  AND2_X1 mux_c0_U4 ( .A1(mux_c0_n265), .A2(final_x_k[63]), .ZN(c0[63]) );
  INV_X1 mux_c0_U3 ( .A(mux_c0_n263), .ZN(mux_c0_n265) );
  INV_X1 mux_c0_U2 ( .A(mux_c0_n263), .ZN(mux_c0_n264) );
  INV_X1 mux_c0_U1 ( .A(done), .ZN(mux_c0_n263) );
  AND2_X1 mux_c1_U67 ( .A1(mux_c1_n264), .A2(final_y[63]), .ZN(c1[63]) );
  AND2_X1 mux_c1_U66 ( .A1(mux_c1_n264), .A2(final_y[62]), .ZN(c1[62]) );
  AND2_X1 mux_c1_U65 ( .A1(mux_c1_n264), .A2(final_y[61]), .ZN(c1[61]) );
  AND2_X1 mux_c1_U64 ( .A1(mux_c1_n264), .A2(final_y[60]), .ZN(c1[60]) );
  AND2_X1 mux_c1_U63 ( .A1(mux_c1_n264), .A2(final_y[59]), .ZN(c1[59]) );
  AND2_X1 mux_c1_U62 ( .A1(mux_c1_n264), .A2(final_y[58]), .ZN(c1[58]) );
  AND2_X1 mux_c1_U61 ( .A1(mux_c1_n264), .A2(final_y[57]), .ZN(c1[57]) );
  AND2_X1 mux_c1_U60 ( .A1(mux_c1_n264), .A2(final_y[56]), .ZN(c1[56]) );
  AND2_X1 mux_c1_U59 ( .A1(mux_c1_n264), .A2(final_y[55]), .ZN(c1[55]) );
  AND2_X1 mux_c1_U58 ( .A1(mux_c1_n263), .A2(final_y[54]), .ZN(c1[54]) );
  AND2_X1 mux_c1_U57 ( .A1(mux_c1_n264), .A2(final_y[53]), .ZN(c1[53]) );
  AND2_X1 mux_c1_U56 ( .A1(mux_c1_n263), .A2(final_y[52]), .ZN(c1[52]) );
  AND2_X1 mux_c1_U55 ( .A1(mux_c1_n264), .A2(final_y[51]), .ZN(c1[51]) );
  AND2_X1 mux_c1_U54 ( .A1(mux_c1_n263), .A2(final_y[50]), .ZN(c1[50]) );
  AND2_X1 mux_c1_U53 ( .A1(mux_c1_n264), .A2(final_y[49]), .ZN(c1[49]) );
  AND2_X1 mux_c1_U52 ( .A1(mux_c1_n263), .A2(final_y[48]), .ZN(c1[48]) );
  AND2_X1 mux_c1_U51 ( .A1(mux_c1_n264), .A2(final_y[47]), .ZN(c1[47]) );
  AND2_X1 mux_c1_U50 ( .A1(mux_c1_n263), .A2(final_y[46]), .ZN(c1[46]) );
  AND2_X1 mux_c1_U49 ( .A1(mux_c1_n264), .A2(final_y[45]), .ZN(c1[45]) );
  AND2_X1 mux_c1_U48 ( .A1(mux_c1_n263), .A2(final_y[44]), .ZN(c1[44]) );
  AND2_X1 mux_c1_U47 ( .A1(mux_c1_n263), .A2(final_y[43]), .ZN(c1[43]) );
  AND2_X1 mux_c1_U46 ( .A1(mux_c1_n263), .A2(final_y[42]), .ZN(c1[42]) );
  AND2_X1 mux_c1_U45 ( .A1(mux_c1_n263), .A2(final_y[41]), .ZN(c1[41]) );
  AND2_X1 mux_c1_U44 ( .A1(mux_c1_n263), .A2(final_y[40]), .ZN(c1[40]) );
  AND2_X1 mux_c1_U43 ( .A1(mux_c1_n263), .A2(final_y[39]), .ZN(c1[39]) );
  AND2_X1 mux_c1_U42 ( .A1(mux_c1_n263), .A2(final_y[38]), .ZN(c1[38]) );
  AND2_X1 mux_c1_U41 ( .A1(mux_c1_n263), .A2(final_y[37]), .ZN(c1[37]) );
  AND2_X1 mux_c1_U40 ( .A1(mux_c1_n263), .A2(final_y[36]), .ZN(c1[36]) );
  AND2_X1 mux_c1_U39 ( .A1(mux_c1_n263), .A2(final_y[35]), .ZN(c1[35]) );
  AND2_X1 mux_c1_U38 ( .A1(mux_c1_n263), .A2(final_y[34]), .ZN(c1[34]) );
  AND2_X1 mux_c1_U37 ( .A1(mux_c1_n263), .A2(final_y[33]), .ZN(c1[33]) );
  AND2_X1 mux_c1_U36 ( .A1(mux_c1_n264), .A2(final_y[32]), .ZN(c1[32]) );
  AND2_X1 mux_c1_U35 ( .A1(mux_c1_n264), .A2(final_y[31]), .ZN(c1[31]) );
  AND2_X1 mux_c1_U34 ( .A1(mux_c1_n264), .A2(final_y[30]), .ZN(c1[30]) );
  AND2_X1 mux_c1_U33 ( .A1(mux_c1_n263), .A2(final_y[29]), .ZN(c1[29]) );
  AND2_X1 mux_c1_U32 ( .A1(mux_c1_n263), .A2(final_y[28]), .ZN(c1[28]) );
  AND2_X1 mux_c1_U31 ( .A1(mux_c1_n264), .A2(final_y[27]), .ZN(c1[27]) );
  AND2_X1 mux_c1_U30 ( .A1(mux_c1_n264), .A2(final_y[26]), .ZN(c1[26]) );
  AND2_X1 mux_c1_U29 ( .A1(mux_c1_n264), .A2(final_y[25]), .ZN(c1[25]) );
  AND2_X1 mux_c1_U28 ( .A1(mux_c1_n263), .A2(final_y[24]), .ZN(c1[24]) );
  AND2_X1 mux_c1_U27 ( .A1(mux_c1_n264), .A2(final_y[23]), .ZN(c1[23]) );
  AND2_X1 mux_c1_U26 ( .A1(mux_c1_n263), .A2(final_y[22]), .ZN(c1[22]) );
  AND2_X1 mux_c1_U25 ( .A1(mux_c1_n263), .A2(final_y[21]), .ZN(c1[21]) );
  AND2_X1 mux_c1_U24 ( .A1(mux_c1_n263), .A2(final_y[20]), .ZN(c1[20]) );
  AND2_X1 mux_c1_U23 ( .A1(mux_c1_n264), .A2(final_y[19]), .ZN(c1[19]) );
  AND2_X1 mux_c1_U22 ( .A1(mux_c1_n264), .A2(final_y[18]), .ZN(c1[18]) );
  AND2_X1 mux_c1_U21 ( .A1(mux_c1_n263), .A2(final_y[17]), .ZN(c1[17]) );
  AND2_X1 mux_c1_U20 ( .A1(mux_c1_n263), .A2(final_y[16]), .ZN(c1[16]) );
  AND2_X1 mux_c1_U19 ( .A1(mux_c1_n264), .A2(final_y[15]), .ZN(c1[15]) );
  AND2_X1 mux_c1_U18 ( .A1(mux_c1_n264), .A2(final_y[14]), .ZN(c1[14]) );
  AND2_X1 mux_c1_U17 ( .A1(mux_c1_n263), .A2(final_y[13]), .ZN(c1[13]) );
  AND2_X1 mux_c1_U16 ( .A1(mux_c1_n264), .A2(final_y[12]), .ZN(c1[12]) );
  AND2_X1 mux_c1_U15 ( .A1(mux_c1_n263), .A2(final_y[11]), .ZN(c1[11]) );
  AND2_X1 mux_c1_U14 ( .A1(mux_c1_n263), .A2(final_y[10]), .ZN(c1[10]) );
  AND2_X1 mux_c1_U13 ( .A1(mux_c1_n264), .A2(final_y[9]), .ZN(c1[9]) );
  AND2_X1 mux_c1_U12 ( .A1(mux_c1_n263), .A2(final_y[8]), .ZN(c1[8]) );
  AND2_X1 mux_c1_U11 ( .A1(mux_c1_n264), .A2(final_y[7]), .ZN(c1[7]) );
  AND2_X1 mux_c1_U10 ( .A1(mux_c1_n264), .A2(final_y[6]), .ZN(c1[6]) );
  AND2_X1 mux_c1_U9 ( .A1(mux_c1_n263), .A2(final_y[5]), .ZN(c1[5]) );
  AND2_X1 mux_c1_U8 ( .A1(mux_c1_n263), .A2(final_y[4]), .ZN(c1[4]) );
  AND2_X1 mux_c1_U7 ( .A1(mux_c1_n264), .A2(final_y[3]), .ZN(c1[3]) );
  AND2_X1 mux_c1_U6 ( .A1(mux_c1_n263), .A2(final_y[2]), .ZN(c1[2]) );
  AND2_X1 mux_c1_U5 ( .A1(mux_c1_n264), .A2(final_y[1]), .ZN(c1[1]) );
  AND2_X1 mux_c1_U4 ( .A1(mux_c1_n264), .A2(final_y[0]), .ZN(c1[0]) );
  INV_X1 mux_c1_U3 ( .A(mux_c1_n262), .ZN(mux_c1_n264) );
  INV_X1 mux_c1_U2 ( .A(mux_c1_n262), .ZN(mux_c1_n263) );
  INV_X1 mux_c1_U1 ( .A(done), .ZN(mux_c1_n262) );
endmodule

