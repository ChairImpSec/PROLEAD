module circuit ( clk, reset, data_in1, data_in2, data_in3, key, 
        data_out1, data_out2, data_out3, done );
  input [63:0] data_in1;
  input [63:0] data_in2;
  input [63:0] data_in3;
  input [79:0] key;
  output [63:0] data_out1;
  output [63:0] data_out2;
  output [63:0] data_out3;
  input clk, reset;
  output done;
  wire   enSboxReg, intDone, final, fsm_n35, fsm_n34, fsm_n33, fsm_n32,
         fsm_n31, fsm_n30, fsm_n29, fsm_n28, fsm_n27, fsm_n26, fsm_n25,
         fsm_n24, fsm_n23, fsm_n22, fsm_n21, fsm_n20, fsm_n19, fsm_n18,
         fsm_n17, fsm_n16, fsm_n15, fsm_n14, fsm_n13, fsm_n12, fsm_n11,
         fsm_n10, fsm_n43, fsm_n42, fsm_n41, fsm_n8, fsm_n7, fsm_ps_state_2_,
         fsm_en_countSerial, fsm_rst_countSerial, fsm_en_countRound,
         fsm_rst_countRound, fsm_cnt_rnd_n35, fsm_cnt_rnd_n34, fsm_cnt_rnd_n33,
         fsm_cnt_rnd_n32, fsm_cnt_rnd_n31, fsm_cnt_rnd_n30, fsm_cnt_rnd_n29,
         fsm_cnt_rnd_n28, fsm_cnt_rnd_n27, fsm_cnt_rnd_n26, fsm_cnt_rnd_n25,
         fsm_cnt_rnd_n1, fsm_cnt_rnd_n18, fsm_cnt_rnd_n17, fsm_cnt_rnd_n16,
         fsm_cnt_rnd_n15, fsm_cnt_rnd_n14, fsm_cnt_ser_n30, fsm_cnt_ser_n25,
         fsm_cnt_ser_n24, fsm_cnt_ser_n23, fsm_cnt_ser_n22, fsm_cnt_ser_n21,
         fsm_cnt_ser_n20, fsm_cnt_ser_n19, fsm_cnt_ser_n29, fsm_cnt_ser_n28,
         fsm_cnt_ser_n27, fsm_cnt_ser_n26, fsm_cnt_ser_n3, fsm_cnt_ser_n1,
         stateFF_n139, stateFF_n138, stateFF_n137, stateFF_n136, stateFF_n135,
         stateFF_state_n11, stateFF_state_n10, stateFF_state_n9,
         stateFF_state_n8, stateFF_state_n7, stateFF_state_gff_1_n41,
         stateFF_state_gff_1_n40, stateFF_state_gff_1_n39,
         stateFF_state_gff_1_n38, stateFF_state_gff_1_n37,
         stateFF_state_gff_1_n36, stateFF_state_gff_1_n35,
         stateFF_state_gff_1_n34, stateFF_state_gff_1_n33,
         stateFF_state_gff_1_n32, stateFF_state_gff_1_n31,
         stateFF_state_gff_1_n30, stateFF_state_gff_1_n29,
         stateFF_state_gff_1_n28, stateFF_state_gff_1_n27,
         stateFF_state_gff_1_n26, stateFF_state_gff_1_n25,
         stateFF_state_gff_1_n24, stateFF_state_gff_1_n23,
         stateFF_state_gff_1_n22, stateFF_state_gff_1_n21,
         stateFF_state_gff_1_n20, stateFF_state_gff_2_n67,
         stateFF_state_gff_2_n66, stateFF_state_gff_2_n65,
         stateFF_state_gff_2_n64, stateFF_state_gff_2_n63,
         stateFF_state_gff_2_n62, stateFF_state_gff_2_n61,
         stateFF_state_gff_2_n60, stateFF_state_gff_2_n59,
         stateFF_state_gff_2_n58, stateFF_state_gff_2_n57,
         stateFF_state_gff_2_n56, stateFF_state_gff_2_n55,
         stateFF_state_gff_2_n54, stateFF_state_gff_2_n35,
         stateFF_state_gff_2_n34, stateFF_state_gff_2_n33,
         stateFF_state_gff_2_n32, stateFF_state_gff_2_n31,
         stateFF_state_gff_2_n30, stateFF_state_gff_2_n29,
         stateFF_state_gff_2_n28, stateFF_state_gff_3_n68,
         stateFF_state_gff_3_n67, stateFF_state_gff_3_n66,
         stateFF_state_gff_3_n65, stateFF_state_gff_3_n64,
         stateFF_state_gff_3_n63, stateFF_state_gff_3_n62,
         stateFF_state_gff_3_n61, stateFF_state_gff_3_n60,
         stateFF_state_gff_3_n59, stateFF_state_gff_3_n58,
         stateFF_state_gff_3_n57, stateFF_state_gff_3_n56,
         stateFF_state_gff_3_n55, stateFF_state_gff_3_n54,
         stateFF_state_gff_3_n35, stateFF_state_gff_3_n34,
         stateFF_state_gff_3_n33, stateFF_state_gff_3_n32,
         stateFF_state_gff_3_n31, stateFF_state_gff_3_n30,
         stateFF_state_gff_3_n29, stateFF_state_gff_3_n28,
         stateFF_state_gff_4_n68, stateFF_state_gff_4_n67,
         stateFF_state_gff_4_n66, stateFF_state_gff_4_n65,
         stateFF_state_gff_4_n64, stateFF_state_gff_4_n63,
         stateFF_state_gff_4_n62, stateFF_state_gff_4_n61,
         stateFF_state_gff_4_n60, stateFF_state_gff_4_n59,
         stateFF_state_gff_4_n58, stateFF_state_gff_4_n57,
         stateFF_state_gff_4_n56, stateFF_state_gff_4_n55,
         stateFF_state_gff_4_n54, stateFF_state_gff_4_n35,
         stateFF_state_gff_4_n34, stateFF_state_gff_4_n33,
         stateFF_state_gff_4_n32, stateFF_state_gff_4_n31,
         stateFF_state_gff_4_n30, stateFF_state_gff_4_n29,
         stateFF_state_gff_4_n28, stateFF_state_gff_5_n68,
         stateFF_state_gff_5_n67, stateFF_state_gff_5_n66,
         stateFF_state_gff_5_n65, stateFF_state_gff_5_n64,
         stateFF_state_gff_5_n63, stateFF_state_gff_5_n62,
         stateFF_state_gff_5_n61, stateFF_state_gff_5_n60,
         stateFF_state_gff_5_n59, stateFF_state_gff_5_n58,
         stateFF_state_gff_5_n57, stateFF_state_gff_5_n56,
         stateFF_state_gff_5_n55, stateFF_state_gff_5_n54,
         stateFF_state_gff_5_n35, stateFF_state_gff_5_n34,
         stateFF_state_gff_5_n33, stateFF_state_gff_5_n32,
         stateFF_state_gff_5_n31, stateFF_state_gff_5_n30,
         stateFF_state_gff_5_n29, stateFF_state_gff_5_n28,
         stateFF_state_gff_6_n69, stateFF_state_gff_6_n68,
         stateFF_state_gff_6_n67, stateFF_state_gff_6_n66,
         stateFF_state_gff_6_n65, stateFF_state_gff_6_n64,
         stateFF_state_gff_6_n63, stateFF_state_gff_6_n62,
         stateFF_state_gff_6_n61, stateFF_state_gff_6_n60,
         stateFF_state_gff_6_n59, stateFF_state_gff_6_n58,
         stateFF_state_gff_6_n57, stateFF_state_gff_6_n56,
         stateFF_state_gff_6_n55, stateFF_state_gff_6_n36,
         stateFF_state_gff_6_n35, stateFF_state_gff_6_n34,
         stateFF_state_gff_6_n33, stateFF_state_gff_6_n32,
         stateFF_state_gff_6_n31, stateFF_state_gff_6_n30,
         stateFF_state_gff_6_n29, stateFF_state_gff_7_n69,
         stateFF_state_gff_7_n68, stateFF_state_gff_7_n67,
         stateFF_state_gff_7_n66, stateFF_state_gff_7_n65,
         stateFF_state_gff_7_n64, stateFF_state_gff_7_n63,
         stateFF_state_gff_7_n62, stateFF_state_gff_7_n61,
         stateFF_state_gff_7_n60, stateFF_state_gff_7_n59,
         stateFF_state_gff_7_n58, stateFF_state_gff_7_n57,
         stateFF_state_gff_7_n56, stateFF_state_gff_7_n55,
         stateFF_state_gff_7_n36, stateFF_state_gff_7_n35,
         stateFF_state_gff_7_n34, stateFF_state_gff_7_n33,
         stateFF_state_gff_7_n32, stateFF_state_gff_7_n31,
         stateFF_state_gff_7_n30, stateFF_state_gff_7_n29,
         stateFF_state_gff_8_n69, stateFF_state_gff_8_n68,
         stateFF_state_gff_8_n67, stateFF_state_gff_8_n66,
         stateFF_state_gff_8_n65, stateFF_state_gff_8_n64,
         stateFF_state_gff_8_n63, stateFF_state_gff_8_n62,
         stateFF_state_gff_8_n61, stateFF_state_gff_8_n60,
         stateFF_state_gff_8_n59, stateFF_state_gff_8_n58,
         stateFF_state_gff_8_n57, stateFF_state_gff_8_n56,
         stateFF_state_gff_8_n55, stateFF_state_gff_8_n36,
         stateFF_state_gff_8_n35, stateFF_state_gff_8_n34,
         stateFF_state_gff_8_n33, stateFF_state_gff_8_n32,
         stateFF_state_gff_8_n31, stateFF_state_gff_8_n30,
         stateFF_state_gff_8_n29, stateFF_state_gff_9_n69,
         stateFF_state_gff_9_n68, stateFF_state_gff_9_n67,
         stateFF_state_gff_9_n66, stateFF_state_gff_9_n65,
         stateFF_state_gff_9_n64, stateFF_state_gff_9_n63,
         stateFF_state_gff_9_n62, stateFF_state_gff_9_n61,
         stateFF_state_gff_9_n60, stateFF_state_gff_9_n59,
         stateFF_state_gff_9_n58, stateFF_state_gff_9_n57,
         stateFF_state_gff_9_n56, stateFF_state_gff_9_n55,
         stateFF_state_gff_9_n36, stateFF_state_gff_9_n35,
         stateFF_state_gff_9_n34, stateFF_state_gff_9_n33,
         stateFF_state_gff_9_n32, stateFF_state_gff_9_n31,
         stateFF_state_gff_9_n30, stateFF_state_gff_9_n29,
         stateFF_state_gff_10_n69, stateFF_state_gff_10_n68,
         stateFF_state_gff_10_n67, stateFF_state_gff_10_n66,
         stateFF_state_gff_10_n65, stateFF_state_gff_10_n64,
         stateFF_state_gff_10_n63, stateFF_state_gff_10_n62,
         stateFF_state_gff_10_n61, stateFF_state_gff_10_n60,
         stateFF_state_gff_10_n59, stateFF_state_gff_10_n58,
         stateFF_state_gff_10_n57, stateFF_state_gff_10_n56,
         stateFF_state_gff_10_n55, stateFF_state_gff_10_n36,
         stateFF_state_gff_10_n35, stateFF_state_gff_10_n34,
         stateFF_state_gff_10_n33, stateFF_state_gff_10_n32,
         stateFF_state_gff_10_n31, stateFF_state_gff_10_n30,
         stateFF_state_gff_10_n29, stateFF_state_gff_11_n69,
         stateFF_state_gff_11_n68, stateFF_state_gff_11_n67,
         stateFF_state_gff_11_n66, stateFF_state_gff_11_n65,
         stateFF_state_gff_11_n64, stateFF_state_gff_11_n63,
         stateFF_state_gff_11_n62, stateFF_state_gff_11_n61,
         stateFF_state_gff_11_n60, stateFF_state_gff_11_n59,
         stateFF_state_gff_11_n58, stateFF_state_gff_11_n57,
         stateFF_state_gff_11_n56, stateFF_state_gff_11_n55,
         stateFF_state_gff_11_n36, stateFF_state_gff_11_n35,
         stateFF_state_gff_11_n34, stateFF_state_gff_11_n33,
         stateFF_state_gff_11_n32, stateFF_state_gff_11_n31,
         stateFF_state_gff_11_n30, stateFF_state_gff_11_n29,
         stateFF_state_gff_12_n69, stateFF_state_gff_12_n68,
         stateFF_state_gff_12_n67, stateFF_state_gff_12_n66,
         stateFF_state_gff_12_n65, stateFF_state_gff_12_n64,
         stateFF_state_gff_12_n63, stateFF_state_gff_12_n62,
         stateFF_state_gff_12_n61, stateFF_state_gff_12_n60,
         stateFF_state_gff_12_n59, stateFF_state_gff_12_n58,
         stateFF_state_gff_12_n57, stateFF_state_gff_12_n56,
         stateFF_state_gff_12_n55, stateFF_state_gff_12_n36,
         stateFF_state_gff_12_n35, stateFF_state_gff_12_n34,
         stateFF_state_gff_12_n33, stateFF_state_gff_12_n32,
         stateFF_state_gff_12_n31, stateFF_state_gff_12_n30,
         stateFF_state_gff_12_n29, stateFF_state_gff_13_n69,
         stateFF_state_gff_13_n68, stateFF_state_gff_13_n67,
         stateFF_state_gff_13_n66, stateFF_state_gff_13_n65,
         stateFF_state_gff_13_n64, stateFF_state_gff_13_n63,
         stateFF_state_gff_13_n62, stateFF_state_gff_13_n61,
         stateFF_state_gff_13_n60, stateFF_state_gff_13_n59,
         stateFF_state_gff_13_n58, stateFF_state_gff_13_n57,
         stateFF_state_gff_13_n56, stateFF_state_gff_13_n55,
         stateFF_state_gff_13_n36, stateFF_state_gff_13_n35,
         stateFF_state_gff_13_n34, stateFF_state_gff_13_n33,
         stateFF_state_gff_13_n32, stateFF_state_gff_13_n31,
         stateFF_state_gff_13_n30, stateFF_state_gff_13_n29,
         stateFF_state_gff_14_n69, stateFF_state_gff_14_n68,
         stateFF_state_gff_14_n67, stateFF_state_gff_14_n66,
         stateFF_state_gff_14_n65, stateFF_state_gff_14_n64,
         stateFF_state_gff_14_n63, stateFF_state_gff_14_n62,
         stateFF_state_gff_14_n61, stateFF_state_gff_14_n60,
         stateFF_state_gff_14_n59, stateFF_state_gff_14_n58,
         stateFF_state_gff_14_n57, stateFF_state_gff_14_n56,
         stateFF_state_gff_14_n55, stateFF_state_gff_14_n36,
         stateFF_state_gff_14_n35, stateFF_state_gff_14_n34,
         stateFF_state_gff_14_n33, stateFF_state_gff_14_n32,
         stateFF_state_gff_14_n31, stateFF_state_gff_14_n30,
         stateFF_state_gff_14_n29, stateFF_state_gff_15_n69,
         stateFF_state_gff_15_n68, stateFF_state_gff_15_n67,
         stateFF_state_gff_15_n66, stateFF_state_gff_15_n65,
         stateFF_state_gff_15_n64, stateFF_state_gff_15_n63,
         stateFF_state_gff_15_n62, stateFF_state_gff_15_n61,
         stateFF_state_gff_15_n60, stateFF_state_gff_15_n59,
         stateFF_state_gff_15_n58, stateFF_state_gff_15_n57,
         stateFF_state_gff_15_n56, stateFF_state_gff_15_n55,
         stateFF_state_gff_15_n36, stateFF_state_gff_15_n35,
         stateFF_state_gff_15_n34, stateFF_state_gff_15_n33,
         stateFF_state_gff_15_n32, stateFF_state_gff_15_n31,
         stateFF_state_gff_15_n30, stateFF_state_gff_15_n29,
         stateFF_state_gff_16_n68, stateFF_state_gff_16_n67,
         stateFF_state_gff_16_n66, stateFF_state_gff_16_n65,
         stateFF_state_gff_16_n64, stateFF_state_gff_16_n63,
         stateFF_state_gff_16_n62, stateFF_state_gff_16_n61,
         stateFF_state_gff_16_n60, stateFF_state_gff_16_n59,
         stateFF_state_gff_16_n58, stateFF_state_gff_16_n57,
         stateFF_state_gff_16_n56, stateFF_state_gff_16_n55,
         stateFF_state_gff_16_n54, stateFF_state_gff_16_n35,
         stateFF_state_gff_16_n34, stateFF_state_gff_16_n33,
         stateFF_state_gff_16_n32, stateFF_state_gff_16_n31,
         stateFF_state_gff_16_n30, stateFF_state_gff_16_n29,
         stateFF_state_gff_16_n28, md1FF_n267, md1FF_n266, md1FF_n265,
         md1FF_n264, md1FF_n263, md1FF_state_n11, md1FF_state_n10,
         md1FF_state_n9, md1FF_state_n8, md1FF_state_n7, md1FF_state_gff_1_n67,
         md1FF_state_gff_1_n66, md1FF_state_gff_1_n65, md1FF_state_gff_1_n64,
         md1FF_state_gff_1_n63, md1FF_state_gff_1_n62, md1FF_state_gff_1_n61,
         md1FF_state_gff_1_n60, md1FF_state_gff_1_n59, md1FF_state_gff_1_n58,
         md1FF_state_gff_1_n57, md1FF_state_gff_1_n56, md1FF_state_gff_1_n55,
         md1FF_state_gff_1_n54, md1FF_state_gff_1_n35, md1FF_state_gff_1_n34,
         md1FF_state_gff_1_n33, md1FF_state_gff_1_n32, md1FF_state_gff_1_n31,
         md1FF_state_gff_1_n30, md1FF_state_gff_1_n29, md1FF_state_gff_1_n28,
         md1FF_state_gff_2_n68, md1FF_state_gff_2_n67, md1FF_state_gff_2_n66,
         md1FF_state_gff_2_n65, md1FF_state_gff_2_n64, md1FF_state_gff_2_n63,
         md1FF_state_gff_2_n62, md1FF_state_gff_2_n61, md1FF_state_gff_2_n60,
         md1FF_state_gff_2_n59, md1FF_state_gff_2_n58, md1FF_state_gff_2_n57,
         md1FF_state_gff_2_n56, md1FF_state_gff_2_n55, md1FF_state_gff_2_n54,
         md1FF_state_gff_2_n35, md1FF_state_gff_2_n34, md1FF_state_gff_2_n33,
         md1FF_state_gff_2_n32, md1FF_state_gff_2_n31, md1FF_state_gff_2_n30,
         md1FF_state_gff_2_n29, md1FF_state_gff_2_n28, md1FF_state_gff_3_n68,
         md1FF_state_gff_3_n67, md1FF_state_gff_3_n66, md1FF_state_gff_3_n65,
         md1FF_state_gff_3_n64, md1FF_state_gff_3_n63, md1FF_state_gff_3_n62,
         md1FF_state_gff_3_n61, md1FF_state_gff_3_n60, md1FF_state_gff_3_n59,
         md1FF_state_gff_3_n58, md1FF_state_gff_3_n57, md1FF_state_gff_3_n56,
         md1FF_state_gff_3_n55, md1FF_state_gff_3_n54, md1FF_state_gff_3_n35,
         md1FF_state_gff_3_n34, md1FF_state_gff_3_n33, md1FF_state_gff_3_n32,
         md1FF_state_gff_3_n31, md1FF_state_gff_3_n30, md1FF_state_gff_3_n29,
         md1FF_state_gff_3_n28, md1FF_state_gff_4_n68, md1FF_state_gff_4_n67,
         md1FF_state_gff_4_n66, md1FF_state_gff_4_n65, md1FF_state_gff_4_n64,
         md1FF_state_gff_4_n63, md1FF_state_gff_4_n62, md1FF_state_gff_4_n61,
         md1FF_state_gff_4_n60, md1FF_state_gff_4_n59, md1FF_state_gff_4_n58,
         md1FF_state_gff_4_n57, md1FF_state_gff_4_n56, md1FF_state_gff_4_n55,
         md1FF_state_gff_4_n54, md1FF_state_gff_4_n35, md1FF_state_gff_4_n34,
         md1FF_state_gff_4_n33, md1FF_state_gff_4_n32, md1FF_state_gff_4_n31,
         md1FF_state_gff_4_n30, md1FF_state_gff_4_n29, md1FF_state_gff_4_n28,
         md1FF_state_gff_5_n69, md1FF_state_gff_5_n68, md1FF_state_gff_5_n67,
         md1FF_state_gff_5_n66, md1FF_state_gff_5_n65, md1FF_state_gff_5_n64,
         md1FF_state_gff_5_n63, md1FF_state_gff_5_n62, md1FF_state_gff_5_n61,
         md1FF_state_gff_5_n60, md1FF_state_gff_5_n59, md1FF_state_gff_5_n58,
         md1FF_state_gff_5_n57, md1FF_state_gff_5_n56, md1FF_state_gff_5_n55,
         md1FF_state_gff_5_n36, md1FF_state_gff_5_n35, md1FF_state_gff_5_n34,
         md1FF_state_gff_5_n33, md1FF_state_gff_5_n32, md1FF_state_gff_5_n31,
         md1FF_state_gff_5_n30, md1FF_state_gff_5_n29, md1FF_state_gff_6_n69,
         md1FF_state_gff_6_n68, md1FF_state_gff_6_n67, md1FF_state_gff_6_n66,
         md1FF_state_gff_6_n65, md1FF_state_gff_6_n64, md1FF_state_gff_6_n63,
         md1FF_state_gff_6_n62, md1FF_state_gff_6_n61, md1FF_state_gff_6_n60,
         md1FF_state_gff_6_n59, md1FF_state_gff_6_n58, md1FF_state_gff_6_n57,
         md1FF_state_gff_6_n56, md1FF_state_gff_6_n55, md1FF_state_gff_6_n36,
         md1FF_state_gff_6_n35, md1FF_state_gff_6_n34, md1FF_state_gff_6_n33,
         md1FF_state_gff_6_n32, md1FF_state_gff_6_n31, md1FF_state_gff_6_n30,
         md1FF_state_gff_6_n29, md1FF_state_gff_7_n69, md1FF_state_gff_7_n68,
         md1FF_state_gff_7_n67, md1FF_state_gff_7_n66, md1FF_state_gff_7_n65,
         md1FF_state_gff_7_n64, md1FF_state_gff_7_n63, md1FF_state_gff_7_n62,
         md1FF_state_gff_7_n61, md1FF_state_gff_7_n60, md1FF_state_gff_7_n59,
         md1FF_state_gff_7_n58, md1FF_state_gff_7_n57, md1FF_state_gff_7_n56,
         md1FF_state_gff_7_n55, md1FF_state_gff_7_n36, md1FF_state_gff_7_n35,
         md1FF_state_gff_7_n34, md1FF_state_gff_7_n33, md1FF_state_gff_7_n32,
         md1FF_state_gff_7_n31, md1FF_state_gff_7_n30, md1FF_state_gff_7_n29,
         md1FF_state_gff_8_n69, md1FF_state_gff_8_n68, md1FF_state_gff_8_n67,
         md1FF_state_gff_8_n66, md1FF_state_gff_8_n65, md1FF_state_gff_8_n64,
         md1FF_state_gff_8_n63, md1FF_state_gff_8_n62, md1FF_state_gff_8_n61,
         md1FF_state_gff_8_n60, md1FF_state_gff_8_n59, md1FF_state_gff_8_n58,
         md1FF_state_gff_8_n57, md1FF_state_gff_8_n56, md1FF_state_gff_8_n55,
         md1FF_state_gff_8_n36, md1FF_state_gff_8_n35, md1FF_state_gff_8_n34,
         md1FF_state_gff_8_n33, md1FF_state_gff_8_n32, md1FF_state_gff_8_n31,
         md1FF_state_gff_8_n30, md1FF_state_gff_8_n29, md1FF_state_gff_9_n69,
         md1FF_state_gff_9_n68, md1FF_state_gff_9_n67, md1FF_state_gff_9_n66,
         md1FF_state_gff_9_n65, md1FF_state_gff_9_n64, md1FF_state_gff_9_n63,
         md1FF_state_gff_9_n62, md1FF_state_gff_9_n61, md1FF_state_gff_9_n60,
         md1FF_state_gff_9_n59, md1FF_state_gff_9_n58, md1FF_state_gff_9_n57,
         md1FF_state_gff_9_n56, md1FF_state_gff_9_n55, md1FF_state_gff_9_n36,
         md1FF_state_gff_9_n35, md1FF_state_gff_9_n34, md1FF_state_gff_9_n33,
         md1FF_state_gff_9_n32, md1FF_state_gff_9_n31, md1FF_state_gff_9_n30,
         md1FF_state_gff_9_n29, md1FF_state_gff_10_n69, md1FF_state_gff_10_n68,
         md1FF_state_gff_10_n67, md1FF_state_gff_10_n66,
         md1FF_state_gff_10_n65, md1FF_state_gff_10_n64,
         md1FF_state_gff_10_n63, md1FF_state_gff_10_n62,
         md1FF_state_gff_10_n61, md1FF_state_gff_10_n60,
         md1FF_state_gff_10_n59, md1FF_state_gff_10_n58,
         md1FF_state_gff_10_n57, md1FF_state_gff_10_n56,
         md1FF_state_gff_10_n55, md1FF_state_gff_10_n36,
         md1FF_state_gff_10_n35, md1FF_state_gff_10_n34,
         md1FF_state_gff_10_n33, md1FF_state_gff_10_n32,
         md1FF_state_gff_10_n31, md1FF_state_gff_10_n30,
         md1FF_state_gff_10_n29, md1FF_state_gff_11_n69,
         md1FF_state_gff_11_n68, md1FF_state_gff_11_n67,
         md1FF_state_gff_11_n66, md1FF_state_gff_11_n65,
         md1FF_state_gff_11_n64, md1FF_state_gff_11_n63,
         md1FF_state_gff_11_n62, md1FF_state_gff_11_n61,
         md1FF_state_gff_11_n60, md1FF_state_gff_11_n59,
         md1FF_state_gff_11_n58, md1FF_state_gff_11_n57,
         md1FF_state_gff_11_n56, md1FF_state_gff_11_n55,
         md1FF_state_gff_11_n36, md1FF_state_gff_11_n35,
         md1FF_state_gff_11_n34, md1FF_state_gff_11_n33,
         md1FF_state_gff_11_n32, md1FF_state_gff_11_n31,
         md1FF_state_gff_11_n30, md1FF_state_gff_11_n29,
         md1FF_state_gff_12_n69, md1FF_state_gff_12_n68,
         md1FF_state_gff_12_n67, md1FF_state_gff_12_n66,
         md1FF_state_gff_12_n65, md1FF_state_gff_12_n64,
         md1FF_state_gff_12_n63, md1FF_state_gff_12_n62,
         md1FF_state_gff_12_n61, md1FF_state_gff_12_n60,
         md1FF_state_gff_12_n59, md1FF_state_gff_12_n58,
         md1FF_state_gff_12_n57, md1FF_state_gff_12_n56,
         md1FF_state_gff_12_n55, md1FF_state_gff_12_n36,
         md1FF_state_gff_12_n35, md1FF_state_gff_12_n34,
         md1FF_state_gff_12_n33, md1FF_state_gff_12_n32,
         md1FF_state_gff_12_n31, md1FF_state_gff_12_n30,
         md1FF_state_gff_12_n29, md1FF_state_gff_13_n69,
         md1FF_state_gff_13_n68, md1FF_state_gff_13_n67,
         md1FF_state_gff_13_n66, md1FF_state_gff_13_n65,
         md1FF_state_gff_13_n64, md1FF_state_gff_13_n63,
         md1FF_state_gff_13_n62, md1FF_state_gff_13_n61,
         md1FF_state_gff_13_n60, md1FF_state_gff_13_n59,
         md1FF_state_gff_13_n58, md1FF_state_gff_13_n57,
         md1FF_state_gff_13_n56, md1FF_state_gff_13_n55,
         md1FF_state_gff_13_n36, md1FF_state_gff_13_n35,
         md1FF_state_gff_13_n34, md1FF_state_gff_13_n33,
         md1FF_state_gff_13_n32, md1FF_state_gff_13_n31,
         md1FF_state_gff_13_n30, md1FF_state_gff_13_n29,
         md1FF_state_gff_14_n69, md1FF_state_gff_14_n68,
         md1FF_state_gff_14_n67, md1FF_state_gff_14_n66,
         md1FF_state_gff_14_n65, md1FF_state_gff_14_n64,
         md1FF_state_gff_14_n63, md1FF_state_gff_14_n62,
         md1FF_state_gff_14_n61, md1FF_state_gff_14_n60,
         md1FF_state_gff_14_n59, md1FF_state_gff_14_n58,
         md1FF_state_gff_14_n57, md1FF_state_gff_14_n56,
         md1FF_state_gff_14_n55, md1FF_state_gff_14_n36,
         md1FF_state_gff_14_n35, md1FF_state_gff_14_n34,
         md1FF_state_gff_14_n33, md1FF_state_gff_14_n32,
         md1FF_state_gff_14_n31, md1FF_state_gff_14_n30,
         md1FF_state_gff_14_n29, md1FF_state_gff_15_n68,
         md1FF_state_gff_15_n67, md1FF_state_gff_15_n66,
         md1FF_state_gff_15_n65, md1FF_state_gff_15_n64,
         md1FF_state_gff_15_n63, md1FF_state_gff_15_n62,
         md1FF_state_gff_15_n61, md1FF_state_gff_15_n60,
         md1FF_state_gff_15_n59, md1FF_state_gff_15_n58,
         md1FF_state_gff_15_n57, md1FF_state_gff_15_n56,
         md1FF_state_gff_15_n55, md1FF_state_gff_15_n54,
         md1FF_state_gff_15_n35, md1FF_state_gff_15_n34,
         md1FF_state_gff_15_n33, md1FF_state_gff_15_n32,
         md1FF_state_gff_15_n31, md1FF_state_gff_15_n30,
         md1FF_state_gff_15_n29, md1FF_state_gff_15_n28,
         md1FF_state_gff_16_n68, md1FF_state_gff_16_n67,
         md1FF_state_gff_16_n66, md1FF_state_gff_16_n65,
         md1FF_state_gff_16_n64, md1FF_state_gff_16_n63,
         md1FF_state_gff_16_n62, md1FF_state_gff_16_n61,
         md1FF_state_gff_16_n60, md1FF_state_gff_16_n59,
         md1FF_state_gff_16_n58, md1FF_state_gff_16_n57,
         md1FF_state_gff_16_n56, md1FF_state_gff_16_n55,
         md1FF_state_gff_16_n54, md1FF_state_gff_16_n35,
         md1FF_state_gff_16_n34, md1FF_state_gff_16_n33,
         md1FF_state_gff_16_n32, md1FF_state_gff_16_n31,
         md1FF_state_gff_16_n30, md1FF_state_gff_16_n29,
         md1FF_state_gff_16_n28, md2FF_n267, md2FF_n266, md2FF_n265,
         md2FF_n264, md2FF_n263, md2FF_state_n11, md2FF_state_n10,
         md2FF_state_n9, md2FF_state_n8, md2FF_state_n7, md2FF_state_gff_1_n67,
         md2FF_state_gff_1_n66, md2FF_state_gff_1_n65, md2FF_state_gff_1_n64,
         md2FF_state_gff_1_n63, md2FF_state_gff_1_n62, md2FF_state_gff_1_n61,
         md2FF_state_gff_1_n60, md2FF_state_gff_1_n59, md2FF_state_gff_1_n58,
         md2FF_state_gff_1_n57, md2FF_state_gff_1_n56, md2FF_state_gff_1_n55,
         md2FF_state_gff_1_n54, md2FF_state_gff_1_n35, md2FF_state_gff_1_n34,
         md2FF_state_gff_1_n33, md2FF_state_gff_1_n32, md2FF_state_gff_1_n31,
         md2FF_state_gff_1_n30, md2FF_state_gff_1_n29, md2FF_state_gff_1_n28,
         md2FF_state_gff_2_n68, md2FF_state_gff_2_n67, md2FF_state_gff_2_n66,
         md2FF_state_gff_2_n65, md2FF_state_gff_2_n64, md2FF_state_gff_2_n63,
         md2FF_state_gff_2_n62, md2FF_state_gff_2_n61, md2FF_state_gff_2_n60,
         md2FF_state_gff_2_n59, md2FF_state_gff_2_n58, md2FF_state_gff_2_n57,
         md2FF_state_gff_2_n56, md2FF_state_gff_2_n55, md2FF_state_gff_2_n54,
         md2FF_state_gff_2_n35, md2FF_state_gff_2_n34, md2FF_state_gff_2_n33,
         md2FF_state_gff_2_n32, md2FF_state_gff_2_n31, md2FF_state_gff_2_n30,
         md2FF_state_gff_2_n29, md2FF_state_gff_2_n28, md2FF_state_gff_3_n68,
         md2FF_state_gff_3_n67, md2FF_state_gff_3_n66, md2FF_state_gff_3_n65,
         md2FF_state_gff_3_n64, md2FF_state_gff_3_n63, md2FF_state_gff_3_n62,
         md2FF_state_gff_3_n61, md2FF_state_gff_3_n60, md2FF_state_gff_3_n59,
         md2FF_state_gff_3_n58, md2FF_state_gff_3_n57, md2FF_state_gff_3_n56,
         md2FF_state_gff_3_n55, md2FF_state_gff_3_n54, md2FF_state_gff_3_n35,
         md2FF_state_gff_3_n34, md2FF_state_gff_3_n33, md2FF_state_gff_3_n32,
         md2FF_state_gff_3_n31, md2FF_state_gff_3_n30, md2FF_state_gff_3_n29,
         md2FF_state_gff_3_n28, md2FF_state_gff_4_n68, md2FF_state_gff_4_n67,
         md2FF_state_gff_4_n66, md2FF_state_gff_4_n65, md2FF_state_gff_4_n64,
         md2FF_state_gff_4_n63, md2FF_state_gff_4_n62, md2FF_state_gff_4_n61,
         md2FF_state_gff_4_n60, md2FF_state_gff_4_n59, md2FF_state_gff_4_n58,
         md2FF_state_gff_4_n57, md2FF_state_gff_4_n56, md2FF_state_gff_4_n55,
         md2FF_state_gff_4_n54, md2FF_state_gff_4_n35, md2FF_state_gff_4_n34,
         md2FF_state_gff_4_n33, md2FF_state_gff_4_n32, md2FF_state_gff_4_n31,
         md2FF_state_gff_4_n30, md2FF_state_gff_4_n29, md2FF_state_gff_4_n28,
         md2FF_state_gff_5_n69, md2FF_state_gff_5_n68, md2FF_state_gff_5_n67,
         md2FF_state_gff_5_n66, md2FF_state_gff_5_n65, md2FF_state_gff_5_n64,
         md2FF_state_gff_5_n63, md2FF_state_gff_5_n62, md2FF_state_gff_5_n61,
         md2FF_state_gff_5_n60, md2FF_state_gff_5_n59, md2FF_state_gff_5_n58,
         md2FF_state_gff_5_n57, md2FF_state_gff_5_n56, md2FF_state_gff_5_n55,
         md2FF_state_gff_5_n36, md2FF_state_gff_5_n35, md2FF_state_gff_5_n34,
         md2FF_state_gff_5_n33, md2FF_state_gff_5_n32, md2FF_state_gff_5_n31,
         md2FF_state_gff_5_n30, md2FF_state_gff_5_n29, md2FF_state_gff_6_n69,
         md2FF_state_gff_6_n68, md2FF_state_gff_6_n67, md2FF_state_gff_6_n66,
         md2FF_state_gff_6_n65, md2FF_state_gff_6_n64, md2FF_state_gff_6_n63,
         md2FF_state_gff_6_n62, md2FF_state_gff_6_n61, md2FF_state_gff_6_n60,
         md2FF_state_gff_6_n59, md2FF_state_gff_6_n58, md2FF_state_gff_6_n57,
         md2FF_state_gff_6_n56, md2FF_state_gff_6_n55, md2FF_state_gff_6_n36,
         md2FF_state_gff_6_n35, md2FF_state_gff_6_n34, md2FF_state_gff_6_n33,
         md2FF_state_gff_6_n32, md2FF_state_gff_6_n31, md2FF_state_gff_6_n30,
         md2FF_state_gff_6_n29, md2FF_state_gff_7_n69, md2FF_state_gff_7_n68,
         md2FF_state_gff_7_n67, md2FF_state_gff_7_n66, md2FF_state_gff_7_n65,
         md2FF_state_gff_7_n64, md2FF_state_gff_7_n63, md2FF_state_gff_7_n62,
         md2FF_state_gff_7_n61, md2FF_state_gff_7_n60, md2FF_state_gff_7_n59,
         md2FF_state_gff_7_n58, md2FF_state_gff_7_n57, md2FF_state_gff_7_n56,
         md2FF_state_gff_7_n55, md2FF_state_gff_7_n36, md2FF_state_gff_7_n35,
         md2FF_state_gff_7_n34, md2FF_state_gff_7_n33, md2FF_state_gff_7_n32,
         md2FF_state_gff_7_n31, md2FF_state_gff_7_n30, md2FF_state_gff_7_n29,
         md2FF_state_gff_8_n69, md2FF_state_gff_8_n68, md2FF_state_gff_8_n67,
         md2FF_state_gff_8_n66, md2FF_state_gff_8_n65, md2FF_state_gff_8_n64,
         md2FF_state_gff_8_n63, md2FF_state_gff_8_n62, md2FF_state_gff_8_n61,
         md2FF_state_gff_8_n60, md2FF_state_gff_8_n59, md2FF_state_gff_8_n58,
         md2FF_state_gff_8_n57, md2FF_state_gff_8_n56, md2FF_state_gff_8_n55,
         md2FF_state_gff_8_n36, md2FF_state_gff_8_n35, md2FF_state_gff_8_n34,
         md2FF_state_gff_8_n33, md2FF_state_gff_8_n32, md2FF_state_gff_8_n31,
         md2FF_state_gff_8_n30, md2FF_state_gff_8_n29, md2FF_state_gff_9_n69,
         md2FF_state_gff_9_n68, md2FF_state_gff_9_n67, md2FF_state_gff_9_n66,
         md2FF_state_gff_9_n65, md2FF_state_gff_9_n64, md2FF_state_gff_9_n63,
         md2FF_state_gff_9_n62, md2FF_state_gff_9_n61, md2FF_state_gff_9_n60,
         md2FF_state_gff_9_n59, md2FF_state_gff_9_n58, md2FF_state_gff_9_n57,
         md2FF_state_gff_9_n56, md2FF_state_gff_9_n55, md2FF_state_gff_9_n36,
         md2FF_state_gff_9_n35, md2FF_state_gff_9_n34, md2FF_state_gff_9_n33,
         md2FF_state_gff_9_n32, md2FF_state_gff_9_n31, md2FF_state_gff_9_n30,
         md2FF_state_gff_9_n29, md2FF_state_gff_10_n69, md2FF_state_gff_10_n68,
         md2FF_state_gff_10_n67, md2FF_state_gff_10_n66,
         md2FF_state_gff_10_n65, md2FF_state_gff_10_n64,
         md2FF_state_gff_10_n63, md2FF_state_gff_10_n62,
         md2FF_state_gff_10_n61, md2FF_state_gff_10_n60,
         md2FF_state_gff_10_n59, md2FF_state_gff_10_n58,
         md2FF_state_gff_10_n57, md2FF_state_gff_10_n56,
         md2FF_state_gff_10_n55, md2FF_state_gff_10_n36,
         md2FF_state_gff_10_n35, md2FF_state_gff_10_n34,
         md2FF_state_gff_10_n33, md2FF_state_gff_10_n32,
         md2FF_state_gff_10_n31, md2FF_state_gff_10_n30,
         md2FF_state_gff_10_n29, md2FF_state_gff_11_n69,
         md2FF_state_gff_11_n68, md2FF_state_gff_11_n67,
         md2FF_state_gff_11_n66, md2FF_state_gff_11_n65,
         md2FF_state_gff_11_n64, md2FF_state_gff_11_n63,
         md2FF_state_gff_11_n62, md2FF_state_gff_11_n61,
         md2FF_state_gff_11_n60, md2FF_state_gff_11_n59,
         md2FF_state_gff_11_n58, md2FF_state_gff_11_n57,
         md2FF_state_gff_11_n56, md2FF_state_gff_11_n55,
         md2FF_state_gff_11_n36, md2FF_state_gff_11_n35,
         md2FF_state_gff_11_n34, md2FF_state_gff_11_n33,
         md2FF_state_gff_11_n32, md2FF_state_gff_11_n31,
         md2FF_state_gff_11_n30, md2FF_state_gff_11_n29,
         md2FF_state_gff_12_n69, md2FF_state_gff_12_n68,
         md2FF_state_gff_12_n67, md2FF_state_gff_12_n66,
         md2FF_state_gff_12_n65, md2FF_state_gff_12_n64,
         md2FF_state_gff_12_n63, md2FF_state_gff_12_n62,
         md2FF_state_gff_12_n61, md2FF_state_gff_12_n60,
         md2FF_state_gff_12_n59, md2FF_state_gff_12_n58,
         md2FF_state_gff_12_n57, md2FF_state_gff_12_n56,
         md2FF_state_gff_12_n55, md2FF_state_gff_12_n36,
         md2FF_state_gff_12_n35, md2FF_state_gff_12_n34,
         md2FF_state_gff_12_n33, md2FF_state_gff_12_n32,
         md2FF_state_gff_12_n31, md2FF_state_gff_12_n30,
         md2FF_state_gff_12_n29, md2FF_state_gff_13_n69,
         md2FF_state_gff_13_n68, md2FF_state_gff_13_n67,
         md2FF_state_gff_13_n66, md2FF_state_gff_13_n65,
         md2FF_state_gff_13_n64, md2FF_state_gff_13_n63,
         md2FF_state_gff_13_n62, md2FF_state_gff_13_n61,
         md2FF_state_gff_13_n60, md2FF_state_gff_13_n59,
         md2FF_state_gff_13_n58, md2FF_state_gff_13_n57,
         md2FF_state_gff_13_n56, md2FF_state_gff_13_n55,
         md2FF_state_gff_13_n36, md2FF_state_gff_13_n35,
         md2FF_state_gff_13_n34, md2FF_state_gff_13_n33,
         md2FF_state_gff_13_n32, md2FF_state_gff_13_n31,
         md2FF_state_gff_13_n30, md2FF_state_gff_13_n29,
         md2FF_state_gff_14_n69, md2FF_state_gff_14_n68,
         md2FF_state_gff_14_n67, md2FF_state_gff_14_n66,
         md2FF_state_gff_14_n65, md2FF_state_gff_14_n64,
         md2FF_state_gff_14_n63, md2FF_state_gff_14_n62,
         md2FF_state_gff_14_n61, md2FF_state_gff_14_n60,
         md2FF_state_gff_14_n59, md2FF_state_gff_14_n58,
         md2FF_state_gff_14_n57, md2FF_state_gff_14_n56,
         md2FF_state_gff_14_n55, md2FF_state_gff_14_n36,
         md2FF_state_gff_14_n35, md2FF_state_gff_14_n34,
         md2FF_state_gff_14_n33, md2FF_state_gff_14_n32,
         md2FF_state_gff_14_n31, md2FF_state_gff_14_n30,
         md2FF_state_gff_14_n29, md2FF_state_gff_15_n68,
         md2FF_state_gff_15_n67, md2FF_state_gff_15_n66,
         md2FF_state_gff_15_n65, md2FF_state_gff_15_n64,
         md2FF_state_gff_15_n63, md2FF_state_gff_15_n62,
         md2FF_state_gff_15_n61, md2FF_state_gff_15_n60,
         md2FF_state_gff_15_n59, md2FF_state_gff_15_n58,
         md2FF_state_gff_15_n57, md2FF_state_gff_15_n56,
         md2FF_state_gff_15_n55, md2FF_state_gff_15_n54,
         md2FF_state_gff_15_n35, md2FF_state_gff_15_n34,
         md2FF_state_gff_15_n33, md2FF_state_gff_15_n32,
         md2FF_state_gff_15_n31, md2FF_state_gff_15_n30,
         md2FF_state_gff_15_n29, md2FF_state_gff_15_n28,
         md2FF_state_gff_16_n68, md2FF_state_gff_16_n67,
         md2FF_state_gff_16_n66, md2FF_state_gff_16_n65,
         md2FF_state_gff_16_n64, md2FF_state_gff_16_n63,
         md2FF_state_gff_16_n62, md2FF_state_gff_16_n61,
         md2FF_state_gff_16_n60, md2FF_state_gff_16_n59,
         md2FF_state_gff_16_n58, md2FF_state_gff_16_n57,
         md2FF_state_gff_16_n56, md2FF_state_gff_16_n55,
         md2FF_state_gff_16_n54, md2FF_state_gff_16_n35,
         md2FF_state_gff_16_n34, md2FF_state_gff_16_n33,
         md2FF_state_gff_16_n32, md2FF_state_gff_16_n31,
         md2FF_state_gff_16_n30, md2FF_state_gff_16_n29,
         md2FF_state_gff_16_n28, keyFF_n183, keyFF_n182, keyFF_n181,
         keyFF_n180, keyFF_n179, keyFF_n178, keyFF_n177, keyFF_n176,
         keyFF_n175, keyFF_n174, keyFF_keystate_n8, keyFF_keystate_n7,
         keyFF_keystate_n6, keyFF_keystate_gff_1_n68, keyFF_keystate_gff_1_n67,
         keyFF_keystate_gff_1_n66, keyFF_keystate_gff_1_n65,
         keyFF_keystate_gff_1_n64, keyFF_keystate_gff_1_n63,
         keyFF_keystate_gff_1_n62, keyFF_keystate_gff_1_n61,
         keyFF_keystate_gff_1_n60, keyFF_keystate_gff_1_n59,
         keyFF_keystate_gff_1_n58, keyFF_keystate_gff_1_n57,
         keyFF_keystate_gff_1_n56, keyFF_keystate_gff_1_n55,
         keyFF_keystate_gff_1_n36, keyFF_keystate_gff_1_n35,
         keyFF_keystate_gff_1_n34, keyFF_keystate_gff_1_n33,
         keyFF_keystate_gff_1_n32, keyFF_keystate_gff_1_n31,
         keyFF_keystate_gff_1_n30, keyFF_keystate_gff_1_n29,
         keyFF_keystate_gff_2_n68, keyFF_keystate_gff_2_n67,
         keyFF_keystate_gff_2_n66, keyFF_keystate_gff_2_n65,
         keyFF_keystate_gff_2_n64, keyFF_keystate_gff_2_n63,
         keyFF_keystate_gff_2_n62, keyFF_keystate_gff_2_n61,
         keyFF_keystate_gff_2_n60, keyFF_keystate_gff_2_n59,
         keyFF_keystate_gff_2_n58, keyFF_keystate_gff_2_n57,
         keyFF_keystate_gff_2_n56, keyFF_keystate_gff_2_n55,
         keyFF_keystate_gff_2_n36, keyFF_keystate_gff_2_n35,
         keyFF_keystate_gff_2_n34, keyFF_keystate_gff_2_n33,
         keyFF_keystate_gff_2_n32, keyFF_keystate_gff_2_n31,
         keyFF_keystate_gff_2_n30, keyFF_keystate_gff_2_n29,
         keyFF_keystate_gff_3_n68, keyFF_keystate_gff_3_n67,
         keyFF_keystate_gff_3_n66, keyFF_keystate_gff_3_n65,
         keyFF_keystate_gff_3_n64, keyFF_keystate_gff_3_n63,
         keyFF_keystate_gff_3_n62, keyFF_keystate_gff_3_n61,
         keyFF_keystate_gff_3_n60, keyFF_keystate_gff_3_n59,
         keyFF_keystate_gff_3_n58, keyFF_keystate_gff_3_n57,
         keyFF_keystate_gff_3_n56, keyFF_keystate_gff_3_n55,
         keyFF_keystate_gff_3_n36, keyFF_keystate_gff_3_n35,
         keyFF_keystate_gff_3_n34, keyFF_keystate_gff_3_n33,
         keyFF_keystate_gff_3_n32, keyFF_keystate_gff_3_n31,
         keyFF_keystate_gff_3_n30, keyFF_keystate_gff_3_n29,
         keyFF_keystate_gff_4_n68, keyFF_keystate_gff_4_n67,
         keyFF_keystate_gff_4_n66, keyFF_keystate_gff_4_n65,
         keyFF_keystate_gff_4_n64, keyFF_keystate_gff_4_n63,
         keyFF_keystate_gff_4_n62, keyFF_keystate_gff_4_n61,
         keyFF_keystate_gff_4_n60, keyFF_keystate_gff_4_n59,
         keyFF_keystate_gff_4_n58, keyFF_keystate_gff_4_n57,
         keyFF_keystate_gff_4_n56, keyFF_keystate_gff_4_n55,
         keyFF_keystate_gff_4_n36, keyFF_keystate_gff_4_n35,
         keyFF_keystate_gff_4_n34, keyFF_keystate_gff_4_n33,
         keyFF_keystate_gff_4_n32, keyFF_keystate_gff_4_n31,
         keyFF_keystate_gff_4_n30, keyFF_keystate_gff_4_n29,
         keyFF_keystate_gff_5_n69, keyFF_keystate_gff_5_n68,
         keyFF_keystate_gff_5_n67, keyFF_keystate_gff_5_n66,
         keyFF_keystate_gff_5_n65, keyFF_keystate_gff_5_n64,
         keyFF_keystate_gff_5_n63, keyFF_keystate_gff_5_n62,
         keyFF_keystate_gff_5_n61, keyFF_keystate_gff_5_n60,
         keyFF_keystate_gff_5_n59, keyFF_keystate_gff_5_n58,
         keyFF_keystate_gff_5_n57, keyFF_keystate_gff_5_n56,
         keyFF_keystate_gff_5_n55, keyFF_keystate_gff_5_n36,
         keyFF_keystate_gff_5_n35, keyFF_keystate_gff_5_n34,
         keyFF_keystate_gff_5_n33, keyFF_keystate_gff_5_n32,
         keyFF_keystate_gff_5_n31, keyFF_keystate_gff_5_n30,
         keyFF_keystate_gff_5_n29, keyFF_keystate_gff_6_n68,
         keyFF_keystate_gff_6_n67, keyFF_keystate_gff_6_n66,
         keyFF_keystate_gff_6_n65, keyFF_keystate_gff_6_n64,
         keyFF_keystate_gff_6_n63, keyFF_keystate_gff_6_n62,
         keyFF_keystate_gff_6_n61, keyFF_keystate_gff_6_n60,
         keyFF_keystate_gff_6_n59, keyFF_keystate_gff_6_n58,
         keyFF_keystate_gff_6_n57, keyFF_keystate_gff_6_n56,
         keyFF_keystate_gff_6_n55, keyFF_keystate_gff_6_n54,
         keyFF_keystate_gff_6_n35, keyFF_keystate_gff_6_n34,
         keyFF_keystate_gff_6_n33, keyFF_keystate_gff_6_n32,
         keyFF_keystate_gff_6_n31, keyFF_keystate_gff_6_n30,
         keyFF_keystate_gff_6_n29, keyFF_keystate_gff_6_n28,
         keyFF_keystate_gff_7_n68, keyFF_keystate_gff_7_n67,
         keyFF_keystate_gff_7_n66, keyFF_keystate_gff_7_n65,
         keyFF_keystate_gff_7_n64, keyFF_keystate_gff_7_n63,
         keyFF_keystate_gff_7_n62, keyFF_keystate_gff_7_n61,
         keyFF_keystate_gff_7_n60, keyFF_keystate_gff_7_n59,
         keyFF_keystate_gff_7_n58, keyFF_keystate_gff_7_n57,
         keyFF_keystate_gff_7_n56, keyFF_keystate_gff_7_n55,
         keyFF_keystate_gff_7_n54, keyFF_keystate_gff_7_n35,
         keyFF_keystate_gff_7_n34, keyFF_keystate_gff_7_n33,
         keyFF_keystate_gff_7_n32, keyFF_keystate_gff_7_n31,
         keyFF_keystate_gff_7_n30, keyFF_keystate_gff_7_n29,
         keyFF_keystate_gff_7_n28, keyFF_keystate_gff_8_n68,
         keyFF_keystate_gff_8_n67, keyFF_keystate_gff_8_n66,
         keyFF_keystate_gff_8_n65, keyFF_keystate_gff_8_n64,
         keyFF_keystate_gff_8_n63, keyFF_keystate_gff_8_n62,
         keyFF_keystate_gff_8_n61, keyFF_keystate_gff_8_n60,
         keyFF_keystate_gff_8_n59, keyFF_keystate_gff_8_n58,
         keyFF_keystate_gff_8_n57, keyFF_keystate_gff_8_n56,
         keyFF_keystate_gff_8_n55, keyFF_keystate_gff_8_n54,
         keyFF_keystate_gff_8_n35, keyFF_keystate_gff_8_n34,
         keyFF_keystate_gff_8_n33, keyFF_keystate_gff_8_n32,
         keyFF_keystate_gff_8_n31, keyFF_keystate_gff_8_n30,
         keyFF_keystate_gff_8_n29, keyFF_keystate_gff_8_n28,
         keyFF_keystate_gff_9_n69, keyFF_keystate_gff_9_n68,
         keyFF_keystate_gff_9_n67, keyFF_keystate_gff_9_n66,
         keyFF_keystate_gff_9_n65, keyFF_keystate_gff_9_n64,
         keyFF_keystate_gff_9_n63, keyFF_keystate_gff_9_n62,
         keyFF_keystate_gff_9_n61, keyFF_keystate_gff_9_n60,
         keyFF_keystate_gff_9_n59, keyFF_keystate_gff_9_n58,
         keyFF_keystate_gff_9_n57, keyFF_keystate_gff_9_n56,
         keyFF_keystate_gff_9_n55, keyFF_keystate_gff_9_n36,
         keyFF_keystate_gff_9_n35, keyFF_keystate_gff_9_n34,
         keyFF_keystate_gff_9_n33, keyFF_keystate_gff_9_n32,
         keyFF_keystate_gff_9_n31, keyFF_keystate_gff_9_n30,
         keyFF_keystate_gff_9_n29, keyFF_keystate_gff_10_n69,
         keyFF_keystate_gff_10_n68, keyFF_keystate_gff_10_n67,
         keyFF_keystate_gff_10_n66, keyFF_keystate_gff_10_n65,
         keyFF_keystate_gff_10_n64, keyFF_keystate_gff_10_n63,
         keyFF_keystate_gff_10_n62, keyFF_keystate_gff_10_n61,
         keyFF_keystate_gff_10_n60, keyFF_keystate_gff_10_n59,
         keyFF_keystate_gff_10_n58, keyFF_keystate_gff_10_n57,
         keyFF_keystate_gff_10_n56, keyFF_keystate_gff_10_n55,
         keyFF_keystate_gff_10_n36, keyFF_keystate_gff_10_n35,
         keyFF_keystate_gff_10_n34, keyFF_keystate_gff_10_n33,
         keyFF_keystate_gff_10_n32, keyFF_keystate_gff_10_n31,
         keyFF_keystate_gff_10_n30, keyFF_keystate_gff_10_n29,
         keyFF_keystate_gff_11_n69, keyFF_keystate_gff_11_n68,
         keyFF_keystate_gff_11_n67, keyFF_keystate_gff_11_n66,
         keyFF_keystate_gff_11_n65, keyFF_keystate_gff_11_n64,
         keyFF_keystate_gff_11_n63, keyFF_keystate_gff_11_n62,
         keyFF_keystate_gff_11_n61, keyFF_keystate_gff_11_n60,
         keyFF_keystate_gff_11_n59, keyFF_keystate_gff_11_n58,
         keyFF_keystate_gff_11_n57, keyFF_keystate_gff_11_n56,
         keyFF_keystate_gff_11_n55, keyFF_keystate_gff_11_n36,
         keyFF_keystate_gff_11_n35, keyFF_keystate_gff_11_n34,
         keyFF_keystate_gff_11_n33, keyFF_keystate_gff_11_n32,
         keyFF_keystate_gff_11_n31, keyFF_keystate_gff_11_n30,
         keyFF_keystate_gff_11_n29, keyFF_keystate_gff_12_n69,
         keyFF_keystate_gff_12_n68, keyFF_keystate_gff_12_n67,
         keyFF_keystate_gff_12_n66, keyFF_keystate_gff_12_n65,
         keyFF_keystate_gff_12_n64, keyFF_keystate_gff_12_n63,
         keyFF_keystate_gff_12_n62, keyFF_keystate_gff_12_n61,
         keyFF_keystate_gff_12_n60, keyFF_keystate_gff_12_n59,
         keyFF_keystate_gff_12_n58, keyFF_keystate_gff_12_n57,
         keyFF_keystate_gff_12_n56, keyFF_keystate_gff_12_n55,
         keyFF_keystate_gff_12_n36, keyFF_keystate_gff_12_n35,
         keyFF_keystate_gff_12_n34, keyFF_keystate_gff_12_n33,
         keyFF_keystate_gff_12_n32, keyFF_keystate_gff_12_n31,
         keyFF_keystate_gff_12_n30, keyFF_keystate_gff_12_n29,
         keyFF_keystate_gff_13_n69, keyFF_keystate_gff_13_n68,
         keyFF_keystate_gff_13_n67, keyFF_keystate_gff_13_n66,
         keyFF_keystate_gff_13_n65, keyFF_keystate_gff_13_n64,
         keyFF_keystate_gff_13_n63, keyFF_keystate_gff_13_n62,
         keyFF_keystate_gff_13_n61, keyFF_keystate_gff_13_n60,
         keyFF_keystate_gff_13_n59, keyFF_keystate_gff_13_n58,
         keyFF_keystate_gff_13_n57, keyFF_keystate_gff_13_n56,
         keyFF_keystate_gff_13_n55, keyFF_keystate_gff_13_n36,
         keyFF_keystate_gff_13_n35, keyFF_keystate_gff_13_n34,
         keyFF_keystate_gff_13_n33, keyFF_keystate_gff_13_n32,
         keyFF_keystate_gff_13_n31, keyFF_keystate_gff_13_n30,
         keyFF_keystate_gff_13_n29, keyFF_keystate_gff_14_n69,
         keyFF_keystate_gff_14_n68, keyFF_keystate_gff_14_n67,
         keyFF_keystate_gff_14_n66, keyFF_keystate_gff_14_n65,
         keyFF_keystate_gff_14_n64, keyFF_keystate_gff_14_n63,
         keyFF_keystate_gff_14_n62, keyFF_keystate_gff_14_n61,
         keyFF_keystate_gff_14_n60, keyFF_keystate_gff_14_n59,
         keyFF_keystate_gff_14_n58, keyFF_keystate_gff_14_n57,
         keyFF_keystate_gff_14_n56, keyFF_keystate_gff_14_n55,
         keyFF_keystate_gff_14_n36, keyFF_keystate_gff_14_n35,
         keyFF_keystate_gff_14_n34, keyFF_keystate_gff_14_n33,
         keyFF_keystate_gff_14_n32, keyFF_keystate_gff_14_n31,
         keyFF_keystate_gff_14_n30, keyFF_keystate_gff_14_n29,
         keyFF_keystate_gff_15_n69, keyFF_keystate_gff_15_n68,
         keyFF_keystate_gff_15_n67, keyFF_keystate_gff_15_n66,
         keyFF_keystate_gff_15_n65, keyFF_keystate_gff_15_n64,
         keyFF_keystate_gff_15_n63, keyFF_keystate_gff_15_n62,
         keyFF_keystate_gff_15_n61, keyFF_keystate_gff_15_n60,
         keyFF_keystate_gff_15_n59, keyFF_keystate_gff_15_n58,
         keyFF_keystate_gff_15_n57, keyFF_keystate_gff_15_n56,
         keyFF_keystate_gff_15_n55, keyFF_keystate_gff_15_n36,
         keyFF_keystate_gff_15_n35, keyFF_keystate_gff_15_n34,
         keyFF_keystate_gff_15_n33, keyFF_keystate_gff_15_n32,
         keyFF_keystate_gff_15_n31, keyFF_keystate_gff_15_n30,
         keyFF_keystate_gff_15_n29, keyFF_keystate_gff_16_n69,
         keyFF_keystate_gff_16_n68, keyFF_keystate_gff_16_n67,
         keyFF_keystate_gff_16_n66, keyFF_keystate_gff_16_n65,
         keyFF_keystate_gff_16_n64, keyFF_keystate_gff_16_n63,
         keyFF_keystate_gff_16_n62, keyFF_keystate_gff_16_n61,
         keyFF_keystate_gff_16_n60, keyFF_keystate_gff_16_n59,
         keyFF_keystate_gff_16_n58, keyFF_keystate_gff_16_n57,
         keyFF_keystate_gff_16_n56, keyFF_keystate_gff_16_n55,
         keyFF_keystate_gff_16_n36, keyFF_keystate_gff_16_n35,
         keyFF_keystate_gff_16_n34, keyFF_keystate_gff_16_n33,
         keyFF_keystate_gff_16_n32, keyFF_keystate_gff_16_n31,
         keyFF_keystate_gff_16_n30, keyFF_keystate_gff_16_n29,
         keyFF_keystate_gff_17_n69, keyFF_keystate_gff_17_n68,
         keyFF_keystate_gff_17_n67, keyFF_keystate_gff_17_n66,
         keyFF_keystate_gff_17_n65, keyFF_keystate_gff_17_n64,
         keyFF_keystate_gff_17_n63, keyFF_keystate_gff_17_n62,
         keyFF_keystate_gff_17_n61, keyFF_keystate_gff_17_n60,
         keyFF_keystate_gff_17_n59, keyFF_keystate_gff_17_n58,
         keyFF_keystate_gff_17_n57, keyFF_keystate_gff_17_n56,
         keyFF_keystate_gff_17_n55, keyFF_keystate_gff_17_n36,
         keyFF_keystate_gff_17_n35, keyFF_keystate_gff_17_n34,
         keyFF_keystate_gff_17_n33, keyFF_keystate_gff_17_n32,
         keyFF_keystate_gff_17_n31, keyFF_keystate_gff_17_n30,
         keyFF_keystate_gff_17_n29, keyFF_keystate_gff_18_n69,
         keyFF_keystate_gff_18_n68, keyFF_keystate_gff_18_n67,
         keyFF_keystate_gff_18_n66, keyFF_keystate_gff_18_n65,
         keyFF_keystate_gff_18_n64, keyFF_keystate_gff_18_n63,
         keyFF_keystate_gff_18_n62, keyFF_keystate_gff_18_n61,
         keyFF_keystate_gff_18_n60, keyFF_keystate_gff_18_n59,
         keyFF_keystate_gff_18_n58, keyFF_keystate_gff_18_n57,
         keyFF_keystate_gff_18_n56, keyFF_keystate_gff_18_n55,
         keyFF_keystate_gff_18_n36, keyFF_keystate_gff_18_n35,
         keyFF_keystate_gff_18_n34, keyFF_keystate_gff_18_n33,
         keyFF_keystate_gff_18_n32, keyFF_keystate_gff_18_n31,
         keyFF_keystate_gff_18_n30, keyFF_keystate_gff_18_n29,
         keyFF_keystate_gff_19_n68, keyFF_keystate_gff_19_n67,
         keyFF_keystate_gff_19_n66, keyFF_keystate_gff_19_n65,
         keyFF_keystate_gff_19_n64, keyFF_keystate_gff_19_n63,
         keyFF_keystate_gff_19_n62, keyFF_keystate_gff_19_n61,
         keyFF_keystate_gff_19_n60, keyFF_keystate_gff_19_n59,
         keyFF_keystate_gff_19_n58, keyFF_keystate_gff_19_n57,
         keyFF_keystate_gff_19_n56, keyFF_keystate_gff_19_n55,
         keyFF_keystate_gff_19_n54, keyFF_keystate_gff_19_n35,
         keyFF_keystate_gff_19_n34, keyFF_keystate_gff_19_n33,
         keyFF_keystate_gff_19_n32, keyFF_keystate_gff_19_n31,
         keyFF_keystate_gff_19_n30, keyFF_keystate_gff_19_n29,
         keyFF_keystate_gff_19_n28, keyFF_keystate_gff_20_n68,
         keyFF_keystate_gff_20_n67, keyFF_keystate_gff_20_n66,
         keyFF_keystate_gff_20_n65, keyFF_keystate_gff_20_n64,
         keyFF_keystate_gff_20_n63, keyFF_keystate_gff_20_n62,
         keyFF_keystate_gff_20_n61, keyFF_keystate_gff_20_n60,
         keyFF_keystate_gff_20_n59, keyFF_keystate_gff_20_n58,
         keyFF_keystate_gff_20_n57, keyFF_keystate_gff_20_n56,
         keyFF_keystate_gff_20_n55, keyFF_keystate_gff_20_n54,
         keyFF_keystate_gff_20_n35, keyFF_keystate_gff_20_n34,
         keyFF_keystate_gff_20_n33, keyFF_keystate_gff_20_n32,
         keyFF_keystate_gff_20_n31, keyFF_keystate_gff_20_n30,
         keyFF_keystate_gff_20_n29, keyFF_keystate_gff_20_n28, sboxInst_n25,
         sboxInst_n24, sboxInst_n23, sboxInst_n22, sboxInst_n21, sboxInst_n20,
         sboxInst_n19, sboxInst_n18, sboxInst_n17, sboxInst_n16, sboxInst_n15,
         sboxInst_n14, sboxInst_n13, sboxInst_n12, sboxInst_n11, sboxInst_n10,
         sboxInst_n9, sboxInst_n8, sboxTI_f1_n13, sboxTI_f1_n12, sboxTI_f1_n11,
         sboxTI_f1_n10, sboxTI_f1_n9, sboxTI_f1_n8, sboxTI_f1_n7, sboxTI_f1_n6,
         sboxTI_f1_n5, sboxTI_f1_n4, sboxTI_f1_n3, sboxTI_f1_n2, sboxTI_f1_n1,
         sboxTI_f2_n11, sboxTI_f2_n10, sboxTI_f2_n9, sboxTI_f2_n8,
         sboxTI_f2_n7, sboxTI_f2_n6, sboxTI_f2_n5, sboxTI_f2_n4, sboxTI_f2_n3,
         sboxTI_f2_n2, sboxTI_f2_n1, sboxTI_f3_n13, sboxTI_f3_n12,
         sboxTI_f3_n11, sboxTI_f3_n10, sboxTI_f3_n9, sboxTI_f3_n8,
         sboxTI_f3_n7, sboxTI_f3_n6, sboxTI_f3_n5, sboxTI_f3_n4, sboxTI_f3_n3,
         sboxTI_f3_n2, sboxTI_f3_n1, sboxTI_g1_n22, sboxTI_g1_n21,
         sboxTI_g1_n20, sboxTI_g1_n19, sboxTI_g1_n18, sboxTI_g1_n17,
         sboxTI_g1_n16, sboxTI_g1_n15, sboxTI_g1_n14, sboxTI_g1_n13,
         sboxTI_g1_n12, sboxTI_g1_n11, sboxTI_g1_n10, sboxTI_g1_n9,
         sboxTI_g1_n8, sboxTI_g1_n7, sboxTI_g1_n6, sboxTI_g1_n5, sboxTI_g1_n4,
         sboxTI_g1_n3, sboxTI_g1_n2, sboxTI_g1_n1, sboxTI_g2_n23,
         sboxTI_g2_n22, sboxTI_g2_n21, sboxTI_g2_n20, sboxTI_g2_n19,
         sboxTI_g2_n18, sboxTI_g2_n17, sboxTI_g2_n16, sboxTI_g2_n15,
         sboxTI_g2_n14, sboxTI_g2_n13, sboxTI_g2_n12, sboxTI_g2_n11,
         sboxTI_g2_n10, sboxTI_g2_n9, sboxTI_g2_n8, sboxTI_g2_n7, sboxTI_g2_n6,
         sboxTI_g2_n5, sboxTI_g2_n4, sboxTI_g2_n3, sboxTI_g2_n2, sboxTI_g2_n1,
         sboxTI_g2_C, sboxTI_g3_n41, sboxTI_g3_n40, sboxTI_g3_n39,
         sboxTI_g3_n38, sboxTI_g3_n37, sboxTI_g3_n36, sboxTI_g3_n35,
         sboxTI_g3_n34, sboxTI_g3_n33, sboxTI_g3_n32, sboxTI_g3_n31,
         sboxTI_g3_n30, sboxTI_g3_n29, sboxTI_g3_n28, sboxTI_g3_n27,
         sboxTI_g3_n26, sboxTI_g3_n25, sboxTI_g3_n24, sboxTI_g3_n23,
         sboxTI_g3_n22, sboxTI_g3_n21, sboxTI_g3_n20, sboxTI_g3_C,
         sboxTI_y3_n13, sboxTI_y3_n12, sboxTI_y3_n11, sboxTI_y3_n10,
         sboxTI_y2_n17, sboxTI_y2_n16, sboxTI_y2_n15, sboxTI_y2_n14,
         sboxTI_y1_n17, sboxTI_y1_n16, sboxTI_y1_n15, sboxTI_y1_n14,
         DataOutReg1_gff_n200, DataOutReg1_gff_n199, DataOutReg1_gff_n198,
         DataOutReg1_gff_n193, DataOutReg1_gff_n192, DataOutReg1_gff_n191,
         DataOutReg1_gff_n190, DataOutReg1_gff_n189, DataOutReg1_gff_n188,
         DataOutReg1_gff_n187, DataOutReg1_gff_n186, DataOutReg1_gff_n185,
         DataOutReg1_gff_n184, DataOutReg1_gff_n183, DataOutReg1_gff_n182,
         DataOutReg1_gff_n181, DataOutReg1_gff_n180, DataOutReg1_gff_n179,
         DataOutReg1_gff_n178, DataOutReg1_gff_n177, DataOutReg1_gff_n176,
         DataOutReg1_gff_n175, DataOutReg1_gff_n174, DataOutReg1_gff_n173,
         DataOutReg1_gff_n172, DataOutReg1_gff_n171, DataOutReg1_gff_n170,
         DataOutReg1_gff_n169, DataOutReg1_gff_n168, DataOutReg1_gff_n167,
         DataOutReg1_gff_n166, DataOutReg1_gff_n165, DataOutReg1_gff_n164,
         DataOutReg1_gff_n163, DataOutReg1_gff_n162, DataOutReg1_gff_n161,
         DataOutReg1_gff_n160, DataOutReg1_gff_n159, DataOutReg1_gff_n158,
         DataOutReg1_gff_n157, DataOutReg1_gff_n156, DataOutReg1_gff_n155,
         DataOutReg1_gff_n154, DataOutReg1_gff_n153, DataOutReg1_gff_n152,
         DataOutReg1_gff_n151, DataOutReg1_gff_n150, DataOutReg1_gff_n149,
         DataOutReg1_gff_n148, DataOutReg1_gff_n147, DataOutReg1_gff_n146,
         DataOutReg1_gff_n145, DataOutReg1_gff_n144, DataOutReg1_gff_n143,
         DataOutReg1_gff_n142, DataOutReg1_gff_n141, DataOutReg1_gff_n140,
         DataOutReg1_gff_n139, DataOutReg1_gff_n138, DataOutReg1_gff_n137,
         DataOutReg1_gff_n136, DataOutReg1_gff_n135, DataOutReg1_gff_n134,
         DataOutReg1_gff_n133, DataOutReg1_gff_n132, DataOutReg1_gff_n131,
         DataOutReg1_gff_n130, DataOutReg2_gff_n392, DataOutReg2_gff_n391,
         DataOutReg2_gff_n262, DataOutReg2_gff_n261, DataOutReg2_gff_n260,
         DataOutReg2_gff_n259, DataOutReg2_gff_n258, DataOutReg2_gff_n257,
         DataOutReg2_gff_n256, DataOutReg2_gff_n255, DataOutReg2_gff_n254,
         DataOutReg2_gff_n253, DataOutReg2_gff_n252, DataOutReg2_gff_n251,
         DataOutReg2_gff_n250, DataOutReg2_gff_n249, DataOutReg2_gff_n248,
         DataOutReg2_gff_n247, DataOutReg2_gff_n246, DataOutReg2_gff_n245,
         DataOutReg2_gff_n244, DataOutReg2_gff_n243, DataOutReg2_gff_n242,
         DataOutReg2_gff_n241, DataOutReg2_gff_n240, DataOutReg2_gff_n239,
         DataOutReg2_gff_n238, DataOutReg2_gff_n237, DataOutReg2_gff_n236,
         DataOutReg2_gff_n235, DataOutReg2_gff_n234, DataOutReg2_gff_n233,
         DataOutReg2_gff_n232, DataOutReg2_gff_n231, DataOutReg2_gff_n230,
         DataOutReg2_gff_n229, DataOutReg2_gff_n228, DataOutReg2_gff_n227,
         DataOutReg2_gff_n226, DataOutReg2_gff_n225, DataOutReg2_gff_n224,
         DataOutReg2_gff_n223, DataOutReg2_gff_n222, DataOutReg2_gff_n221,
         DataOutReg2_gff_n220, DataOutReg2_gff_n219, DataOutReg2_gff_n218,
         DataOutReg2_gff_n217, DataOutReg2_gff_n216, DataOutReg2_gff_n215,
         DataOutReg2_gff_n214, DataOutReg2_gff_n213, DataOutReg2_gff_n212,
         DataOutReg2_gff_n211, DataOutReg2_gff_n210, DataOutReg2_gff_n209,
         DataOutReg2_gff_n208, DataOutReg2_gff_n207, DataOutReg2_gff_n206,
         DataOutReg2_gff_n205, DataOutReg2_gff_n204, DataOutReg2_gff_n203,
         DataOutReg2_gff_n202, DataOutReg2_gff_n201, DataOutReg2_gff_n200,
         DataOutReg2_gff_n199, DataOutReg3_gff_n393, DataOutReg3_gff_n392,
         DataOutReg3_gff_n391, DataOutReg3_gff_n262, DataOutReg3_gff_n261,
         DataOutReg3_gff_n260, DataOutReg3_gff_n259, DataOutReg3_gff_n258,
         DataOutReg3_gff_n257, DataOutReg3_gff_n256, DataOutReg3_gff_n255,
         DataOutReg3_gff_n254, DataOutReg3_gff_n253, DataOutReg3_gff_n252,
         DataOutReg3_gff_n251, DataOutReg3_gff_n250, DataOutReg3_gff_n249,
         DataOutReg3_gff_n248, DataOutReg3_gff_n247, DataOutReg3_gff_n246,
         DataOutReg3_gff_n245, DataOutReg3_gff_n244, DataOutReg3_gff_n243,
         DataOutReg3_gff_n242, DataOutReg3_gff_n241, DataOutReg3_gff_n240,
         DataOutReg3_gff_n239, DataOutReg3_gff_n238, DataOutReg3_gff_n237,
         DataOutReg3_gff_n236, DataOutReg3_gff_n235, DataOutReg3_gff_n234,
         DataOutReg3_gff_n233, DataOutReg3_gff_n232, DataOutReg3_gff_n231,
         DataOutReg3_gff_n230, DataOutReg3_gff_n229, DataOutReg3_gff_n228,
         DataOutReg3_gff_n227, DataOutReg3_gff_n226, DataOutReg3_gff_n225,
         DataOutReg3_gff_n224, DataOutReg3_gff_n223, DataOutReg3_gff_n222,
         DataOutReg3_gff_n221, DataOutReg3_gff_n220, DataOutReg3_gff_n219,
         DataOutReg3_gff_n218, DataOutReg3_gff_n217, DataOutReg3_gff_n216,
         DataOutReg3_gff_n215, DataOutReg3_gff_n214, DataOutReg3_gff_n213,
         DataOutReg3_gff_n212, DataOutReg3_gff_n211, DataOutReg3_gff_n210,
         DataOutReg3_gff_n209, DataOutReg3_gff_n208, DataOutReg3_gff_n207,
         DataOutReg3_gff_n206, DataOutReg3_gff_n205, DataOutReg3_gff_n204,
         DataOutReg3_gff_n203, DataOutReg3_gff_n202, DataOutReg3_gff_n201,
         DataOutReg3_gff_n200, DataOutReg3_gff_n199;
  wire   [2:0] ctrlData;
  wire   [4:0] counter;
  wire   [3:0] state;
  wire   [3:0] md1Reg;
  wire   [3:0] md2Reg;
  wire   [3:0] sboxOut;
  wire   [3:0] roundkey;
  wire   [3:1] keyRegKS;
  wire   [3:0] sboxIn1;
  wire   [3:0] fsm_countSerial;
  wire   [63:0] stateFF_permOut;
  wire   [63:0] stateFF_inputPar;
  wire   [63:0] md1FF_permOut;
  wire   [63:0] md1FF_inputPar;
  wire   [63:0] md2FF_permOut;
  wire   [63:0] md2FF_inputPar;
  wire   [75:3] keyFF_outputPar;
  wire   [79:0] keyFF_inputPar;
  wire   [3:0] sboxTI_g1Reg;
  wire   [3:0] sboxTI_g2Reg;
  wire   [3:0] sboxTI_g3Reg;
  wire   [3:0] sboxTI_g3Out;
  wire   [3:0] sboxTI_g2Out;
  wire   [3:0] sboxTI_g1Out;

  XOR2_X2 U9 ( .A(roundkey[2]), .B(state[2]), .Z(sboxIn1[2]) );
  XOR2_X1 U10 ( .A(roundkey[3]), .B(state[3]), .Z(sboxIn1[3]) );
  XOR2_X1 U11 ( .A(roundkey[0]), .B(state[0]), .Z(sboxIn1[0]) );
  XOR2_X1 U12 ( .A(roundkey[1]), .B(state[1]), .Z(sboxIn1[1]) );
  NOR2_X1 fsm_U40 ( .A1(reset), .A2(fsm_n34), .ZN(fsm_n43) );
  NOR2_X1 fsm_U39 ( .A1(final), .A2(fsm_n33), .ZN(fsm_n34) );
  NAND2_X1 fsm_U38 ( .A1(fsm_n32), .A2(fsm_n31), .ZN(fsm_n33) );
  NAND2_X1 fsm_U37 ( .A1(fsm_n7), .A2(fsm_n30), .ZN(fsm_n31) );
  NAND2_X1 fsm_U36 ( .A1(fsm_n29), .A2(fsm_en_countSerial), .ZN(fsm_n32) );
  NOR2_X1 fsm_U35 ( .A1(fsm_n8), .A2(fsm_n28), .ZN(final) );
  NAND2_X1 fsm_U34 ( .A1(fsm_n27), .A2(fsm_n26), .ZN(fsm_rst_countRound) );
  NOR2_X1 fsm_U33 ( .A1(reset), .A2(fsm_n25), .ZN(fsm_n41) );
  NOR2_X1 fsm_U32 ( .A1(enSboxReg), .A2(fsm_n24), .ZN(fsm_n25) );
  AND2_X1 fsm_U31 ( .A1(ctrlData[0]), .A2(fsm_n23), .ZN(fsm_n24) );
  NAND2_X1 fsm_U30 ( .A1(fsm_n22), .A2(fsm_n26), .ZN(fsm_rst_countSerial) );
  NAND2_X1 fsm_U29 ( .A1(fsm_n7), .A2(fsm_n35), .ZN(fsm_n26) );
  NOR2_X1 fsm_U28 ( .A1(fsm_n21), .A2(enSboxReg), .ZN(fsm_n22) );
  NOR2_X1 fsm_U27 ( .A1(reset), .A2(fsm_n20), .ZN(fsm_n42) );
  NOR2_X1 fsm_U26 ( .A1(fsm_n21), .A2(fsm_n19), .ZN(fsm_n20) );
  NOR2_X1 fsm_U25 ( .A1(fsm_n23), .A2(fsm_n18), .ZN(fsm_n19) );
  INV_X1 fsm_U24 ( .A(ctrlData[0]), .ZN(fsm_n18) );
  NAND2_X1 fsm_U23 ( .A1(counter[0]), .A2(fsm_n17), .ZN(fsm_n23) );
  NOR2_X1 fsm_U22 ( .A1(fsm_n16), .A2(fsm_n15), .ZN(fsm_n17) );
  NAND2_X1 fsm_U21 ( .A1(counter[2]), .A2(fsm_n14), .ZN(fsm_n15) );
  NOR2_X1 fsm_U20 ( .A1(fsm_n7), .A2(fsm_n13), .ZN(fsm_n14) );
  INV_X1 fsm_U19 ( .A(counter[4]), .ZN(fsm_n13) );
  NAND2_X1 fsm_U18 ( .A1(counter[1]), .A2(counter[3]), .ZN(fsm_n16) );
  INV_X1 fsm_U17 ( .A(fsm_n28), .ZN(fsm_n21) );
  AND2_X1 fsm_U16 ( .A1(fsm_n7), .A2(ctrlData[0]), .ZN(ctrlData[2]) );
  INV_X2 fsm_U15 ( .A(fsm_n27), .ZN(ctrlData[1]) );
  NOR2_X1 fsm_U14 ( .A1(fsm_en_countSerial), .A2(ctrlData[0]), .ZN(fsm_n27) );
  NOR2_X4 fsm_U13 ( .A1(fsm_n28), .A2(fsm_n35), .ZN(intDone) );
  AND2_X1 fsm_U12 ( .A1(enSboxReg), .A2(fsm_n29), .ZN(fsm_en_countRound) );
  NOR2_X1 fsm_U11 ( .A1(fsm_n12), .A2(fsm_n11), .ZN(fsm_n29) );
  NAND2_X1 fsm_U10 ( .A1(fsm_countSerial[0]), .A2(fsm_countSerial[1]), .ZN(
        fsm_n11) );
  NAND2_X1 fsm_U9 ( .A1(fsm_countSerial[2]), .A2(fsm_countSerial[3]), .ZN(
        fsm_n12) );
  NOR2_X2 fsm_U8 ( .A1(fsm_n7), .A2(fsm_n10), .ZN(enSboxReg) );
  INV_X1 fsm_U7 ( .A(fsm_n30), .ZN(fsm_n10) );
  NOR2_X4 fsm_U6 ( .A1(fsm_ps_state_2_), .A2(fsm_n8), .ZN(ctrlData[0]) );
  NAND2_X1 fsm_U5 ( .A1(fsm_ps_state_2_), .A2(fsm_n7), .ZN(fsm_n28) );
  OR2_X1 fsm_U4 ( .A1(enSboxReg), .A2(intDone), .ZN(fsm_en_countSerial) );
  NOR2_X1 fsm_U3 ( .A1(fsm_n35), .A2(fsm_ps_state_2_), .ZN(fsm_n30) );
DFF_X1 fsm_ps_state_reg_1_ ( .D(fsm_n41), .CK(clk), .Q(), .QN(fsm_n7) );
DFF_X1 fsm_ps_state_reg_2_ ( .D(fsm_n42), .CK(clk), .Q(fsm_ps_state_2_) , .QN() );
  DFF_X1 fsm_ps_state_reg_0_ ( .D(fsm_n43), .CK(clk), .Q(fsm_n35), .QN(fsm_n8)
         );
  NOR2_X1 fsm_cnt_rnd_U17 ( .A1(fsm_cnt_rnd_n34), .A2(fsm_cnt_rnd_n33), .ZN(
        fsm_cnt_rnd_n18) );
  XNOR2_X1 fsm_cnt_rnd_U16 ( .A(counter[0]), .B(fsm_en_countRound), .ZN(
        fsm_cnt_rnd_n34) );
  NOR2_X1 fsm_cnt_rnd_U15 ( .A1(fsm_cnt_rnd_n33), .A2(fsm_cnt_rnd_n32), .ZN(
        fsm_cnt_rnd_n17) );
  XOR2_X1 fsm_cnt_rnd_U14 ( .A(counter[1]), .B(fsm_cnt_rnd_n31), .Z(
        fsm_cnt_rnd_n32) );
  NOR2_X1 fsm_cnt_rnd_U13 ( .A1(fsm_cnt_rnd_n30), .A2(fsm_cnt_rnd_n33), .ZN(
        fsm_cnt_rnd_n16) );
  XNOR2_X1 fsm_cnt_rnd_U12 ( .A(fsm_cnt_rnd_n29), .B(counter[2]), .ZN(
        fsm_cnt_rnd_n30) );
  NOR2_X1 fsm_cnt_rnd_U11 ( .A1(fsm_cnt_rnd_n28), .A2(fsm_cnt_rnd_n33), .ZN(
        fsm_cnt_rnd_n15) );
  XNOR2_X1 fsm_cnt_rnd_U10 ( .A(fsm_cnt_rnd_n27), .B(fsm_cnt_rnd_n1), .ZN(
        fsm_cnt_rnd_n28) );
  NOR2_X1 fsm_cnt_rnd_U9 ( .A1(fsm_cnt_rnd_n26), .A2(fsm_cnt_rnd_n33), .ZN(
        fsm_cnt_rnd_n14) );
  INV_X1 fsm_cnt_rnd_U8 ( .A(fsm_rst_countRound), .ZN(fsm_cnt_rnd_n33) );
  XNOR2_X1 fsm_cnt_rnd_U7 ( .A(fsm_cnt_rnd_n25), .B(counter[4]), .ZN(
        fsm_cnt_rnd_n26) );
  NOR2_X1 fsm_cnt_rnd_U6 ( .A1(fsm_cnt_rnd_n1), .A2(fsm_cnt_rnd_n27), .ZN(
        fsm_cnt_rnd_n25) );
  NAND2_X1 fsm_cnt_rnd_U5 ( .A1(fsm_cnt_rnd_n29), .A2(counter[2]), .ZN(
        fsm_cnt_rnd_n27) );
  NOR2_X1 fsm_cnt_rnd_U4 ( .A1(fsm_cnt_rnd_n31), .A2(fsm_cnt_rnd_n35), .ZN(
        fsm_cnt_rnd_n29) );
  NAND2_X1 fsm_cnt_rnd_U3 ( .A1(counter[0]), .A2(fsm_en_countRound), .ZN(
        fsm_cnt_rnd_n31) );
  DFF_X1 fsm_cnt_rnd_count_reg_4_ ( .D(fsm_cnt_rnd_n14), .CK(clk), .Q(
        counter[4]) , .QN() ); 
  DFF_X1 fsm_cnt_rnd_count_reg_3_ ( .D(fsm_cnt_rnd_n15), .CK(clk), .Q(
        counter[3]), .QN(fsm_cnt_rnd_n1) );
  DFF_X1 fsm_cnt_rnd_count_reg_2_ ( .D(fsm_cnt_rnd_n16), .CK(clk), .Q(
        counter[2]) , .QN() ); 
  DFF_X1 fsm_cnt_rnd_count_reg_1_ ( .D(fsm_cnt_rnd_n17), .CK(clk), .Q(
        counter[1]), .QN(fsm_cnt_rnd_n35) );
  DFF_X1 fsm_cnt_rnd_count_reg_0_ ( .D(fsm_cnt_rnd_n18), .CK(clk), .Q(
        counter[0]) , .QN() ); 
  NOR2_X1 fsm_cnt_ser_U14 ( .A1(fsm_cnt_ser_n30), .A2(fsm_cnt_ser_n25), .ZN(
        fsm_cnt_ser_n26) );
  XNOR2_X1 fsm_cnt_ser_U13 ( .A(fsm_countSerial[3]), .B(fsm_cnt_ser_n24), .ZN(
        fsm_cnt_ser_n30) );
  NOR2_X1 fsm_cnt_ser_U12 ( .A1(fsm_cnt_ser_n1), .A2(fsm_cnt_ser_n23), .ZN(
        fsm_cnt_ser_n24) );
  NOR2_X1 fsm_cnt_ser_U11 ( .A1(fsm_cnt_ser_n25), .A2(fsm_cnt_ser_n22), .ZN(
        fsm_cnt_ser_n28) );
  XNOR2_X1 fsm_cnt_ser_U10 ( .A(fsm_cnt_ser_n3), .B(fsm_cnt_ser_n21), .ZN(
        fsm_cnt_ser_n22) );
  NOR2_X1 fsm_cnt_ser_U9 ( .A1(fsm_cnt_ser_n25), .A2(fsm_cnt_ser_n20), .ZN(
        fsm_cnt_ser_n27) );
  XNOR2_X1 fsm_cnt_ser_U8 ( .A(fsm_cnt_ser_n1), .B(fsm_cnt_ser_n23), .ZN(
        fsm_cnt_ser_n20) );
  OR2_X1 fsm_cnt_ser_U7 ( .A1(fsm_cnt_ser_n3), .A2(fsm_cnt_ser_n21), .ZN(
        fsm_cnt_ser_n23) );
  NAND2_X1 fsm_cnt_ser_U6 ( .A1(fsm_countSerial[0]), .A2(fsm_en_countSerial), 
        .ZN(fsm_cnt_ser_n21) );
  NOR2_X1 fsm_cnt_ser_U5 ( .A1(fsm_cnt_ser_n19), .A2(fsm_cnt_ser_n25), .ZN(
        fsm_cnt_ser_n29) );
  INV_X1 fsm_cnt_ser_U4 ( .A(fsm_rst_countSerial), .ZN(fsm_cnt_ser_n25) );
  XNOR2_X1 fsm_cnt_ser_U3 ( .A(fsm_countSerial[0]), .B(fsm_en_countSerial), 
        .ZN(fsm_cnt_ser_n19) );
  DFF_X1 fsm_cnt_ser_count_reg_3_ ( .D(fsm_cnt_ser_n26), .CK(clk), .Q(
        fsm_countSerial[3]) , .QN() ); 
  DFF_X1 fsm_cnt_ser_count_reg_2_ ( .D(fsm_cnt_ser_n27), .CK(clk), .Q(
        fsm_countSerial[2]), .QN(fsm_cnt_ser_n1) );
  DFF_X1 fsm_cnt_ser_count_reg_1_ ( .D(fsm_cnt_ser_n28), .CK(clk), .Q(
        fsm_countSerial[1]), .QN(fsm_cnt_ser_n3) );
  DFF_X1 fsm_cnt_ser_count_reg_0_ ( .D(fsm_cnt_ser_n29), .CK(clk), .Q(
        fsm_countSerial[0]) , .QN() ); 
  MUX2_X1 stateFF_U70 ( .A(stateFF_permOut[9]), .B(data_in1[9]), .S(
        stateFF_n139), .Z(stateFF_inputPar[9]) );
  MUX2_X1 stateFF_U69 ( .A(stateFF_permOut[8]), .B(data_in1[8]), .S(
        stateFF_n138), .Z(stateFF_inputPar[8]) );
  MUX2_X1 stateFF_U68 ( .A(stateFF_permOut[7]), .B(data_in1[7]), .S(
        stateFF_n139), .Z(stateFF_inputPar[7]) );
  MUX2_X1 stateFF_U67 ( .A(stateFF_permOut[6]), .B(data_in1[6]), .S(
        stateFF_n138), .Z(stateFF_inputPar[6]) );
  MUX2_X1 stateFF_U66 ( .A(stateFF_permOut[5]), .B(data_in1[5]), .S(
        stateFF_n137), .Z(stateFF_inputPar[5]) );
  MUX2_X1 stateFF_U65 ( .A(stateFF_permOut[4]), .B(data_in1[4]), .S(
        stateFF_n137), .Z(stateFF_inputPar[4]) );
  MUX2_X1 stateFF_U64 ( .A(stateFF_permOut[3]), .B(data_in1[3]), .S(
        stateFF_n137), .Z(stateFF_inputPar[3]) );
  MUX2_X1 stateFF_U63 ( .A(stateFF_permOut[2]), .B(data_in1[2]), .S(
        stateFF_n137), .Z(stateFF_inputPar[2]) );
  MUX2_X1 stateFF_U62 ( .A(stateFF_permOut[1]), .B(data_in1[1]), .S(
        stateFF_n137), .Z(stateFF_inputPar[1]) );
  MUX2_X1 stateFF_U61 ( .A(stateFF_permOut[0]), .B(data_in1[0]), .S(
        stateFF_n137), .Z(stateFF_inputPar[0]) );
  MUX2_X1 stateFF_U60 ( .A(stateFF_permOut[63]), .B(data_in1[63]), .S(
        stateFF_n137), .Z(stateFF_inputPar[63]) );
  MUX2_X1 stateFF_U59 ( .A(stateFF_permOut[62]), .B(data_in1[62]), .S(
        stateFF_n137), .Z(stateFF_inputPar[62]) );
  MUX2_X1 stateFF_U58 ( .A(stateFF_permOut[61]), .B(data_in1[61]), .S(
        stateFF_n137), .Z(stateFF_inputPar[61]) );
  MUX2_X1 stateFF_U57 ( .A(stateFF_permOut[60]), .B(data_in1[60]), .S(
        stateFF_n137), .Z(stateFF_inputPar[60]) );
  MUX2_X1 stateFF_U56 ( .A(stateFF_permOut[59]), .B(data_in1[59]), .S(
        stateFF_n137), .Z(stateFF_inputPar[59]) );
  MUX2_X1 stateFF_U55 ( .A(stateFF_permOut[58]), .B(data_in1[58]), .S(
        stateFF_n137), .Z(stateFF_inputPar[58]) );
  MUX2_X1 stateFF_U54 ( .A(stateFF_permOut[57]), .B(data_in1[57]), .S(
        stateFF_n139), .Z(stateFF_inputPar[57]) );
  MUX2_X1 stateFF_U53 ( .A(stateFF_permOut[56]), .B(data_in1[56]), .S(
        stateFF_n138), .Z(stateFF_inputPar[56]) );
  MUX2_X1 stateFF_U52 ( .A(stateFF_permOut[55]), .B(data_in1[55]), .S(
        stateFF_n139), .Z(stateFF_inputPar[55]) );
  MUX2_X1 stateFF_U51 ( .A(stateFF_permOut[54]), .B(data_in1[54]), .S(
        stateFF_n138), .Z(stateFF_inputPar[54]) );
  MUX2_X1 stateFF_U50 ( .A(stateFF_permOut[53]), .B(data_in1[53]), .S(
        stateFF_n139), .Z(stateFF_inputPar[53]) );
  MUX2_X1 stateFF_U49 ( .A(stateFF_permOut[52]), .B(data_in1[52]), .S(
        stateFF_n137), .Z(stateFF_inputPar[52]) );
  MUX2_X1 stateFF_U48 ( .A(stateFF_permOut[51]), .B(data_in1[51]), .S(
        stateFF_n136), .Z(stateFF_inputPar[51]) );
  MUX2_X1 stateFF_U47 ( .A(stateFF_permOut[50]), .B(data_in1[50]), .S(
        stateFF_n139), .Z(stateFF_inputPar[50]) );
  MUX2_X1 stateFF_U46 ( .A(stateFF_permOut[49]), .B(data_in1[49]), .S(
        stateFF_n138), .Z(stateFF_inputPar[49]) );
  MUX2_X1 stateFF_U45 ( .A(stateFF_permOut[48]), .B(data_in1[48]), .S(
        stateFF_n138), .Z(stateFF_inputPar[48]) );
  MUX2_X1 stateFF_U44 ( .A(stateFF_permOut[47]), .B(data_in1[47]), .S(
        stateFF_n137), .Z(stateFF_inputPar[47]) );
  INV_X1 stateFF_U43 ( .A(stateFF_n135), .ZN(stateFF_n137) );
  MUX2_X1 stateFF_U42 ( .A(stateFF_permOut[46]), .B(data_in1[46]), .S(
        stateFF_n136), .Z(stateFF_inputPar[46]) );
  MUX2_X1 stateFF_U41 ( .A(stateFF_permOut[45]), .B(data_in1[45]), .S(
        stateFF_n138), .Z(stateFF_inputPar[45]) );
  MUX2_X1 stateFF_U40 ( .A(stateFF_permOut[44]), .B(data_in1[44]), .S(
        stateFF_n138), .Z(stateFF_inputPar[44]) );
  MUX2_X1 stateFF_U39 ( .A(stateFF_permOut[43]), .B(data_in1[43]), .S(
        stateFF_n138), .Z(stateFF_inputPar[43]) );
  MUX2_X1 stateFF_U38 ( .A(stateFF_permOut[42]), .B(data_in1[42]), .S(
        stateFF_n138), .Z(stateFF_inputPar[42]) );
  MUX2_X1 stateFF_U37 ( .A(stateFF_permOut[41]), .B(data_in1[41]), .S(
        stateFF_n138), .Z(stateFF_inputPar[41]) );
  MUX2_X1 stateFF_U36 ( .A(stateFF_permOut[40]), .B(data_in1[40]), .S(
        stateFF_n138), .Z(stateFF_inputPar[40]) );
  MUX2_X1 stateFF_U35 ( .A(stateFF_permOut[39]), .B(data_in1[39]), .S(
        stateFF_n138), .Z(stateFF_inputPar[39]) );
  MUX2_X1 stateFF_U34 ( .A(stateFF_permOut[38]), .B(data_in1[38]), .S(
        stateFF_n138), .Z(stateFF_inputPar[38]) );
  MUX2_X1 stateFF_U33 ( .A(stateFF_permOut[37]), .B(data_in1[37]), .S(
        stateFF_n138), .Z(stateFF_inputPar[37]) );
  MUX2_X1 stateFF_U32 ( .A(stateFF_permOut[36]), .B(data_in1[36]), .S(
        stateFF_n138), .Z(stateFF_inputPar[36]) );
  MUX2_X1 stateFF_U31 ( .A(stateFF_permOut[35]), .B(data_in1[35]), .S(
        stateFF_n138), .Z(stateFF_inputPar[35]) );
  MUX2_X1 stateFF_U30 ( .A(stateFF_permOut[34]), .B(data_in1[34]), .S(
        stateFF_n138), .Z(stateFF_inputPar[34]) );
  INV_X1 stateFF_U29 ( .A(stateFF_n135), .ZN(stateFF_n138) );
  MUX2_X1 stateFF_U28 ( .A(stateFF_permOut[33]), .B(data_in1[33]), .S(
        stateFF_n139), .Z(stateFF_inputPar[33]) );
  MUX2_X1 stateFF_U27 ( .A(stateFF_permOut[32]), .B(data_in1[32]), .S(
        stateFF_n139), .Z(stateFF_inputPar[32]) );
  MUX2_X1 stateFF_U26 ( .A(stateFF_permOut[31]), .B(data_in1[31]), .S(
        stateFF_n139), .Z(stateFF_inputPar[31]) );
  MUX2_X1 stateFF_U25 ( .A(stateFF_permOut[30]), .B(data_in1[30]), .S(
        stateFF_n139), .Z(stateFF_inputPar[30]) );
  MUX2_X1 stateFF_U24 ( .A(stateFF_permOut[29]), .B(data_in1[29]), .S(
        stateFF_n139), .Z(stateFF_inputPar[29]) );
  MUX2_X1 stateFF_U23 ( .A(stateFF_permOut[28]), .B(data_in1[28]), .S(
        stateFF_n139), .Z(stateFF_inputPar[28]) );
  MUX2_X1 stateFF_U22 ( .A(stateFF_permOut[27]), .B(data_in1[27]), .S(
        stateFF_n139), .Z(stateFF_inputPar[27]) );
  MUX2_X1 stateFF_U21 ( .A(stateFF_permOut[26]), .B(data_in1[26]), .S(
        stateFF_n139), .Z(stateFF_inputPar[26]) );
  MUX2_X1 stateFF_U20 ( .A(stateFF_permOut[25]), .B(data_in1[25]), .S(
        stateFF_n139), .Z(stateFF_inputPar[25]) );
  MUX2_X1 stateFF_U19 ( .A(stateFF_permOut[24]), .B(data_in1[24]), .S(
        stateFF_n139), .Z(stateFF_inputPar[24]) );
  MUX2_X1 stateFF_U18 ( .A(stateFF_permOut[23]), .B(data_in1[23]), .S(
        stateFF_n139), .Z(stateFF_inputPar[23]) );
  MUX2_X1 stateFF_U17 ( .A(stateFF_permOut[22]), .B(data_in1[22]), .S(
        stateFF_n139), .Z(stateFF_inputPar[22]) );
  INV_X1 stateFF_U16 ( .A(stateFF_n135), .ZN(stateFF_n139) );
  MUX2_X1 stateFF_U15 ( .A(stateFF_permOut[21]), .B(data_in1[21]), .S(
        stateFF_n136), .Z(stateFF_inputPar[21]) );
  MUX2_X1 stateFF_U14 ( .A(stateFF_permOut[20]), .B(data_in1[20]), .S(
        stateFF_n136), .Z(stateFF_inputPar[20]) );
  MUX2_X1 stateFF_U13 ( .A(stateFF_permOut[19]), .B(data_in1[19]), .S(
        stateFF_n136), .Z(stateFF_inputPar[19]) );
  MUX2_X1 stateFF_U12 ( .A(stateFF_permOut[18]), .B(data_in1[18]), .S(
        stateFF_n136), .Z(stateFF_inputPar[18]) );
  MUX2_X1 stateFF_U11 ( .A(stateFF_permOut[17]), .B(data_in1[17]), .S(
        stateFF_n136), .Z(stateFF_inputPar[17]) );
  MUX2_X1 stateFF_U10 ( .A(stateFF_permOut[16]), .B(data_in1[16]), .S(
        stateFF_n136), .Z(stateFF_inputPar[16]) );
  MUX2_X1 stateFF_U9 ( .A(stateFF_permOut[15]), .B(data_in1[15]), .S(
        stateFF_n136), .Z(stateFF_inputPar[15]) );
  MUX2_X1 stateFF_U8 ( .A(stateFF_permOut[14]), .B(data_in1[14]), .S(
        stateFF_n136), .Z(stateFF_inputPar[14]) );
  MUX2_X1 stateFF_U7 ( .A(stateFF_permOut[13]), .B(data_in1[13]), .S(
        stateFF_n136), .Z(stateFF_inputPar[13]) );
  MUX2_X1 stateFF_U6 ( .A(stateFF_permOut[12]), .B(data_in1[12]), .S(
        stateFF_n136), .Z(stateFF_inputPar[12]) );
  MUX2_X1 stateFF_U5 ( .A(stateFF_permOut[11]), .B(data_in1[11]), .S(
        stateFF_n136), .Z(stateFF_inputPar[11]) );
  MUX2_X1 stateFF_U4 ( .A(stateFF_permOut[10]), .B(data_in1[10]), .S(
        stateFF_n136), .Z(stateFF_inputPar[10]) );
  INV_X1 stateFF_U3 ( .A(stateFF_n135), .ZN(stateFF_n136) );
  INV_X1 stateFF_U2 ( .A(ctrlData[2]), .ZN(stateFF_n135) );
  INV_X1 stateFF_state_U5 ( .A(ctrlData[1]), .ZN(stateFF_state_n8) );
  INV_X2 stateFF_state_U4 ( .A(stateFF_state_n11), .ZN(stateFF_state_n10) );
  INV_X2 stateFF_state_U3 ( .A(stateFF_state_n11), .ZN(stateFF_state_n9) );
  INV_X1 stateFF_state_U2 ( .A(ctrlData[0]), .ZN(stateFF_state_n11) );
  INV_X1 stateFF_state_U1 ( .A(stateFF_state_n8), .ZN(stateFF_state_n7) );
  NAND2_X1 stateFF_state_gff_1_U19 ( .A1(stateFF_state_gff_1_n41), .A2(
        stateFF_state_gff_1_n40), .ZN(stateFF_state_gff_1_n25) );
  NAND2_X1 stateFF_state_gff_1_U18 ( .A1(stateFF_state_gff_1_n39), .A2(
        stateFF_permOut[16]), .ZN(stateFF_state_gff_1_n40) );
  MUX2_X1 stateFF_state_gff_1_U17 ( .A(stateFF_state_gff_1_n21), .B(
        stateFF_state_gff_1_n38), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_1_n41) );
  NAND2_X1 stateFF_state_gff_1_U16 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[1]), .ZN(stateFF_state_gff_1_n38) );
  NAND2_X1 stateFF_state_gff_1_U15 ( .A1(stateFF_state_gff_1_n37), .A2(
        stateFF_state_gff_1_n36), .ZN(stateFF_state_gff_1_n27) );
  NAND2_X1 stateFF_state_gff_1_U14 ( .A1(stateFF_state_gff_1_n39), .A2(
        stateFF_permOut[48]), .ZN(stateFF_state_gff_1_n36) );
  MUX2_X1 stateFF_state_gff_1_U13 ( .A(stateFF_state_gff_1_n23), .B(
        stateFF_state_gff_1_n35), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_1_n37) );
  NAND2_X1 stateFF_state_gff_1_U12 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[3]), .ZN(stateFF_state_gff_1_n35) );
  NAND2_X1 stateFF_state_gff_1_U11 ( .A1(stateFF_state_gff_1_n34), .A2(
        stateFF_state_gff_1_n33), .ZN(stateFF_state_gff_1_n24) );
  NAND2_X1 stateFF_state_gff_1_U10 ( .A1(stateFF_state_gff_1_n39), .A2(
        stateFF_permOut[0]), .ZN(stateFF_state_gff_1_n33) );
  MUX2_X1 stateFF_state_gff_1_U9 ( .A(stateFF_state_gff_1_n20), .B(
        stateFF_state_gff_1_n32), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_1_n34) );
  NAND2_X1 stateFF_state_gff_1_U8 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[0]), .ZN(stateFF_state_gff_1_n32) );
  NAND2_X1 stateFF_state_gff_1_U7 ( .A1(stateFF_state_gff_1_n31), .A2(
        stateFF_state_gff_1_n30), .ZN(stateFF_state_gff_1_n26) );
  NAND2_X1 stateFF_state_gff_1_U6 ( .A1(stateFF_state_gff_1_n39), .A2(
        stateFF_permOut[32]), .ZN(stateFF_state_gff_1_n30) );
  NOR2_X1 stateFF_state_gff_1_U5 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_1_n29), .ZN(stateFF_state_gff_1_n39) );
  INV_X1 stateFF_state_gff_1_U4 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_1_n29) );
  MUX2_X1 stateFF_state_gff_1_U3 ( .A(stateFF_state_gff_1_n22), .B(
        stateFF_state_gff_1_n28), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_1_n31) );
  NAND2_X1 stateFF_state_gff_1_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[2]), .ZN(stateFF_state_gff_1_n28) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_1_n24), .CK(clk), .Q(stateFF_permOut[1]), .QN(
        stateFF_state_gff_1_n20) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_1_n25), .CK(clk), .Q(stateFF_permOut[17]), .QN(
        stateFF_state_gff_1_n21) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_1_n26), .CK(clk), .Q(stateFF_permOut[33]), .QN(
        stateFF_state_gff_1_n22) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_1_n27), .CK(clk), .Q(stateFF_permOut[49]), .QN(
        stateFF_state_gff_1_n23) );
  NAND2_X1 stateFF_state_gff_2_U19 ( .A1(stateFF_state_gff_2_n67), .A2(
        stateFF_state_gff_2_n66), .ZN(stateFF_state_gff_2_n28) );
  NAND2_X1 stateFF_state_gff_2_U18 ( .A1(stateFF_state_gff_2_n65), .A2(
        stateFF_permOut[49]), .ZN(stateFF_state_gff_2_n66) );
  MUX2_X1 stateFF_state_gff_2_U17 ( .A(stateFF_state_gff_2_n32), .B(
        stateFF_state_gff_2_n64), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_2_n67) );
  NAND2_X1 stateFF_state_gff_2_U16 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[7]), .ZN(stateFF_state_gff_2_n64) );
  NAND2_X1 stateFF_state_gff_2_U15 ( .A1(stateFF_state_gff_2_n63), .A2(
        stateFF_state_gff_2_n62), .ZN(stateFF_state_gff_2_n29) );
  NAND2_X1 stateFF_state_gff_2_U14 ( .A1(stateFF_state_gff_2_n65), .A2(
        stateFF_permOut[33]), .ZN(stateFF_state_gff_2_n62) );
  MUX2_X1 stateFF_state_gff_2_U13 ( .A(stateFF_state_gff_2_n33), .B(
        stateFF_state_gff_2_n61), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_2_n63) );
  NAND2_X1 stateFF_state_gff_2_U12 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[6]), .ZN(stateFF_state_gff_2_n61) );
  NAND2_X1 stateFF_state_gff_2_U11 ( .A1(stateFF_state_gff_2_n60), .A2(
        stateFF_state_gff_2_n59), .ZN(stateFF_state_gff_2_n30) );
  NAND2_X1 stateFF_state_gff_2_U10 ( .A1(stateFF_state_gff_2_n65), .A2(
        stateFF_permOut[17]), .ZN(stateFF_state_gff_2_n59) );
  MUX2_X1 stateFF_state_gff_2_U9 ( .A(stateFF_state_gff_2_n34), .B(
        stateFF_state_gff_2_n58), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_2_n60) );
  NAND2_X1 stateFF_state_gff_2_U8 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[5]), .ZN(stateFF_state_gff_2_n58) );
  NAND2_X1 stateFF_state_gff_2_U7 ( .A1(stateFF_state_gff_2_n57), .A2(
        stateFF_state_gff_2_n56), .ZN(stateFF_state_gff_2_n31) );
  NAND2_X1 stateFF_state_gff_2_U6 ( .A1(stateFF_state_gff_2_n65), .A2(
        stateFF_permOut[1]), .ZN(stateFF_state_gff_2_n56) );
  NOR2_X1 stateFF_state_gff_2_U5 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_2_n55), .ZN(stateFF_state_gff_2_n65) );
  INV_X1 stateFF_state_gff_2_U4 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_2_n55) );
  MUX2_X1 stateFF_state_gff_2_U3 ( .A(stateFF_state_gff_2_n35), .B(
        stateFF_state_gff_2_n54), .S(stateFF_state_n7), .Z(
        stateFF_state_gff_2_n57) );
  NAND2_X1 stateFF_state_gff_2_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[4]), .ZN(stateFF_state_gff_2_n54) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_2_n31), .CK(clk), .Q(stateFF_permOut[2]), .QN(
        stateFF_state_gff_2_n35) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_2_n30), .CK(clk), .Q(stateFF_permOut[18]), .QN(
        stateFF_state_gff_2_n34) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_2_n29), .CK(clk), .Q(stateFF_permOut[34]), .QN(
        stateFF_state_gff_2_n33) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_2_n28), .CK(clk), .Q(stateFF_permOut[50]), .QN(
        stateFF_state_gff_2_n32) );
  NAND2_X1 stateFF_state_gff_3_U20 ( .A1(stateFF_state_gff_3_n68), .A2(
        stateFF_state_gff_3_n67), .ZN(stateFF_state_gff_3_n30) );
  NAND2_X1 stateFF_state_gff_3_U19 ( .A1(stateFF_state_gff_3_n66), .A2(
        stateFF_permOut[18]), .ZN(stateFF_state_gff_3_n67) );
  MUX2_X1 stateFF_state_gff_3_U18 ( .A(stateFF_state_gff_3_n34), .B(
        stateFF_state_gff_3_n65), .S(stateFF_state_gff_3_n64), .Z(
        stateFF_state_gff_3_n68) );
  NAND2_X1 stateFF_state_gff_3_U17 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[9]), .ZN(stateFF_state_gff_3_n65) );
  NAND2_X1 stateFF_state_gff_3_U16 ( .A1(stateFF_state_gff_3_n63), .A2(
        stateFF_state_gff_3_n62), .ZN(stateFF_state_gff_3_n31) );
  NAND2_X1 stateFF_state_gff_3_U15 ( .A1(stateFF_state_gff_3_n66), .A2(
        stateFF_permOut[2]), .ZN(stateFF_state_gff_3_n62) );
  MUX2_X1 stateFF_state_gff_3_U14 ( .A(stateFF_state_gff_3_n35), .B(
        stateFF_state_gff_3_n61), .S(stateFF_state_gff_3_n64), .Z(
        stateFF_state_gff_3_n63) );
  NAND2_X1 stateFF_state_gff_3_U13 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[8]), .ZN(stateFF_state_gff_3_n61) );
  NAND2_X1 stateFF_state_gff_3_U12 ( .A1(stateFF_state_gff_3_n60), .A2(
        stateFF_state_gff_3_n59), .ZN(stateFF_state_gff_3_n28) );
  NAND2_X1 stateFF_state_gff_3_U11 ( .A1(stateFF_state_gff_3_n66), .A2(
        stateFF_permOut[50]), .ZN(stateFF_state_gff_3_n59) );
  MUX2_X1 stateFF_state_gff_3_U10 ( .A(stateFF_state_gff_3_n32), .B(
        stateFF_state_gff_3_n58), .S(stateFF_state_gff_3_n64), .Z(
        stateFF_state_gff_3_n60) );
  NAND2_X1 stateFF_state_gff_3_U9 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[11]), .ZN(stateFF_state_gff_3_n58) );
  NAND2_X1 stateFF_state_gff_3_U8 ( .A1(stateFF_state_gff_3_n57), .A2(
        stateFF_state_gff_3_n56), .ZN(stateFF_state_gff_3_n29) );
  NAND2_X1 stateFF_state_gff_3_U7 ( .A1(stateFF_state_gff_3_n66), .A2(
        stateFF_permOut[34]), .ZN(stateFF_state_gff_3_n56) );
  NOR2_X1 stateFF_state_gff_3_U6 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_3_n55), .ZN(stateFF_state_gff_3_n66) );
  MUX2_X1 stateFF_state_gff_3_U5 ( .A(stateFF_state_gff_3_n33), .B(
        stateFF_state_gff_3_n54), .S(stateFF_state_gff_3_n64), .Z(
        stateFF_state_gff_3_n57) );
  INV_X1 stateFF_state_gff_3_U4 ( .A(stateFF_state_gff_3_n55), .ZN(
        stateFF_state_gff_3_n64) );
  INV_X1 stateFF_state_gff_3_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_3_n55) );
  NAND2_X1 stateFF_state_gff_3_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[10]), .ZN(stateFF_state_gff_3_n54) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_3_n31), .CK(clk), .Q(stateFF_permOut[3]), .QN(
        stateFF_state_gff_3_n35) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_3_n30), .CK(clk), .Q(stateFF_permOut[19]), .QN(
        stateFF_state_gff_3_n34) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_3_n29), .CK(clk), .Q(stateFF_permOut[35]), .QN(
        stateFF_state_gff_3_n33) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_3_n28), .CK(clk), .Q(stateFF_permOut[51]), .QN(
        stateFF_state_gff_3_n32) );
  NAND2_X1 stateFF_state_gff_4_U20 ( .A1(stateFF_state_gff_4_n68), .A2(
        stateFF_state_gff_4_n67), .ZN(stateFF_state_gff_4_n28) );
  NAND2_X1 stateFF_state_gff_4_U19 ( .A1(stateFF_state_gff_4_n66), .A2(
        stateFF_permOut[51]), .ZN(stateFF_state_gff_4_n67) );
  MUX2_X1 stateFF_state_gff_4_U18 ( .A(stateFF_state_gff_4_n32), .B(
        stateFF_state_gff_4_n65), .S(stateFF_state_gff_4_n64), .Z(
        stateFF_state_gff_4_n68) );
  NAND2_X1 stateFF_state_gff_4_U17 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[15]), .ZN(stateFF_state_gff_4_n65) );
  NAND2_X1 stateFF_state_gff_4_U16 ( .A1(stateFF_state_gff_4_n63), .A2(
        stateFF_state_gff_4_n62), .ZN(stateFF_state_gff_4_n29) );
  NAND2_X1 stateFF_state_gff_4_U15 ( .A1(stateFF_state_gff_4_n66), .A2(
        stateFF_permOut[35]), .ZN(stateFF_state_gff_4_n62) );
  MUX2_X1 stateFF_state_gff_4_U14 ( .A(stateFF_state_gff_4_n33), .B(
        stateFF_state_gff_4_n61), .S(stateFF_state_gff_4_n64), .Z(
        stateFF_state_gff_4_n63) );
  NAND2_X1 stateFF_state_gff_4_U13 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[14]), .ZN(stateFF_state_gff_4_n61) );
  NAND2_X1 stateFF_state_gff_4_U12 ( .A1(stateFF_state_gff_4_n60), .A2(
        stateFF_state_gff_4_n59), .ZN(stateFF_state_gff_4_n30) );
  NAND2_X1 stateFF_state_gff_4_U11 ( .A1(stateFF_state_gff_4_n66), .A2(
        stateFF_permOut[19]), .ZN(stateFF_state_gff_4_n59) );
  MUX2_X1 stateFF_state_gff_4_U10 ( .A(stateFF_state_gff_4_n34), .B(
        stateFF_state_gff_4_n58), .S(stateFF_state_gff_4_n64), .Z(
        stateFF_state_gff_4_n60) );
  NAND2_X1 stateFF_state_gff_4_U9 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[13]), .ZN(stateFF_state_gff_4_n58) );
  NAND2_X1 stateFF_state_gff_4_U8 ( .A1(stateFF_state_gff_4_n57), .A2(
        stateFF_state_gff_4_n56), .ZN(stateFF_state_gff_4_n31) );
  NAND2_X1 stateFF_state_gff_4_U7 ( .A1(stateFF_state_gff_4_n66), .A2(
        stateFF_permOut[3]), .ZN(stateFF_state_gff_4_n56) );
  NOR2_X1 stateFF_state_gff_4_U6 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_4_n55), .ZN(stateFF_state_gff_4_n66) );
  MUX2_X1 stateFF_state_gff_4_U5 ( .A(stateFF_state_gff_4_n35), .B(
        stateFF_state_gff_4_n54), .S(stateFF_state_gff_4_n64), .Z(
        stateFF_state_gff_4_n57) );
  INV_X1 stateFF_state_gff_4_U4 ( .A(stateFF_state_gff_4_n55), .ZN(
        stateFF_state_gff_4_n64) );
  INV_X1 stateFF_state_gff_4_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_4_n55) );
  NAND2_X1 stateFF_state_gff_4_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[12]), .ZN(stateFF_state_gff_4_n54) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_4_n31), .CK(clk), .Q(stateFF_permOut[4]), .QN(
        stateFF_state_gff_4_n35) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_4_n30), .CK(clk), .Q(stateFF_permOut[20]), .QN(
        stateFF_state_gff_4_n34) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_4_n29), .CK(clk), .Q(stateFF_permOut[36]), .QN(
        stateFF_state_gff_4_n33) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_4_n28), .CK(clk), .Q(stateFF_permOut[52]), .QN(
        stateFF_state_gff_4_n32) );
  NAND2_X1 stateFF_state_gff_5_U20 ( .A1(stateFF_state_gff_5_n68), .A2(
        stateFF_state_gff_5_n67), .ZN(stateFF_state_gff_5_n28) );
  NAND2_X1 stateFF_state_gff_5_U19 ( .A1(stateFF_state_gff_5_n66), .A2(
        stateFF_permOut[52]), .ZN(stateFF_state_gff_5_n67) );
  MUX2_X1 stateFF_state_gff_5_U18 ( .A(stateFF_state_gff_5_n32), .B(
        stateFF_state_gff_5_n65), .S(stateFF_state_gff_5_n64), .Z(
        stateFF_state_gff_5_n68) );
  NAND2_X1 stateFF_state_gff_5_U17 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[19]), .ZN(stateFF_state_gff_5_n65) );
  NAND2_X1 stateFF_state_gff_5_U16 ( .A1(stateFF_state_gff_5_n63), .A2(
        stateFF_state_gff_5_n62), .ZN(stateFF_state_gff_5_n29) );
  NAND2_X1 stateFF_state_gff_5_U15 ( .A1(stateFF_state_gff_5_n66), .A2(
        stateFF_permOut[36]), .ZN(stateFF_state_gff_5_n62) );
  MUX2_X1 stateFF_state_gff_5_U14 ( .A(stateFF_state_gff_5_n33), .B(
        stateFF_state_gff_5_n61), .S(stateFF_state_gff_5_n64), .Z(
        stateFF_state_gff_5_n63) );
  NAND2_X1 stateFF_state_gff_5_U13 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[18]), .ZN(stateFF_state_gff_5_n61) );
  NAND2_X1 stateFF_state_gff_5_U12 ( .A1(stateFF_state_gff_5_n60), .A2(
        stateFF_state_gff_5_n59), .ZN(stateFF_state_gff_5_n30) );
  NAND2_X1 stateFF_state_gff_5_U11 ( .A1(stateFF_state_gff_5_n66), .A2(
        stateFF_permOut[20]), .ZN(stateFF_state_gff_5_n59) );
  MUX2_X1 stateFF_state_gff_5_U10 ( .A(stateFF_state_gff_5_n34), .B(
        stateFF_state_gff_5_n58), .S(stateFF_state_gff_5_n64), .Z(
        stateFF_state_gff_5_n60) );
  NAND2_X1 stateFF_state_gff_5_U9 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[17]), .ZN(stateFF_state_gff_5_n58) );
  NAND2_X1 stateFF_state_gff_5_U8 ( .A1(stateFF_state_gff_5_n57), .A2(
        stateFF_state_gff_5_n56), .ZN(stateFF_state_gff_5_n31) );
  NAND2_X1 stateFF_state_gff_5_U7 ( .A1(stateFF_state_gff_5_n66), .A2(
        stateFF_permOut[4]), .ZN(stateFF_state_gff_5_n56) );
  NOR2_X1 stateFF_state_gff_5_U6 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_5_n55), .ZN(stateFF_state_gff_5_n66) );
  MUX2_X1 stateFF_state_gff_5_U5 ( .A(stateFF_state_gff_5_n35), .B(
        stateFF_state_gff_5_n54), .S(stateFF_state_gff_5_n64), .Z(
        stateFF_state_gff_5_n57) );
  INV_X1 stateFF_state_gff_5_U4 ( .A(stateFF_state_gff_5_n55), .ZN(
        stateFF_state_gff_5_n64) );
  INV_X1 stateFF_state_gff_5_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_5_n55) );
  NAND2_X1 stateFF_state_gff_5_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[16]), .ZN(stateFF_state_gff_5_n54) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_5_n31), .CK(clk), .Q(stateFF_permOut[5]), .QN(
        stateFF_state_gff_5_n35) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_5_n30), .CK(clk), .Q(stateFF_permOut[21]), .QN(
        stateFF_state_gff_5_n34) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_5_n29), .CK(clk), .Q(stateFF_permOut[37]), .QN(
        stateFF_state_gff_5_n33) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_5_n28), .CK(clk), .Q(stateFF_permOut[53]), .QN(
        stateFF_state_gff_5_n32) );
  NAND2_X1 stateFF_state_gff_6_U20 ( .A1(stateFF_state_gff_6_n69), .A2(
        stateFF_state_gff_6_n68), .ZN(stateFF_state_gff_6_n29) );
  NAND2_X1 stateFF_state_gff_6_U19 ( .A1(stateFF_state_gff_6_n67), .A2(
        stateFF_permOut[53]), .ZN(stateFF_state_gff_6_n68) );
  MUX2_X1 stateFF_state_gff_6_U18 ( .A(stateFF_state_gff_6_n33), .B(
        stateFF_state_gff_6_n66), .S(stateFF_state_gff_6_n65), .Z(
        stateFF_state_gff_6_n69) );
  NAND2_X1 stateFF_state_gff_6_U17 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[23]), .ZN(stateFF_state_gff_6_n66) );
  NAND2_X1 stateFF_state_gff_6_U16 ( .A1(stateFF_state_gff_6_n64), .A2(
        stateFF_state_gff_6_n63), .ZN(stateFF_state_gff_6_n30) );
  NAND2_X1 stateFF_state_gff_6_U15 ( .A1(stateFF_state_gff_6_n67), .A2(
        stateFF_permOut[37]), .ZN(stateFF_state_gff_6_n63) );
  MUX2_X1 stateFF_state_gff_6_U14 ( .A(stateFF_state_gff_6_n34), .B(
        stateFF_state_gff_6_n62), .S(stateFF_state_gff_6_n65), .Z(
        stateFF_state_gff_6_n64) );
  NAND2_X1 stateFF_state_gff_6_U13 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[22]), .ZN(stateFF_state_gff_6_n62) );
  NAND2_X1 stateFF_state_gff_6_U12 ( .A1(stateFF_state_gff_6_n61), .A2(
        stateFF_state_gff_6_n60), .ZN(stateFF_state_gff_6_n31) );
  NAND2_X1 stateFF_state_gff_6_U11 ( .A1(stateFF_state_gff_6_n67), .A2(
        stateFF_permOut[21]), .ZN(stateFF_state_gff_6_n60) );
  MUX2_X1 stateFF_state_gff_6_U10 ( .A(stateFF_state_gff_6_n35), .B(
        stateFF_state_gff_6_n59), .S(stateFF_state_gff_6_n65), .Z(
        stateFF_state_gff_6_n61) );
  NAND2_X1 stateFF_state_gff_6_U9 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[21]), .ZN(stateFF_state_gff_6_n59) );
  NAND2_X1 stateFF_state_gff_6_U8 ( .A1(stateFF_state_gff_6_n58), .A2(
        stateFF_state_gff_6_n57), .ZN(stateFF_state_gff_6_n32) );
  NAND2_X1 stateFF_state_gff_6_U7 ( .A1(stateFF_state_gff_6_n67), .A2(
        stateFF_permOut[5]), .ZN(stateFF_state_gff_6_n57) );
  NOR2_X1 stateFF_state_gff_6_U6 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_6_n56), .ZN(stateFF_state_gff_6_n67) );
  MUX2_X1 stateFF_state_gff_6_U5 ( .A(stateFF_state_gff_6_n36), .B(
        stateFF_state_gff_6_n55), .S(stateFF_state_gff_6_n65), .Z(
        stateFF_state_gff_6_n58) );
  INV_X1 stateFF_state_gff_6_U4 ( .A(stateFF_state_gff_6_n56), .ZN(
        stateFF_state_gff_6_n65) );
  INV_X1 stateFF_state_gff_6_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_6_n56) );
  NAND2_X1 stateFF_state_gff_6_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[20]), .ZN(stateFF_state_gff_6_n55) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_6_n32), .CK(clk), .Q(stateFF_permOut[6]), .QN(
        stateFF_state_gff_6_n36) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_6_n31), .CK(clk), .Q(stateFF_permOut[22]), .QN(
        stateFF_state_gff_6_n35) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_6_n30), .CK(clk), .Q(stateFF_permOut[38]), .QN(
        stateFF_state_gff_6_n34) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_6_n29), .CK(clk), .Q(stateFF_permOut[54]), .QN(
        stateFF_state_gff_6_n33) );
  NAND2_X1 stateFF_state_gff_7_U20 ( .A1(stateFF_state_gff_7_n69), .A2(
        stateFF_state_gff_7_n68), .ZN(stateFF_state_gff_7_n29) );
  NAND2_X1 stateFF_state_gff_7_U19 ( .A1(stateFF_state_gff_7_n67), .A2(
        stateFF_permOut[54]), .ZN(stateFF_state_gff_7_n68) );
  MUX2_X1 stateFF_state_gff_7_U18 ( .A(stateFF_state_gff_7_n33), .B(
        stateFF_state_gff_7_n66), .S(stateFF_state_gff_7_n65), .Z(
        stateFF_state_gff_7_n69) );
  NAND2_X1 stateFF_state_gff_7_U17 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[27]), .ZN(stateFF_state_gff_7_n66) );
  NAND2_X1 stateFF_state_gff_7_U16 ( .A1(stateFF_state_gff_7_n64), .A2(
        stateFF_state_gff_7_n63), .ZN(stateFF_state_gff_7_n30) );
  NAND2_X1 stateFF_state_gff_7_U15 ( .A1(stateFF_state_gff_7_n67), .A2(
        stateFF_permOut[38]), .ZN(stateFF_state_gff_7_n63) );
  MUX2_X1 stateFF_state_gff_7_U14 ( .A(stateFF_state_gff_7_n34), .B(
        stateFF_state_gff_7_n62), .S(stateFF_state_gff_7_n65), .Z(
        stateFF_state_gff_7_n64) );
  NAND2_X1 stateFF_state_gff_7_U13 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[26]), .ZN(stateFF_state_gff_7_n62) );
  NAND2_X1 stateFF_state_gff_7_U12 ( .A1(stateFF_state_gff_7_n61), .A2(
        stateFF_state_gff_7_n60), .ZN(stateFF_state_gff_7_n31) );
  NAND2_X1 stateFF_state_gff_7_U11 ( .A1(stateFF_state_gff_7_n67), .A2(
        stateFF_permOut[22]), .ZN(stateFF_state_gff_7_n60) );
  MUX2_X1 stateFF_state_gff_7_U10 ( .A(stateFF_state_gff_7_n35), .B(
        stateFF_state_gff_7_n59), .S(stateFF_state_gff_7_n65), .Z(
        stateFF_state_gff_7_n61) );
  NAND2_X1 stateFF_state_gff_7_U9 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[25]), .ZN(stateFF_state_gff_7_n59) );
  NAND2_X1 stateFF_state_gff_7_U8 ( .A1(stateFF_state_gff_7_n58), .A2(
        stateFF_state_gff_7_n57), .ZN(stateFF_state_gff_7_n32) );
  NAND2_X1 stateFF_state_gff_7_U7 ( .A1(stateFF_state_gff_7_n67), .A2(
        stateFF_permOut[6]), .ZN(stateFF_state_gff_7_n57) );
  NOR2_X1 stateFF_state_gff_7_U6 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_7_n56), .ZN(stateFF_state_gff_7_n67) );
  MUX2_X1 stateFF_state_gff_7_U5 ( .A(stateFF_state_gff_7_n36), .B(
        stateFF_state_gff_7_n55), .S(stateFF_state_gff_7_n65), .Z(
        stateFF_state_gff_7_n58) );
  INV_X1 stateFF_state_gff_7_U4 ( .A(stateFF_state_gff_7_n56), .ZN(
        stateFF_state_gff_7_n65) );
  INV_X1 stateFF_state_gff_7_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_7_n56) );
  NAND2_X1 stateFF_state_gff_7_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[24]), .ZN(stateFF_state_gff_7_n55) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_7_n32), .CK(clk), .Q(stateFF_permOut[7]), .QN(
        stateFF_state_gff_7_n36) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_7_n31), .CK(clk), .Q(stateFF_permOut[23]), .QN(
        stateFF_state_gff_7_n35) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_7_n30), .CK(clk), .Q(stateFF_permOut[39]), .QN(
        stateFF_state_gff_7_n34) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_7_n29), .CK(clk), .Q(stateFF_permOut[55]), .QN(
        stateFF_state_gff_7_n33) );
  NAND2_X1 stateFF_state_gff_8_U20 ( .A1(stateFF_state_gff_8_n69), .A2(
        stateFF_state_gff_8_n68), .ZN(stateFF_state_gff_8_n29) );
  NAND2_X1 stateFF_state_gff_8_U19 ( .A1(stateFF_state_gff_8_n67), .A2(
        stateFF_permOut[55]), .ZN(stateFF_state_gff_8_n68) );
  MUX2_X1 stateFF_state_gff_8_U18 ( .A(stateFF_state_gff_8_n33), .B(
        stateFF_state_gff_8_n66), .S(stateFF_state_gff_8_n65), .Z(
        stateFF_state_gff_8_n69) );
  NAND2_X1 stateFF_state_gff_8_U17 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[31]), .ZN(stateFF_state_gff_8_n66) );
  NAND2_X1 stateFF_state_gff_8_U16 ( .A1(stateFF_state_gff_8_n64), .A2(
        stateFF_state_gff_8_n63), .ZN(stateFF_state_gff_8_n30) );
  NAND2_X1 stateFF_state_gff_8_U15 ( .A1(stateFF_state_gff_8_n67), .A2(
        stateFF_permOut[39]), .ZN(stateFF_state_gff_8_n63) );
  MUX2_X1 stateFF_state_gff_8_U14 ( .A(stateFF_state_gff_8_n34), .B(
        stateFF_state_gff_8_n62), .S(stateFF_state_gff_8_n65), .Z(
        stateFF_state_gff_8_n64) );
  NAND2_X1 stateFF_state_gff_8_U13 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[30]), .ZN(stateFF_state_gff_8_n62) );
  NAND2_X1 stateFF_state_gff_8_U12 ( .A1(stateFF_state_gff_8_n61), .A2(
        stateFF_state_gff_8_n60), .ZN(stateFF_state_gff_8_n31) );
  NAND2_X1 stateFF_state_gff_8_U11 ( .A1(stateFF_state_gff_8_n67), .A2(
        stateFF_permOut[23]), .ZN(stateFF_state_gff_8_n60) );
  MUX2_X1 stateFF_state_gff_8_U10 ( .A(stateFF_state_gff_8_n35), .B(
        stateFF_state_gff_8_n59), .S(stateFF_state_gff_8_n65), .Z(
        stateFF_state_gff_8_n61) );
  NAND2_X1 stateFF_state_gff_8_U9 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[29]), .ZN(stateFF_state_gff_8_n59) );
  NAND2_X1 stateFF_state_gff_8_U8 ( .A1(stateFF_state_gff_8_n58), .A2(
        stateFF_state_gff_8_n57), .ZN(stateFF_state_gff_8_n32) );
  NAND2_X1 stateFF_state_gff_8_U7 ( .A1(stateFF_state_gff_8_n67), .A2(
        stateFF_permOut[7]), .ZN(stateFF_state_gff_8_n57) );
  NOR2_X1 stateFF_state_gff_8_U6 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_8_n56), .ZN(stateFF_state_gff_8_n67) );
  MUX2_X1 stateFF_state_gff_8_U5 ( .A(stateFF_state_gff_8_n36), .B(
        stateFF_state_gff_8_n55), .S(stateFF_state_gff_8_n65), .Z(
        stateFF_state_gff_8_n58) );
  INV_X1 stateFF_state_gff_8_U4 ( .A(stateFF_state_gff_8_n56), .ZN(
        stateFF_state_gff_8_n65) );
  INV_X1 stateFF_state_gff_8_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_8_n56) );
  NAND2_X1 stateFF_state_gff_8_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[28]), .ZN(stateFF_state_gff_8_n55) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_8_n32), .CK(clk), .Q(stateFF_permOut[8]), .QN(
        stateFF_state_gff_8_n36) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_8_n31), .CK(clk), .Q(stateFF_permOut[24]), .QN(
        stateFF_state_gff_8_n35) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_8_n30), .CK(clk), .Q(stateFF_permOut[40]), .QN(
        stateFF_state_gff_8_n34) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_8_n29), .CK(clk), .Q(stateFF_permOut[56]), .QN(
        stateFF_state_gff_8_n33) );
  NAND2_X1 stateFF_state_gff_9_U20 ( .A1(stateFF_state_gff_9_n69), .A2(
        stateFF_state_gff_9_n68), .ZN(stateFF_state_gff_9_n29) );
  NAND2_X1 stateFF_state_gff_9_U19 ( .A1(stateFF_state_gff_9_n67), .A2(
        stateFF_permOut[56]), .ZN(stateFF_state_gff_9_n68) );
  MUX2_X1 stateFF_state_gff_9_U18 ( .A(stateFF_state_gff_9_n33), .B(
        stateFF_state_gff_9_n66), .S(stateFF_state_gff_9_n65), .Z(
        stateFF_state_gff_9_n69) );
  NAND2_X1 stateFF_state_gff_9_U17 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[35]), .ZN(stateFF_state_gff_9_n66) );
  NAND2_X1 stateFF_state_gff_9_U16 ( .A1(stateFF_state_gff_9_n64), .A2(
        stateFF_state_gff_9_n63), .ZN(stateFF_state_gff_9_n30) );
  NAND2_X1 stateFF_state_gff_9_U15 ( .A1(stateFF_state_gff_9_n67), .A2(
        stateFF_permOut[40]), .ZN(stateFF_state_gff_9_n63) );
  MUX2_X1 stateFF_state_gff_9_U14 ( .A(stateFF_state_gff_9_n34), .B(
        stateFF_state_gff_9_n62), .S(stateFF_state_gff_9_n65), .Z(
        stateFF_state_gff_9_n64) );
  NAND2_X1 stateFF_state_gff_9_U13 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[34]), .ZN(stateFF_state_gff_9_n62) );
  NAND2_X1 stateFF_state_gff_9_U12 ( .A1(stateFF_state_gff_9_n61), .A2(
        stateFF_state_gff_9_n60), .ZN(stateFF_state_gff_9_n31) );
  NAND2_X1 stateFF_state_gff_9_U11 ( .A1(stateFF_state_gff_9_n67), .A2(
        stateFF_permOut[24]), .ZN(stateFF_state_gff_9_n60) );
  MUX2_X1 stateFF_state_gff_9_U10 ( .A(stateFF_state_gff_9_n35), .B(
        stateFF_state_gff_9_n59), .S(stateFF_state_gff_9_n65), .Z(
        stateFF_state_gff_9_n61) );
  NAND2_X1 stateFF_state_gff_9_U9 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[33]), .ZN(stateFF_state_gff_9_n59) );
  NAND2_X1 stateFF_state_gff_9_U8 ( .A1(stateFF_state_gff_9_n58), .A2(
        stateFF_state_gff_9_n57), .ZN(stateFF_state_gff_9_n32) );
  NAND2_X1 stateFF_state_gff_9_U7 ( .A1(stateFF_state_gff_9_n67), .A2(
        stateFF_permOut[8]), .ZN(stateFF_state_gff_9_n57) );
  NOR2_X1 stateFF_state_gff_9_U6 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_9_n56), .ZN(stateFF_state_gff_9_n67) );
  MUX2_X1 stateFF_state_gff_9_U5 ( .A(stateFF_state_gff_9_n36), .B(
        stateFF_state_gff_9_n55), .S(stateFF_state_gff_9_n65), .Z(
        stateFF_state_gff_9_n58) );
  INV_X1 stateFF_state_gff_9_U4 ( .A(stateFF_state_gff_9_n56), .ZN(
        stateFF_state_gff_9_n65) );
  INV_X1 stateFF_state_gff_9_U3 ( .A(ctrlData[1]), .ZN(stateFF_state_gff_9_n56) );
  NAND2_X1 stateFF_state_gff_9_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[32]), .ZN(stateFF_state_gff_9_n55) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_9_n32), .CK(clk), .Q(stateFF_permOut[9]), .QN(
        stateFF_state_gff_9_n36) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_9_n31), .CK(clk), .Q(stateFF_permOut[25]), .QN(
        stateFF_state_gff_9_n35) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_9_n30), .CK(clk), .Q(stateFF_permOut[41]), .QN(
        stateFF_state_gff_9_n34) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_9_n29), .CK(clk), .Q(stateFF_permOut[57]), .QN(
        stateFF_state_gff_9_n33) );
  NAND2_X1 stateFF_state_gff_10_U20 ( .A1(stateFF_state_gff_10_n69), .A2(
        stateFF_state_gff_10_n68), .ZN(stateFF_state_gff_10_n29) );
  NAND2_X1 stateFF_state_gff_10_U19 ( .A1(stateFF_state_gff_10_n67), .A2(
        stateFF_permOut[57]), .ZN(stateFF_state_gff_10_n68) );
  MUX2_X1 stateFF_state_gff_10_U18 ( .A(stateFF_state_gff_10_n33), .B(
        stateFF_state_gff_10_n66), .S(stateFF_state_gff_10_n65), .Z(
        stateFF_state_gff_10_n69) );
  NAND2_X1 stateFF_state_gff_10_U17 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[39]), .ZN(stateFF_state_gff_10_n66) );
  NAND2_X1 stateFF_state_gff_10_U16 ( .A1(stateFF_state_gff_10_n64), .A2(
        stateFF_state_gff_10_n63), .ZN(stateFF_state_gff_10_n30) );
  NAND2_X1 stateFF_state_gff_10_U15 ( .A1(stateFF_state_gff_10_n67), .A2(
        stateFF_permOut[41]), .ZN(stateFF_state_gff_10_n63) );
  MUX2_X1 stateFF_state_gff_10_U14 ( .A(stateFF_state_gff_10_n34), .B(
        stateFF_state_gff_10_n62), .S(stateFF_state_gff_10_n65), .Z(
        stateFF_state_gff_10_n64) );
  NAND2_X1 stateFF_state_gff_10_U13 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[38]), .ZN(stateFF_state_gff_10_n62) );
  NAND2_X1 stateFF_state_gff_10_U12 ( .A1(stateFF_state_gff_10_n61), .A2(
        stateFF_state_gff_10_n60), .ZN(stateFF_state_gff_10_n31) );
  NAND2_X1 stateFF_state_gff_10_U11 ( .A1(stateFF_state_gff_10_n67), .A2(
        stateFF_permOut[25]), .ZN(stateFF_state_gff_10_n60) );
  MUX2_X1 stateFF_state_gff_10_U10 ( .A(stateFF_state_gff_10_n35), .B(
        stateFF_state_gff_10_n59), .S(stateFF_state_gff_10_n65), .Z(
        stateFF_state_gff_10_n61) );
  NAND2_X1 stateFF_state_gff_10_U9 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[37]), .ZN(stateFF_state_gff_10_n59) );
  NAND2_X1 stateFF_state_gff_10_U8 ( .A1(stateFF_state_gff_10_n58), .A2(
        stateFF_state_gff_10_n57), .ZN(stateFF_state_gff_10_n32) );
  NAND2_X1 stateFF_state_gff_10_U7 ( .A1(stateFF_state_gff_10_n67), .A2(
        stateFF_permOut[9]), .ZN(stateFF_state_gff_10_n57) );
  NOR2_X1 stateFF_state_gff_10_U6 ( .A1(stateFF_state_n10), .A2(
        stateFF_state_gff_10_n56), .ZN(stateFF_state_gff_10_n67) );
  MUX2_X1 stateFF_state_gff_10_U5 ( .A(stateFF_state_gff_10_n36), .B(
        stateFF_state_gff_10_n55), .S(stateFF_state_gff_10_n65), .Z(
        stateFF_state_gff_10_n58) );
  INV_X1 stateFF_state_gff_10_U4 ( .A(stateFF_state_gff_10_n56), .ZN(
        stateFF_state_gff_10_n65) );
  INV_X1 stateFF_state_gff_10_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_10_n56) );
  NAND2_X1 stateFF_state_gff_10_U2 ( .A1(stateFF_state_n10), .A2(
        stateFF_inputPar[36]), .ZN(stateFF_state_gff_10_n55) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_10_n32), .CK(clk), .Q(stateFF_permOut[10]), .QN(
        stateFF_state_gff_10_n36) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_10_n31), .CK(clk), .Q(stateFF_permOut[26]), .QN(
        stateFF_state_gff_10_n35) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_10_n30), .CK(clk), .Q(stateFF_permOut[42]), .QN(
        stateFF_state_gff_10_n34) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_10_n29), .CK(clk), .Q(stateFF_permOut[58]), .QN(
        stateFF_state_gff_10_n33) );
  NAND2_X1 stateFF_state_gff_11_U20 ( .A1(stateFF_state_gff_11_n69), .A2(
        stateFF_state_gff_11_n68), .ZN(stateFF_state_gff_11_n29) );
  NAND2_X1 stateFF_state_gff_11_U19 ( .A1(stateFF_state_gff_11_n67), .A2(
        stateFF_permOut[58]), .ZN(stateFF_state_gff_11_n68) );
  MUX2_X1 stateFF_state_gff_11_U18 ( .A(stateFF_state_gff_11_n33), .B(
        stateFF_state_gff_11_n66), .S(stateFF_state_gff_11_n65), .Z(
        stateFF_state_gff_11_n69) );
  NAND2_X1 stateFF_state_gff_11_U17 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[43]), .ZN(stateFF_state_gff_11_n66) );
  NAND2_X1 stateFF_state_gff_11_U16 ( .A1(stateFF_state_gff_11_n64), .A2(
        stateFF_state_gff_11_n63), .ZN(stateFF_state_gff_11_n30) );
  NAND2_X1 stateFF_state_gff_11_U15 ( .A1(stateFF_state_gff_11_n67), .A2(
        stateFF_permOut[42]), .ZN(stateFF_state_gff_11_n63) );
  MUX2_X1 stateFF_state_gff_11_U14 ( .A(stateFF_state_gff_11_n34), .B(
        stateFF_state_gff_11_n62), .S(stateFF_state_gff_11_n65), .Z(
        stateFF_state_gff_11_n64) );
  NAND2_X1 stateFF_state_gff_11_U13 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[42]), .ZN(stateFF_state_gff_11_n62) );
  NAND2_X1 stateFF_state_gff_11_U12 ( .A1(stateFF_state_gff_11_n61), .A2(
        stateFF_state_gff_11_n60), .ZN(stateFF_state_gff_11_n31) );
  NAND2_X1 stateFF_state_gff_11_U11 ( .A1(stateFF_state_gff_11_n67), .A2(
        stateFF_permOut[26]), .ZN(stateFF_state_gff_11_n60) );
  MUX2_X1 stateFF_state_gff_11_U10 ( .A(stateFF_state_gff_11_n35), .B(
        stateFF_state_gff_11_n59), .S(stateFF_state_gff_11_n65), .Z(
        stateFF_state_gff_11_n61) );
  NAND2_X1 stateFF_state_gff_11_U9 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[41]), .ZN(stateFF_state_gff_11_n59) );
  NAND2_X1 stateFF_state_gff_11_U8 ( .A1(stateFF_state_gff_11_n58), .A2(
        stateFF_state_gff_11_n57), .ZN(stateFF_state_gff_11_n32) );
  NAND2_X1 stateFF_state_gff_11_U7 ( .A1(stateFF_state_gff_11_n67), .A2(
        stateFF_permOut[10]), .ZN(stateFF_state_gff_11_n57) );
  NOR2_X1 stateFF_state_gff_11_U6 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_11_n56), .ZN(stateFF_state_gff_11_n67) );
  MUX2_X1 stateFF_state_gff_11_U5 ( .A(stateFF_state_gff_11_n36), .B(
        stateFF_state_gff_11_n55), .S(stateFF_state_gff_11_n65), .Z(
        stateFF_state_gff_11_n58) );
  INV_X1 stateFF_state_gff_11_U4 ( .A(stateFF_state_gff_11_n56), .ZN(
        stateFF_state_gff_11_n65) );
  INV_X1 stateFF_state_gff_11_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_11_n56) );
  NAND2_X1 stateFF_state_gff_11_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[40]), .ZN(stateFF_state_gff_11_n55) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_11_n32), .CK(clk), .Q(stateFF_permOut[11]), .QN(
        stateFF_state_gff_11_n36) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_11_n31), .CK(clk), .Q(stateFF_permOut[27]), .QN(
        stateFF_state_gff_11_n35) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_11_n30), .CK(clk), .Q(stateFF_permOut[43]), .QN(
        stateFF_state_gff_11_n34) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_11_n29), .CK(clk), .Q(stateFF_permOut[59]), .QN(
        stateFF_state_gff_11_n33) );
  NAND2_X1 stateFF_state_gff_12_U20 ( .A1(stateFF_state_gff_12_n69), .A2(
        stateFF_state_gff_12_n68), .ZN(stateFF_state_gff_12_n29) );
  NAND2_X1 stateFF_state_gff_12_U19 ( .A1(stateFF_state_gff_12_n67), .A2(
        stateFF_permOut[59]), .ZN(stateFF_state_gff_12_n68) );
  MUX2_X1 stateFF_state_gff_12_U18 ( .A(stateFF_state_gff_12_n33), .B(
        stateFF_state_gff_12_n66), .S(stateFF_state_gff_12_n65), .Z(
        stateFF_state_gff_12_n69) );
  NAND2_X1 stateFF_state_gff_12_U17 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[47]), .ZN(stateFF_state_gff_12_n66) );
  NAND2_X1 stateFF_state_gff_12_U16 ( .A1(stateFF_state_gff_12_n64), .A2(
        stateFF_state_gff_12_n63), .ZN(stateFF_state_gff_12_n30) );
  NAND2_X1 stateFF_state_gff_12_U15 ( .A1(stateFF_state_gff_12_n67), .A2(
        stateFF_permOut[43]), .ZN(stateFF_state_gff_12_n63) );
  MUX2_X1 stateFF_state_gff_12_U14 ( .A(stateFF_state_gff_12_n34), .B(
        stateFF_state_gff_12_n62), .S(stateFF_state_gff_12_n65), .Z(
        stateFF_state_gff_12_n64) );
  NAND2_X1 stateFF_state_gff_12_U13 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[46]), .ZN(stateFF_state_gff_12_n62) );
  NAND2_X1 stateFF_state_gff_12_U12 ( .A1(stateFF_state_gff_12_n61), .A2(
        stateFF_state_gff_12_n60), .ZN(stateFF_state_gff_12_n31) );
  NAND2_X1 stateFF_state_gff_12_U11 ( .A1(stateFF_state_gff_12_n67), .A2(
        stateFF_permOut[27]), .ZN(stateFF_state_gff_12_n60) );
  MUX2_X1 stateFF_state_gff_12_U10 ( .A(stateFF_state_gff_12_n35), .B(
        stateFF_state_gff_12_n59), .S(stateFF_state_gff_12_n65), .Z(
        stateFF_state_gff_12_n61) );
  NAND2_X1 stateFF_state_gff_12_U9 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[45]), .ZN(stateFF_state_gff_12_n59) );
  NAND2_X1 stateFF_state_gff_12_U8 ( .A1(stateFF_state_gff_12_n58), .A2(
        stateFF_state_gff_12_n57), .ZN(stateFF_state_gff_12_n32) );
  NAND2_X1 stateFF_state_gff_12_U7 ( .A1(stateFF_state_gff_12_n67), .A2(
        stateFF_permOut[11]), .ZN(stateFF_state_gff_12_n57) );
  NOR2_X1 stateFF_state_gff_12_U6 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_12_n56), .ZN(stateFF_state_gff_12_n67) );
  MUX2_X1 stateFF_state_gff_12_U5 ( .A(stateFF_state_gff_12_n36), .B(
        stateFF_state_gff_12_n55), .S(stateFF_state_gff_12_n65), .Z(
        stateFF_state_gff_12_n58) );
  INV_X1 stateFF_state_gff_12_U4 ( .A(stateFF_state_gff_12_n56), .ZN(
        stateFF_state_gff_12_n65) );
  INV_X1 stateFF_state_gff_12_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_12_n56) );
  NAND2_X1 stateFF_state_gff_12_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[44]), .ZN(stateFF_state_gff_12_n55) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_12_n32), .CK(clk), .Q(stateFF_permOut[12]), .QN(
        stateFF_state_gff_12_n36) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_12_n31), .CK(clk), .Q(stateFF_permOut[28]), .QN(
        stateFF_state_gff_12_n35) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_12_n30), .CK(clk), .Q(stateFF_permOut[44]), .QN(
        stateFF_state_gff_12_n34) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_12_n29), .CK(clk), .Q(stateFF_permOut[60]), .QN(
        stateFF_state_gff_12_n33) );
  NAND2_X1 stateFF_state_gff_13_U20 ( .A1(stateFF_state_gff_13_n69), .A2(
        stateFF_state_gff_13_n68), .ZN(stateFF_state_gff_13_n29) );
  NAND2_X1 stateFF_state_gff_13_U19 ( .A1(stateFF_state_gff_13_n67), .A2(
        stateFF_permOut[60]), .ZN(stateFF_state_gff_13_n68) );
  MUX2_X1 stateFF_state_gff_13_U18 ( .A(stateFF_state_gff_13_n33), .B(
        stateFF_state_gff_13_n66), .S(stateFF_state_gff_13_n65), .Z(
        stateFF_state_gff_13_n69) );
  NAND2_X1 stateFF_state_gff_13_U17 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[51]), .ZN(stateFF_state_gff_13_n66) );
  NAND2_X1 stateFF_state_gff_13_U16 ( .A1(stateFF_state_gff_13_n64), .A2(
        stateFF_state_gff_13_n63), .ZN(stateFF_state_gff_13_n30) );
  NAND2_X1 stateFF_state_gff_13_U15 ( .A1(stateFF_state_gff_13_n67), .A2(
        stateFF_permOut[44]), .ZN(stateFF_state_gff_13_n63) );
  MUX2_X1 stateFF_state_gff_13_U14 ( .A(stateFF_state_gff_13_n34), .B(
        stateFF_state_gff_13_n62), .S(stateFF_state_gff_13_n65), .Z(
        stateFF_state_gff_13_n64) );
  NAND2_X1 stateFF_state_gff_13_U13 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[50]), .ZN(stateFF_state_gff_13_n62) );
  NAND2_X1 stateFF_state_gff_13_U12 ( .A1(stateFF_state_gff_13_n61), .A2(
        stateFF_state_gff_13_n60), .ZN(stateFF_state_gff_13_n31) );
  NAND2_X1 stateFF_state_gff_13_U11 ( .A1(stateFF_state_gff_13_n67), .A2(
        stateFF_permOut[28]), .ZN(stateFF_state_gff_13_n60) );
  MUX2_X1 stateFF_state_gff_13_U10 ( .A(stateFF_state_gff_13_n35), .B(
        stateFF_state_gff_13_n59), .S(stateFF_state_gff_13_n65), .Z(
        stateFF_state_gff_13_n61) );
  NAND2_X1 stateFF_state_gff_13_U9 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[49]), .ZN(stateFF_state_gff_13_n59) );
  NAND2_X1 stateFF_state_gff_13_U8 ( .A1(stateFF_state_gff_13_n58), .A2(
        stateFF_state_gff_13_n57), .ZN(stateFF_state_gff_13_n32) );
  NAND2_X1 stateFF_state_gff_13_U7 ( .A1(stateFF_state_gff_13_n67), .A2(
        stateFF_permOut[12]), .ZN(stateFF_state_gff_13_n57) );
  NOR2_X1 stateFF_state_gff_13_U6 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_13_n56), .ZN(stateFF_state_gff_13_n67) );
  MUX2_X1 stateFF_state_gff_13_U5 ( .A(stateFF_state_gff_13_n36), .B(
        stateFF_state_gff_13_n55), .S(stateFF_state_gff_13_n65), .Z(
        stateFF_state_gff_13_n58) );
  INV_X1 stateFF_state_gff_13_U4 ( .A(stateFF_state_gff_13_n56), .ZN(
        stateFF_state_gff_13_n65) );
  INV_X1 stateFF_state_gff_13_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_13_n56) );
  NAND2_X1 stateFF_state_gff_13_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[48]), .ZN(stateFF_state_gff_13_n55) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_13_n32), .CK(clk), .Q(stateFF_permOut[13]), .QN(
        stateFF_state_gff_13_n36) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_13_n31), .CK(clk), .Q(stateFF_permOut[29]), .QN(
        stateFF_state_gff_13_n35) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_13_n30), .CK(clk), .Q(stateFF_permOut[45]), .QN(
        stateFF_state_gff_13_n34) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_13_n29), .CK(clk), .Q(stateFF_permOut[61]), .QN(
        stateFF_state_gff_13_n33) );
  NAND2_X1 stateFF_state_gff_14_U20 ( .A1(stateFF_state_gff_14_n69), .A2(
        stateFF_state_gff_14_n68), .ZN(stateFF_state_gff_14_n29) );
  NAND2_X1 stateFF_state_gff_14_U19 ( .A1(stateFF_state_gff_14_n67), .A2(
        stateFF_permOut[61]), .ZN(stateFF_state_gff_14_n68) );
  MUX2_X1 stateFF_state_gff_14_U18 ( .A(stateFF_state_gff_14_n33), .B(
        stateFF_state_gff_14_n66), .S(stateFF_state_gff_14_n65), .Z(
        stateFF_state_gff_14_n69) );
  NAND2_X1 stateFF_state_gff_14_U17 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[55]), .ZN(stateFF_state_gff_14_n66) );
  NAND2_X1 stateFF_state_gff_14_U16 ( .A1(stateFF_state_gff_14_n64), .A2(
        stateFF_state_gff_14_n63), .ZN(stateFF_state_gff_14_n30) );
  NAND2_X1 stateFF_state_gff_14_U15 ( .A1(stateFF_state_gff_14_n67), .A2(
        stateFF_permOut[45]), .ZN(stateFF_state_gff_14_n63) );
  MUX2_X1 stateFF_state_gff_14_U14 ( .A(stateFF_state_gff_14_n34), .B(
        stateFF_state_gff_14_n62), .S(stateFF_state_gff_14_n65), .Z(
        stateFF_state_gff_14_n64) );
  NAND2_X1 stateFF_state_gff_14_U13 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[54]), .ZN(stateFF_state_gff_14_n62) );
  NAND2_X1 stateFF_state_gff_14_U12 ( .A1(stateFF_state_gff_14_n61), .A2(
        stateFF_state_gff_14_n60), .ZN(stateFF_state_gff_14_n31) );
  NAND2_X1 stateFF_state_gff_14_U11 ( .A1(stateFF_state_gff_14_n67), .A2(
        stateFF_permOut[29]), .ZN(stateFF_state_gff_14_n60) );
  MUX2_X1 stateFF_state_gff_14_U10 ( .A(stateFF_state_gff_14_n35), .B(
        stateFF_state_gff_14_n59), .S(stateFF_state_gff_14_n65), .Z(
        stateFF_state_gff_14_n61) );
  NAND2_X1 stateFF_state_gff_14_U9 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[53]), .ZN(stateFF_state_gff_14_n59) );
  NAND2_X1 stateFF_state_gff_14_U8 ( .A1(stateFF_state_gff_14_n58), .A2(
        stateFF_state_gff_14_n57), .ZN(stateFF_state_gff_14_n32) );
  NAND2_X1 stateFF_state_gff_14_U7 ( .A1(stateFF_state_gff_14_n67), .A2(
        stateFF_permOut[13]), .ZN(stateFF_state_gff_14_n57) );
  NOR2_X1 stateFF_state_gff_14_U6 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_14_n56), .ZN(stateFF_state_gff_14_n67) );
  MUX2_X1 stateFF_state_gff_14_U5 ( .A(stateFF_state_gff_14_n36), .B(
        stateFF_state_gff_14_n55), .S(stateFF_state_gff_14_n65), .Z(
        stateFF_state_gff_14_n58) );
  INV_X1 stateFF_state_gff_14_U4 ( .A(stateFF_state_gff_14_n56), .ZN(
        stateFF_state_gff_14_n65) );
  INV_X1 stateFF_state_gff_14_U3 ( .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_14_n56) );
  NAND2_X1 stateFF_state_gff_14_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[52]), .ZN(stateFF_state_gff_14_n55) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_14_n32), .CK(clk), .Q(stateFF_permOut[14]), .QN(
        stateFF_state_gff_14_n36) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_14_n31), .CK(clk), .Q(stateFF_permOut[30]), .QN(
        stateFF_state_gff_14_n35) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_14_n30), .CK(clk), .Q(stateFF_permOut[46]), .QN(
        stateFF_state_gff_14_n34) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_14_n29), .CK(clk), .Q(stateFF_permOut[62]), .QN(
        stateFF_state_gff_14_n33) );
  NAND2_X1 stateFF_state_gff_15_U20 ( .A1(stateFF_state_gff_15_n69), .A2(
        stateFF_state_gff_15_n68), .ZN(stateFF_state_gff_15_n29) );
  NAND2_X1 stateFF_state_gff_15_U19 ( .A1(stateFF_state_gff_15_n67), .A2(
        stateFF_permOut[62]), .ZN(stateFF_state_gff_15_n68) );
  MUX2_X1 stateFF_state_gff_15_U18 ( .A(stateFF_state_gff_15_n33), .B(
        stateFF_state_gff_15_n66), .S(stateFF_state_gff_15_n65), .Z(
        stateFF_state_gff_15_n69) );
  NAND2_X1 stateFF_state_gff_15_U17 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[59]), .ZN(stateFF_state_gff_15_n66) );
  NAND2_X1 stateFF_state_gff_15_U16 ( .A1(stateFF_state_gff_15_n64), .A2(
        stateFF_state_gff_15_n63), .ZN(stateFF_state_gff_15_n30) );
  NAND2_X1 stateFF_state_gff_15_U15 ( .A1(stateFF_state_gff_15_n67), .A2(
        stateFF_permOut[46]), .ZN(stateFF_state_gff_15_n63) );
  MUX2_X1 stateFF_state_gff_15_U14 ( .A(stateFF_state_gff_15_n34), .B(
        stateFF_state_gff_15_n62), .S(stateFF_state_gff_15_n65), .Z(
        stateFF_state_gff_15_n64) );
  NAND2_X1 stateFF_state_gff_15_U13 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[58]), .ZN(stateFF_state_gff_15_n62) );
  NAND2_X1 stateFF_state_gff_15_U12 ( .A1(stateFF_state_gff_15_n61), .A2(
        stateFF_state_gff_15_n60), .ZN(stateFF_state_gff_15_n31) );
  NAND2_X1 stateFF_state_gff_15_U11 ( .A1(stateFF_state_gff_15_n67), .A2(
        stateFF_permOut[30]), .ZN(stateFF_state_gff_15_n60) );
  MUX2_X1 stateFF_state_gff_15_U10 ( .A(stateFF_state_gff_15_n35), .B(
        stateFF_state_gff_15_n59), .S(stateFF_state_gff_15_n65), .Z(
        stateFF_state_gff_15_n61) );
  NAND2_X1 stateFF_state_gff_15_U9 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[57]), .ZN(stateFF_state_gff_15_n59) );
  NAND2_X1 stateFF_state_gff_15_U8 ( .A1(stateFF_state_gff_15_n58), .A2(
        stateFF_state_gff_15_n57), .ZN(stateFF_state_gff_15_n32) );
  NAND2_X1 stateFF_state_gff_15_U7 ( .A1(stateFF_state_gff_15_n67), .A2(
        stateFF_permOut[14]), .ZN(stateFF_state_gff_15_n57) );
  NOR2_X1 stateFF_state_gff_15_U6 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_15_n56), .ZN(stateFF_state_gff_15_n67) );
  MUX2_X1 stateFF_state_gff_15_U5 ( .A(stateFF_state_gff_15_n36), .B(
        stateFF_state_gff_15_n55), .S(stateFF_state_gff_15_n65), .Z(
        stateFF_state_gff_15_n58) );
  INV_X1 stateFF_state_gff_15_U4 ( .A(stateFF_state_gff_15_n56), .ZN(
        stateFF_state_gff_15_n65) );
  INV_X1 stateFF_state_gff_15_U3 ( .A(ctrlData[1]), .ZN(
        stateFF_state_gff_15_n56) );
  NAND2_X1 stateFF_state_gff_15_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[56]), .ZN(stateFF_state_gff_15_n55) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_15_n32), .CK(clk), .Q(stateFF_permOut[15]), .QN(
        stateFF_state_gff_15_n36) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_15_n31), .CK(clk), .Q(stateFF_permOut[31]), .QN(
        stateFF_state_gff_15_n35) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_15_n30), .CK(clk), .Q(stateFF_permOut[47]), .QN(
        stateFF_state_gff_15_n34) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_15_n29), .CK(clk), .Q(stateFF_permOut[63]), .QN(
        stateFF_state_gff_15_n33) );
  NAND2_X1 stateFF_state_gff_16_U20 ( .A1(stateFF_state_gff_16_n68), .A2(
        stateFF_state_gff_16_n67), .ZN(stateFF_state_gff_16_n28) );
  NAND2_X1 stateFF_state_gff_16_U19 ( .A1(stateFF_state_gff_16_n66), .A2(
        stateFF_permOut[63]), .ZN(stateFF_state_gff_16_n67) );
  MUX2_X1 stateFF_state_gff_16_U18 ( .A(stateFF_state_gff_16_n32), .B(
        stateFF_state_gff_16_n65), .S(stateFF_state_gff_16_n64), .Z(
        stateFF_state_gff_16_n68) );
  NAND2_X1 stateFF_state_gff_16_U17 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[63]), .ZN(stateFF_state_gff_16_n65) );
  NAND2_X1 stateFF_state_gff_16_U16 ( .A1(stateFF_state_gff_16_n63), .A2(
        stateFF_state_gff_16_n62), .ZN(stateFF_state_gff_16_n29) );
  NAND2_X1 stateFF_state_gff_16_U15 ( .A1(stateFF_state_gff_16_n66), .A2(
        stateFF_permOut[47]), .ZN(stateFF_state_gff_16_n62) );
  MUX2_X1 stateFF_state_gff_16_U14 ( .A(stateFF_state_gff_16_n33), .B(
        stateFF_state_gff_16_n61), .S(stateFF_state_gff_16_n64), .Z(
        stateFF_state_gff_16_n63) );
  NAND2_X1 stateFF_state_gff_16_U13 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[62]), .ZN(stateFF_state_gff_16_n61) );
  NAND2_X1 stateFF_state_gff_16_U12 ( .A1(stateFF_state_gff_16_n60), .A2(
        stateFF_state_gff_16_n59), .ZN(stateFF_state_gff_16_n30) );
  NAND2_X1 stateFF_state_gff_16_U11 ( .A1(stateFF_state_gff_16_n66), .A2(
        stateFF_permOut[31]), .ZN(stateFF_state_gff_16_n59) );
  MUX2_X1 stateFF_state_gff_16_U10 ( .A(stateFF_state_gff_16_n34), .B(
        stateFF_state_gff_16_n58), .S(stateFF_state_gff_16_n64), .Z(
        stateFF_state_gff_16_n60) );
  NAND2_X1 stateFF_state_gff_16_U9 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[61]), .ZN(stateFF_state_gff_16_n58) );
  NAND2_X1 stateFF_state_gff_16_U8 ( .A1(stateFF_state_gff_16_n57), .A2(
        stateFF_state_gff_16_n56), .ZN(stateFF_state_gff_16_n31) );
  NAND2_X1 stateFF_state_gff_16_U7 ( .A1(stateFF_state_gff_16_n66), .A2(
        stateFF_permOut[15]), .ZN(stateFF_state_gff_16_n56) );
  NOR2_X1 stateFF_state_gff_16_U6 ( .A1(stateFF_state_n9), .A2(
        stateFF_state_gff_16_n55), .ZN(stateFF_state_gff_16_n66) );
  MUX2_X1 stateFF_state_gff_16_U5 ( .A(stateFF_state_gff_16_n35), .B(
        stateFF_state_gff_16_n54), .S(stateFF_state_gff_16_n64), .Z(
        stateFF_state_gff_16_n57) );
  INV_X1 stateFF_state_gff_16_U4 ( .A(stateFF_state_gff_16_n55), .ZN(
        stateFF_state_gff_16_n64) );
  INV_X1 stateFF_state_gff_16_U3 ( .A(ctrlData[1]), .ZN(
        stateFF_state_gff_16_n55) );
  NAND2_X1 stateFF_state_gff_16_U2 ( .A1(stateFF_state_n9), .A2(
        stateFF_inputPar[60]), .ZN(stateFF_state_gff_16_n54) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_0_ ( .D(
        stateFF_state_gff_16_n31), .CK(clk), .Q(state[0]), .QN(
        stateFF_state_gff_16_n35) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_1_ ( .D(
        stateFF_state_gff_16_n30), .CK(clk), .Q(state[1]), .QN(
        stateFF_state_gff_16_n34) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_2_ ( .D(
        stateFF_state_gff_16_n29), .CK(clk), .Q(state[2]), .QN(
        stateFF_state_gff_16_n33) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_3_ ( .D(
        stateFF_state_gff_16_n28), .CK(clk), .Q(state[3]), .QN(
        stateFF_state_gff_16_n32) );
  MUX2_X1 md1FF_U70 ( .A(md1FF_permOut[9]), .B(data_in2[9]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[9]) );
  MUX2_X1 md1FF_U69 ( .A(md1FF_permOut[8]), .B(data_in2[8]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[8]) );
  MUX2_X1 md1FF_U68 ( .A(md1FF_permOut[7]), .B(data_in2[7]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[7]) );
  MUX2_X1 md1FF_U67 ( .A(md1FF_permOut[6]), .B(data_in2[6]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[6]) );
  MUX2_X1 md1FF_U66 ( .A(md1FF_permOut[5]), .B(data_in2[5]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[5]) );
  MUX2_X1 md1FF_U65 ( .A(md1FF_permOut[4]), .B(data_in2[4]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[4]) );
  MUX2_X1 md1FF_U64 ( .A(md1FF_permOut[63]), .B(data_in2[63]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[63]) );
  MUX2_X1 md1FF_U63 ( .A(md1FF_permOut[62]), .B(data_in2[62]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[62]) );
  MUX2_X1 md1FF_U62 ( .A(md1FF_permOut[61]), .B(data_in2[61]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[61]) );
  MUX2_X1 md1FF_U61 ( .A(md1FF_permOut[60]), .B(data_in2[60]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[60]) );
  MUX2_X1 md1FF_U60 ( .A(md1FF_permOut[59]), .B(data_in2[59]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[59]) );
  MUX2_X1 md1FF_U59 ( .A(md1FF_permOut[58]), .B(data_in2[58]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[58]) );
  MUX2_X1 md1FF_U58 ( .A(md1FF_permOut[57]), .B(data_in2[57]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[57]) );
  MUX2_X1 md1FF_U57 ( .A(md1FF_permOut[56]), .B(data_in2[56]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[56]) );
  MUX2_X1 md1FF_U56 ( .A(md1FF_permOut[55]), .B(data_in2[55]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[55]) );
  MUX2_X1 md1FF_U55 ( .A(md1FF_permOut[54]), .B(data_in2[54]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[54]) );
  MUX2_X1 md1FF_U54 ( .A(md1FF_permOut[53]), .B(data_in2[53]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[53]) );
  MUX2_X1 md1FF_U53 ( .A(md1FF_permOut[52]), .B(data_in2[52]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[52]) );
  MUX2_X1 md1FF_U52 ( .A(md1FF_permOut[51]), .B(data_in2[51]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[51]) );
  MUX2_X1 md1FF_U51 ( .A(md1FF_permOut[50]), .B(data_in2[50]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[50]) );
  MUX2_X1 md1FF_U50 ( .A(md1FF_permOut[49]), .B(data_in2[49]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[49]) );
  MUX2_X1 md1FF_U49 ( .A(md1FF_permOut[48]), .B(data_in2[48]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[48]) );
  MUX2_X1 md1FF_U48 ( .A(md1FF_permOut[47]), .B(data_in2[47]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[47]) );
  MUX2_X1 md1FF_U47 ( .A(md1FF_permOut[46]), .B(data_in2[46]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[46]) );
  MUX2_X1 md1FF_U46 ( .A(md1FF_permOut[45]), .B(data_in2[45]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[45]) );
  MUX2_X1 md1FF_U45 ( .A(md1FF_permOut[44]), .B(data_in2[44]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[44]) );
  MUX2_X1 md1FF_U44 ( .A(md1FF_permOut[43]), .B(data_in2[43]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[43]) );
  MUX2_X1 md1FF_U43 ( .A(md1FF_permOut[42]), .B(data_in2[42]), .S(md1FF_n265), 
        .Z(md1FF_inputPar[42]) );
  INV_X1 md1FF_U42 ( .A(md1FF_n263), .ZN(md1FF_n265) );
  MUX2_X1 md1FF_U41 ( .A(md1FF_permOut[41]), .B(data_in2[41]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[41]) );
  MUX2_X1 md1FF_U40 ( .A(md1FF_permOut[40]), .B(data_in2[40]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[40]) );
  MUX2_X1 md1FF_U39 ( .A(md1FF_permOut[39]), .B(data_in2[39]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[39]) );
  MUX2_X1 md1FF_U38 ( .A(md1FF_permOut[38]), .B(data_in2[38]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[38]) );
  MUX2_X1 md1FF_U37 ( .A(md1FF_permOut[37]), .B(data_in2[37]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[37]) );
  MUX2_X1 md1FF_U36 ( .A(md1FF_permOut[36]), .B(data_in2[36]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[36]) );
  MUX2_X1 md1FF_U35 ( .A(md1FF_permOut[35]), .B(data_in2[35]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[35]) );
  MUX2_X1 md1FF_U34 ( .A(md1FF_permOut[34]), .B(data_in2[34]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[34]) );
  MUX2_X1 md1FF_U33 ( .A(md1FF_permOut[33]), .B(data_in2[33]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[33]) );
  MUX2_X1 md1FF_U32 ( .A(md1FF_permOut[32]), .B(data_in2[32]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[32]) );
  MUX2_X1 md1FF_U31 ( .A(md1FF_permOut[31]), .B(data_in2[31]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[31]) );
  MUX2_X1 md1FF_U30 ( .A(md1FF_permOut[30]), .B(data_in2[30]), .S(md1FF_n266), 
        .Z(md1FF_inputPar[30]) );
  INV_X1 md1FF_U29 ( .A(md1FF_n263), .ZN(md1FF_n266) );
  MUX2_X1 md1FF_U28 ( .A(md1FF_permOut[29]), .B(data_in2[29]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[29]) );
  MUX2_X1 md1FF_U27 ( .A(md1FF_permOut[28]), .B(data_in2[28]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[28]) );
  MUX2_X1 md1FF_U26 ( .A(md1FF_permOut[27]), .B(data_in2[27]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[27]) );
  MUX2_X1 md1FF_U25 ( .A(md1FF_permOut[26]), .B(data_in2[26]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[26]) );
  MUX2_X1 md1FF_U24 ( .A(md1FF_permOut[25]), .B(data_in2[25]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[25]) );
  MUX2_X1 md1FF_U23 ( .A(md1FF_permOut[24]), .B(data_in2[24]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[24]) );
  MUX2_X1 md1FF_U22 ( .A(md1FF_permOut[23]), .B(data_in2[23]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[23]) );
  MUX2_X1 md1FF_U21 ( .A(md1FF_permOut[22]), .B(data_in2[22]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[22]) );
  MUX2_X1 md1FF_U20 ( .A(md1FF_permOut[21]), .B(data_in2[21]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[21]) );
  MUX2_X1 md1FF_U19 ( .A(md1FF_permOut[20]), .B(data_in2[20]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[20]) );
  MUX2_X1 md1FF_U18 ( .A(md1FF_permOut[19]), .B(data_in2[19]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[19]) );
  MUX2_X1 md1FF_U17 ( .A(md1FF_permOut[18]), .B(data_in2[18]), .S(md1FF_n267), 
        .Z(md1FF_inputPar[18]) );
  INV_X1 md1FF_U16 ( .A(md1FF_n263), .ZN(md1FF_n267) );
  MUX2_X1 md1FF_U15 ( .A(md1FF_permOut[17]), .B(data_in2[17]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[17]) );
  MUX2_X1 md1FF_U14 ( .A(md1FF_permOut[16]), .B(data_in2[16]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[16]) );
  MUX2_X1 md1FF_U13 ( .A(md1FF_permOut[15]), .B(data_in2[15]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[15]) );
  MUX2_X1 md1FF_U12 ( .A(md1FF_permOut[14]), .B(data_in2[14]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[14]) );
  MUX2_X1 md1FF_U11 ( .A(md1FF_permOut[13]), .B(data_in2[13]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[13]) );
  MUX2_X1 md1FF_U10 ( .A(md1FF_permOut[12]), .B(data_in2[12]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[12]) );
  MUX2_X1 md1FF_U9 ( .A(md1FF_permOut[11]), .B(data_in2[11]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[11]) );
  MUX2_X1 md1FF_U8 ( .A(md1FF_permOut[10]), .B(data_in2[10]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[10]) );
  MUX2_X1 md1FF_U7 ( .A(md1FF_permOut[3]), .B(data_in2[3]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[3]) );
  MUX2_X1 md1FF_U6 ( .A(md1FF_permOut[2]), .B(data_in2[2]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[2]) );
  MUX2_X1 md1FF_U5 ( .A(md1FF_permOut[1]), .B(data_in2[1]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[1]) );
  MUX2_X1 md1FF_U4 ( .A(md1FF_permOut[0]), .B(data_in2[0]), .S(md1FF_n264), 
        .Z(md1FF_inputPar[0]) );
  INV_X1 md1FF_U3 ( .A(md1FF_n263), .ZN(md1FF_n264) );
  INV_X1 md1FF_U2 ( .A(ctrlData[2]), .ZN(md1FF_n263) );
  INV_X2 md1FF_state_U5 ( .A(md1FF_state_n11), .ZN(md1FF_state_n10) );
  INV_X2 md1FF_state_U4 ( .A(md1FF_state_n11), .ZN(md1FF_state_n9) );
  INV_X1 md1FF_state_U3 ( .A(ctrlData[0]), .ZN(md1FF_state_n11) );
  INV_X1 md1FF_state_U2 ( .A(ctrlData[1]), .ZN(md1FF_state_n8) );
  INV_X1 md1FF_state_U1 ( .A(md1FF_state_n8), .ZN(md1FF_state_n7) );
  NAND2_X1 md1FF_state_gff_1_U19 ( .A1(md1FF_state_gff_1_n67), .A2(
        md1FF_state_gff_1_n66), .ZN(md1FF_state_gff_1_n28) );
  NAND2_X1 md1FF_state_gff_1_U18 ( .A1(md1FF_state_gff_1_n65), .A2(
        md1FF_permOut[48]), .ZN(md1FF_state_gff_1_n66) );
  MUX2_X1 md1FF_state_gff_1_U17 ( .A(md1FF_state_gff_1_n32), .B(
        md1FF_state_gff_1_n64), .S(md1FF_state_n7), .Z(md1FF_state_gff_1_n67)
         );
  NAND2_X1 md1FF_state_gff_1_U16 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[3]), 
        .ZN(md1FF_state_gff_1_n64) );
  NAND2_X1 md1FF_state_gff_1_U15 ( .A1(md1FF_state_gff_1_n63), .A2(
        md1FF_state_gff_1_n62), .ZN(md1FF_state_gff_1_n30) );
  NAND2_X1 md1FF_state_gff_1_U14 ( .A1(md1FF_state_gff_1_n65), .A2(
        md1FF_permOut[16]), .ZN(md1FF_state_gff_1_n62) );
  MUX2_X1 md1FF_state_gff_1_U13 ( .A(md1FF_state_gff_1_n34), .B(
        md1FF_state_gff_1_n61), .S(md1FF_state_n7), .Z(md1FF_state_gff_1_n63)
         );
  NAND2_X1 md1FF_state_gff_1_U12 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[1]), 
        .ZN(md1FF_state_gff_1_n61) );
  NAND2_X1 md1FF_state_gff_1_U11 ( .A1(md1FF_state_gff_1_n60), .A2(
        md1FF_state_gff_1_n59), .ZN(md1FF_state_gff_1_n31) );
  NAND2_X1 md1FF_state_gff_1_U10 ( .A1(md1FF_state_gff_1_n65), .A2(
        md1FF_permOut[0]), .ZN(md1FF_state_gff_1_n59) );
  MUX2_X1 md1FF_state_gff_1_U9 ( .A(md1FF_state_gff_1_n35), .B(
        md1FF_state_gff_1_n58), .S(md1FF_state_n7), .Z(md1FF_state_gff_1_n60)
         );
  NAND2_X1 md1FF_state_gff_1_U8 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[0]), 
        .ZN(md1FF_state_gff_1_n58) );
  NAND2_X1 md1FF_state_gff_1_U7 ( .A1(md1FF_state_gff_1_n57), .A2(
        md1FF_state_gff_1_n56), .ZN(md1FF_state_gff_1_n29) );
  NAND2_X1 md1FF_state_gff_1_U6 ( .A1(md1FF_state_gff_1_n65), .A2(
        md1FF_permOut[32]), .ZN(md1FF_state_gff_1_n56) );
  NOR2_X1 md1FF_state_gff_1_U5 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_1_n55), .ZN(md1FF_state_gff_1_n65) );
  INV_X1 md1FF_state_gff_1_U4 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_1_n55)
         );
  MUX2_X1 md1FF_state_gff_1_U3 ( .A(md1FF_state_gff_1_n33), .B(
        md1FF_state_gff_1_n54), .S(md1FF_state_n7), .Z(md1FF_state_gff_1_n57)
         );
  NAND2_X1 md1FF_state_gff_1_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[2]), 
        .ZN(md1FF_state_gff_1_n54) );
  DFF_X1 md1FF_state_gff_1_s_current_state_reg_0_ ( .D(md1FF_state_gff_1_n31), 
        .CK(clk), .Q(md1FF_permOut[1]), .QN(md1FF_state_gff_1_n35) );
  DFF_X1 md1FF_state_gff_1_s_current_state_reg_1_ ( .D(md1FF_state_gff_1_n30), 
        .CK(clk), .Q(md1FF_permOut[17]), .QN(md1FF_state_gff_1_n34) );
  DFF_X1 md1FF_state_gff_1_s_current_state_reg_2_ ( .D(md1FF_state_gff_1_n29), 
        .CK(clk), .Q(md1FF_permOut[33]), .QN(md1FF_state_gff_1_n33) );
  DFF_X1 md1FF_state_gff_1_s_current_state_reg_3_ ( .D(md1FF_state_gff_1_n28), 
        .CK(clk), .Q(md1FF_permOut[49]), .QN(md1FF_state_gff_1_n32) );
  NAND2_X1 md1FF_state_gff_2_U20 ( .A1(md1FF_state_gff_2_n68), .A2(
        md1FF_state_gff_2_n67), .ZN(md1FF_state_gff_2_n28) );
  NAND2_X1 md1FF_state_gff_2_U19 ( .A1(md1FF_state_gff_2_n66), .A2(
        md1FF_permOut[49]), .ZN(md1FF_state_gff_2_n67) );
  MUX2_X1 md1FF_state_gff_2_U18 ( .A(md1FF_state_gff_2_n32), .B(
        md1FF_state_gff_2_n65), .S(md1FF_state_gff_2_n64), .Z(
        md1FF_state_gff_2_n68) );
  NAND2_X1 md1FF_state_gff_2_U17 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[7]), 
        .ZN(md1FF_state_gff_2_n65) );
  NAND2_X1 md1FF_state_gff_2_U16 ( .A1(md1FF_state_gff_2_n63), .A2(
        md1FF_state_gff_2_n62), .ZN(md1FF_state_gff_2_n29) );
  NAND2_X1 md1FF_state_gff_2_U15 ( .A1(md1FF_state_gff_2_n66), .A2(
        md1FF_permOut[33]), .ZN(md1FF_state_gff_2_n62) );
  MUX2_X1 md1FF_state_gff_2_U14 ( .A(md1FF_state_gff_2_n33), .B(
        md1FF_state_gff_2_n61), .S(md1FF_state_gff_2_n64), .Z(
        md1FF_state_gff_2_n63) );
  NAND2_X1 md1FF_state_gff_2_U13 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[6]), 
        .ZN(md1FF_state_gff_2_n61) );
  NAND2_X1 md1FF_state_gff_2_U12 ( .A1(md1FF_state_gff_2_n60), .A2(
        md1FF_state_gff_2_n59), .ZN(md1FF_state_gff_2_n30) );
  NAND2_X1 md1FF_state_gff_2_U11 ( .A1(md1FF_state_gff_2_n66), .A2(
        md1FF_permOut[17]), .ZN(md1FF_state_gff_2_n59) );
  MUX2_X1 md1FF_state_gff_2_U10 ( .A(md1FF_state_gff_2_n34), .B(
        md1FF_state_gff_2_n58), .S(md1FF_state_gff_2_n64), .Z(
        md1FF_state_gff_2_n60) );
  NAND2_X1 md1FF_state_gff_2_U9 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[5]), 
        .ZN(md1FF_state_gff_2_n58) );
  NAND2_X1 md1FF_state_gff_2_U8 ( .A1(md1FF_state_gff_2_n57), .A2(
        md1FF_state_gff_2_n56), .ZN(md1FF_state_gff_2_n31) );
  NAND2_X1 md1FF_state_gff_2_U7 ( .A1(md1FF_state_gff_2_n66), .A2(
        md1FF_permOut[1]), .ZN(md1FF_state_gff_2_n56) );
  NOR2_X1 md1FF_state_gff_2_U6 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_2_n55), .ZN(md1FF_state_gff_2_n66) );
  MUX2_X1 md1FF_state_gff_2_U5 ( .A(md1FF_state_gff_2_n35), .B(
        md1FF_state_gff_2_n54), .S(md1FF_state_gff_2_n64), .Z(
        md1FF_state_gff_2_n57) );
  INV_X1 md1FF_state_gff_2_U4 ( .A(md1FF_state_gff_2_n55), .ZN(
        md1FF_state_gff_2_n64) );
  INV_X1 md1FF_state_gff_2_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_2_n55)
         );
  NAND2_X1 md1FF_state_gff_2_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[4]), 
        .ZN(md1FF_state_gff_2_n54) );
  DFF_X1 md1FF_state_gff_2_s_current_state_reg_0_ ( .D(md1FF_state_gff_2_n31), 
        .CK(clk), .Q(md1FF_permOut[2]), .QN(md1FF_state_gff_2_n35) );
  DFF_X1 md1FF_state_gff_2_s_current_state_reg_1_ ( .D(md1FF_state_gff_2_n30), 
        .CK(clk), .Q(md1FF_permOut[18]), .QN(md1FF_state_gff_2_n34) );
  DFF_X1 md1FF_state_gff_2_s_current_state_reg_2_ ( .D(md1FF_state_gff_2_n29), 
        .CK(clk), .Q(md1FF_permOut[34]), .QN(md1FF_state_gff_2_n33) );
  DFF_X1 md1FF_state_gff_2_s_current_state_reg_3_ ( .D(md1FF_state_gff_2_n28), 
        .CK(clk), .Q(md1FF_permOut[50]), .QN(md1FF_state_gff_2_n32) );
  NAND2_X1 md1FF_state_gff_3_U20 ( .A1(md1FF_state_gff_3_n68), .A2(
        md1FF_state_gff_3_n67), .ZN(md1FF_state_gff_3_n30) );
  NAND2_X1 md1FF_state_gff_3_U19 ( .A1(md1FF_state_gff_3_n66), .A2(
        md1FF_permOut[18]), .ZN(md1FF_state_gff_3_n67) );
  MUX2_X1 md1FF_state_gff_3_U18 ( .A(md1FF_state_gff_3_n34), .B(
        md1FF_state_gff_3_n65), .S(md1FF_state_gff_3_n64), .Z(
        md1FF_state_gff_3_n68) );
  NAND2_X1 md1FF_state_gff_3_U17 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[9]), .ZN(md1FF_state_gff_3_n65) );
  NAND2_X1 md1FF_state_gff_3_U16 ( .A1(md1FF_state_gff_3_n63), .A2(
        md1FF_state_gff_3_n62), .ZN(md1FF_state_gff_3_n31) );
  NAND2_X1 md1FF_state_gff_3_U15 ( .A1(md1FF_state_gff_3_n66), .A2(
        md1FF_permOut[2]), .ZN(md1FF_state_gff_3_n62) );
  MUX2_X1 md1FF_state_gff_3_U14 ( .A(md1FF_state_gff_3_n35), .B(
        md1FF_state_gff_3_n61), .S(md1FF_state_gff_3_n64), .Z(
        md1FF_state_gff_3_n63) );
  NAND2_X1 md1FF_state_gff_3_U13 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[8]), .ZN(md1FF_state_gff_3_n61) );
  NAND2_X1 md1FF_state_gff_3_U12 ( .A1(md1FF_state_gff_3_n60), .A2(
        md1FF_state_gff_3_n59), .ZN(md1FF_state_gff_3_n28) );
  NAND2_X1 md1FF_state_gff_3_U11 ( .A1(md1FF_state_gff_3_n66), .A2(
        md1FF_permOut[50]), .ZN(md1FF_state_gff_3_n59) );
  MUX2_X1 md1FF_state_gff_3_U10 ( .A(md1FF_state_gff_3_n32), .B(
        md1FF_state_gff_3_n58), .S(md1FF_state_gff_3_n64), .Z(
        md1FF_state_gff_3_n60) );
  NAND2_X1 md1FF_state_gff_3_U9 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[11]), .ZN(md1FF_state_gff_3_n58) );
  NAND2_X1 md1FF_state_gff_3_U8 ( .A1(md1FF_state_gff_3_n57), .A2(
        md1FF_state_gff_3_n56), .ZN(md1FF_state_gff_3_n29) );
  NAND2_X1 md1FF_state_gff_3_U7 ( .A1(md1FF_state_gff_3_n66), .A2(
        md1FF_permOut[34]), .ZN(md1FF_state_gff_3_n56) );
  NOR2_X1 md1FF_state_gff_3_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_3_n55), .ZN(md1FF_state_gff_3_n66) );
  MUX2_X1 md1FF_state_gff_3_U5 ( .A(md1FF_state_gff_3_n33), .B(
        md1FF_state_gff_3_n54), .S(md1FF_state_gff_3_n64), .Z(
        md1FF_state_gff_3_n57) );
  INV_X1 md1FF_state_gff_3_U4 ( .A(md1FF_state_gff_3_n55), .ZN(
        md1FF_state_gff_3_n64) );
  INV_X1 md1FF_state_gff_3_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_3_n55)
         );
  NAND2_X1 md1FF_state_gff_3_U2 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[10]), .ZN(md1FF_state_gff_3_n54) );
  DFF_X1 md1FF_state_gff_3_s_current_state_reg_0_ ( .D(md1FF_state_gff_3_n31), 
        .CK(clk), .Q(md1FF_permOut[3]), .QN(md1FF_state_gff_3_n35) );
  DFF_X1 md1FF_state_gff_3_s_current_state_reg_1_ ( .D(md1FF_state_gff_3_n30), 
        .CK(clk), .Q(md1FF_permOut[19]), .QN(md1FF_state_gff_3_n34) );
  DFF_X1 md1FF_state_gff_3_s_current_state_reg_2_ ( .D(md1FF_state_gff_3_n29), 
        .CK(clk), .Q(md1FF_permOut[35]), .QN(md1FF_state_gff_3_n33) );
  DFF_X1 md1FF_state_gff_3_s_current_state_reg_3_ ( .D(md1FF_state_gff_3_n28), 
        .CK(clk), .Q(md1FF_permOut[51]), .QN(md1FF_state_gff_3_n32) );
  NAND2_X1 md1FF_state_gff_4_U20 ( .A1(md1FF_state_gff_4_n68), .A2(
        md1FF_state_gff_4_n67), .ZN(md1FF_state_gff_4_n28) );
  NAND2_X1 md1FF_state_gff_4_U19 ( .A1(md1FF_state_gff_4_n66), .A2(
        md1FF_permOut[51]), .ZN(md1FF_state_gff_4_n67) );
  MUX2_X1 md1FF_state_gff_4_U18 ( .A(md1FF_state_gff_4_n32), .B(
        md1FF_state_gff_4_n65), .S(md1FF_state_gff_4_n64), .Z(
        md1FF_state_gff_4_n68) );
  NAND2_X1 md1FF_state_gff_4_U17 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[15]), .ZN(md1FF_state_gff_4_n65) );
  NAND2_X1 md1FF_state_gff_4_U16 ( .A1(md1FF_state_gff_4_n63), .A2(
        md1FF_state_gff_4_n62), .ZN(md1FF_state_gff_4_n29) );
  NAND2_X1 md1FF_state_gff_4_U15 ( .A1(md1FF_state_gff_4_n66), .A2(
        md1FF_permOut[35]), .ZN(md1FF_state_gff_4_n62) );
  MUX2_X1 md1FF_state_gff_4_U14 ( .A(md1FF_state_gff_4_n33), .B(
        md1FF_state_gff_4_n61), .S(md1FF_state_gff_4_n64), .Z(
        md1FF_state_gff_4_n63) );
  NAND2_X1 md1FF_state_gff_4_U13 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[14]), .ZN(md1FF_state_gff_4_n61) );
  NAND2_X1 md1FF_state_gff_4_U12 ( .A1(md1FF_state_gff_4_n60), .A2(
        md1FF_state_gff_4_n59), .ZN(md1FF_state_gff_4_n30) );
  NAND2_X1 md1FF_state_gff_4_U11 ( .A1(md1FF_state_gff_4_n66), .A2(
        md1FF_permOut[19]), .ZN(md1FF_state_gff_4_n59) );
  MUX2_X1 md1FF_state_gff_4_U10 ( .A(md1FF_state_gff_4_n34), .B(
        md1FF_state_gff_4_n58), .S(md1FF_state_gff_4_n64), .Z(
        md1FF_state_gff_4_n60) );
  NAND2_X1 md1FF_state_gff_4_U9 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[13]), .ZN(md1FF_state_gff_4_n58) );
  NAND2_X1 md1FF_state_gff_4_U8 ( .A1(md1FF_state_gff_4_n57), .A2(
        md1FF_state_gff_4_n56), .ZN(md1FF_state_gff_4_n31) );
  NAND2_X1 md1FF_state_gff_4_U7 ( .A1(md1FF_state_gff_4_n66), .A2(
        md1FF_permOut[3]), .ZN(md1FF_state_gff_4_n56) );
  NOR2_X1 md1FF_state_gff_4_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_4_n55), .ZN(md1FF_state_gff_4_n66) );
  MUX2_X1 md1FF_state_gff_4_U5 ( .A(md1FF_state_gff_4_n35), .B(
        md1FF_state_gff_4_n54), .S(md1FF_state_gff_4_n64), .Z(
        md1FF_state_gff_4_n57) );
  INV_X1 md1FF_state_gff_4_U4 ( .A(md1FF_state_gff_4_n55), .ZN(
        md1FF_state_gff_4_n64) );
  INV_X1 md1FF_state_gff_4_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_4_n55)
         );
  NAND2_X1 md1FF_state_gff_4_U2 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[12]), .ZN(md1FF_state_gff_4_n54) );
  DFF_X1 md1FF_state_gff_4_s_current_state_reg_0_ ( .D(md1FF_state_gff_4_n31), 
        .CK(clk), .Q(md1FF_permOut[4]), .QN(md1FF_state_gff_4_n35) );
  DFF_X1 md1FF_state_gff_4_s_current_state_reg_1_ ( .D(md1FF_state_gff_4_n30), 
        .CK(clk), .Q(md1FF_permOut[20]), .QN(md1FF_state_gff_4_n34) );
  DFF_X1 md1FF_state_gff_4_s_current_state_reg_2_ ( .D(md1FF_state_gff_4_n29), 
        .CK(clk), .Q(md1FF_permOut[36]), .QN(md1FF_state_gff_4_n33) );
  DFF_X1 md1FF_state_gff_4_s_current_state_reg_3_ ( .D(md1FF_state_gff_4_n28), 
        .CK(clk), .Q(md1FF_permOut[52]), .QN(md1FF_state_gff_4_n32) );
  NAND2_X1 md1FF_state_gff_5_U20 ( .A1(md1FF_state_gff_5_n69), .A2(
        md1FF_state_gff_5_n68), .ZN(md1FF_state_gff_5_n29) );
  NAND2_X1 md1FF_state_gff_5_U19 ( .A1(md1FF_state_gff_5_n67), .A2(
        md1FF_permOut[52]), .ZN(md1FF_state_gff_5_n68) );
  MUX2_X1 md1FF_state_gff_5_U18 ( .A(md1FF_state_gff_5_n33), .B(
        md1FF_state_gff_5_n66), .S(md1FF_state_gff_5_n65), .Z(
        md1FF_state_gff_5_n69) );
  NAND2_X1 md1FF_state_gff_5_U17 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[19]), .ZN(md1FF_state_gff_5_n66) );
  NAND2_X1 md1FF_state_gff_5_U16 ( .A1(md1FF_state_gff_5_n64), .A2(
        md1FF_state_gff_5_n63), .ZN(md1FF_state_gff_5_n30) );
  NAND2_X1 md1FF_state_gff_5_U15 ( .A1(md1FF_state_gff_5_n67), .A2(
        md1FF_permOut[36]), .ZN(md1FF_state_gff_5_n63) );
  MUX2_X1 md1FF_state_gff_5_U14 ( .A(md1FF_state_gff_5_n34), .B(
        md1FF_state_gff_5_n62), .S(md1FF_state_gff_5_n65), .Z(
        md1FF_state_gff_5_n64) );
  NAND2_X1 md1FF_state_gff_5_U13 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[18]), .ZN(md1FF_state_gff_5_n62) );
  NAND2_X1 md1FF_state_gff_5_U12 ( .A1(md1FF_state_gff_5_n61), .A2(
        md1FF_state_gff_5_n60), .ZN(md1FF_state_gff_5_n31) );
  NAND2_X1 md1FF_state_gff_5_U11 ( .A1(md1FF_state_gff_5_n67), .A2(
        md1FF_permOut[20]), .ZN(md1FF_state_gff_5_n60) );
  MUX2_X1 md1FF_state_gff_5_U10 ( .A(md1FF_state_gff_5_n35), .B(
        md1FF_state_gff_5_n59), .S(md1FF_state_gff_5_n65), .Z(
        md1FF_state_gff_5_n61) );
  NAND2_X1 md1FF_state_gff_5_U9 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[17]), .ZN(md1FF_state_gff_5_n59) );
  NAND2_X1 md1FF_state_gff_5_U8 ( .A1(md1FF_state_gff_5_n58), .A2(
        md1FF_state_gff_5_n57), .ZN(md1FF_state_gff_5_n32) );
  NAND2_X1 md1FF_state_gff_5_U7 ( .A1(md1FF_state_gff_5_n67), .A2(
        md1FF_permOut[4]), .ZN(md1FF_state_gff_5_n57) );
  NOR2_X1 md1FF_state_gff_5_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_5_n56), .ZN(md1FF_state_gff_5_n67) );
  MUX2_X1 md1FF_state_gff_5_U5 ( .A(md1FF_state_gff_5_n36), .B(
        md1FF_state_gff_5_n55), .S(md1FF_state_gff_5_n65), .Z(
        md1FF_state_gff_5_n58) );
  INV_X1 md1FF_state_gff_5_U4 ( .A(md1FF_state_gff_5_n56), .ZN(
        md1FF_state_gff_5_n65) );
  INV_X1 md1FF_state_gff_5_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_5_n56)
         );
  NAND2_X1 md1FF_state_gff_5_U2 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[16]), .ZN(md1FF_state_gff_5_n55) );
  DFF_X1 md1FF_state_gff_5_s_current_state_reg_0_ ( .D(md1FF_state_gff_5_n32), 
        .CK(clk), .Q(md1FF_permOut[5]), .QN(md1FF_state_gff_5_n36) );
  DFF_X1 md1FF_state_gff_5_s_current_state_reg_1_ ( .D(md1FF_state_gff_5_n31), 
        .CK(clk), .Q(md1FF_permOut[21]), .QN(md1FF_state_gff_5_n35) );
  DFF_X1 md1FF_state_gff_5_s_current_state_reg_2_ ( .D(md1FF_state_gff_5_n30), 
        .CK(clk), .Q(md1FF_permOut[37]), .QN(md1FF_state_gff_5_n34) );
  DFF_X1 md1FF_state_gff_5_s_current_state_reg_3_ ( .D(md1FF_state_gff_5_n29), 
        .CK(clk), .Q(md1FF_permOut[53]), .QN(md1FF_state_gff_5_n33) );
  NAND2_X1 md1FF_state_gff_6_U20 ( .A1(md1FF_state_gff_6_n69), .A2(
        md1FF_state_gff_6_n68), .ZN(md1FF_state_gff_6_n29) );
  NAND2_X1 md1FF_state_gff_6_U19 ( .A1(md1FF_state_gff_6_n67), .A2(
        md1FF_permOut[53]), .ZN(md1FF_state_gff_6_n68) );
  MUX2_X1 md1FF_state_gff_6_U18 ( .A(md1FF_state_gff_6_n33), .B(
        md1FF_state_gff_6_n66), .S(md1FF_state_gff_6_n65), .Z(
        md1FF_state_gff_6_n69) );
  NAND2_X1 md1FF_state_gff_6_U17 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[23]), .ZN(md1FF_state_gff_6_n66) );
  NAND2_X1 md1FF_state_gff_6_U16 ( .A1(md1FF_state_gff_6_n64), .A2(
        md1FF_state_gff_6_n63), .ZN(md1FF_state_gff_6_n30) );
  NAND2_X1 md1FF_state_gff_6_U15 ( .A1(md1FF_state_gff_6_n67), .A2(
        md1FF_permOut[37]), .ZN(md1FF_state_gff_6_n63) );
  MUX2_X1 md1FF_state_gff_6_U14 ( .A(md1FF_state_gff_6_n34), .B(
        md1FF_state_gff_6_n62), .S(md1FF_state_gff_6_n65), .Z(
        md1FF_state_gff_6_n64) );
  NAND2_X1 md1FF_state_gff_6_U13 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[22]), .ZN(md1FF_state_gff_6_n62) );
  NAND2_X1 md1FF_state_gff_6_U12 ( .A1(md1FF_state_gff_6_n61), .A2(
        md1FF_state_gff_6_n60), .ZN(md1FF_state_gff_6_n31) );
  NAND2_X1 md1FF_state_gff_6_U11 ( .A1(md1FF_state_gff_6_n67), .A2(
        md1FF_permOut[21]), .ZN(md1FF_state_gff_6_n60) );
  MUX2_X1 md1FF_state_gff_6_U10 ( .A(md1FF_state_gff_6_n35), .B(
        md1FF_state_gff_6_n59), .S(md1FF_state_gff_6_n65), .Z(
        md1FF_state_gff_6_n61) );
  NAND2_X1 md1FF_state_gff_6_U9 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[21]), .ZN(md1FF_state_gff_6_n59) );
  NAND2_X1 md1FF_state_gff_6_U8 ( .A1(md1FF_state_gff_6_n58), .A2(
        md1FF_state_gff_6_n57), .ZN(md1FF_state_gff_6_n32) );
  NAND2_X1 md1FF_state_gff_6_U7 ( .A1(md1FF_state_gff_6_n67), .A2(
        md1FF_permOut[5]), .ZN(md1FF_state_gff_6_n57) );
  NOR2_X1 md1FF_state_gff_6_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_6_n56), .ZN(md1FF_state_gff_6_n67) );
  MUX2_X1 md1FF_state_gff_6_U5 ( .A(md1FF_state_gff_6_n36), .B(
        md1FF_state_gff_6_n55), .S(md1FF_state_gff_6_n65), .Z(
        md1FF_state_gff_6_n58) );
  INV_X1 md1FF_state_gff_6_U4 ( .A(md1FF_state_gff_6_n56), .ZN(
        md1FF_state_gff_6_n65) );
  INV_X1 md1FF_state_gff_6_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_6_n56)
         );
  NAND2_X1 md1FF_state_gff_6_U2 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[20]), .ZN(md1FF_state_gff_6_n55) );
  DFF_X1 md1FF_state_gff_6_s_current_state_reg_0_ ( .D(md1FF_state_gff_6_n32), 
        .CK(clk), .Q(md1FF_permOut[6]), .QN(md1FF_state_gff_6_n36) );
  DFF_X1 md1FF_state_gff_6_s_current_state_reg_1_ ( .D(md1FF_state_gff_6_n31), 
        .CK(clk), .Q(md1FF_permOut[22]), .QN(md1FF_state_gff_6_n35) );
  DFF_X1 md1FF_state_gff_6_s_current_state_reg_2_ ( .D(md1FF_state_gff_6_n30), 
        .CK(clk), .Q(md1FF_permOut[38]), .QN(md1FF_state_gff_6_n34) );
  DFF_X1 md1FF_state_gff_6_s_current_state_reg_3_ ( .D(md1FF_state_gff_6_n29), 
        .CK(clk), .Q(md1FF_permOut[54]), .QN(md1FF_state_gff_6_n33) );
  NAND2_X1 md1FF_state_gff_7_U20 ( .A1(md1FF_state_gff_7_n69), .A2(
        md1FF_state_gff_7_n68), .ZN(md1FF_state_gff_7_n29) );
  NAND2_X1 md1FF_state_gff_7_U19 ( .A1(md1FF_state_gff_7_n67), .A2(
        md1FF_permOut[54]), .ZN(md1FF_state_gff_7_n68) );
  MUX2_X1 md1FF_state_gff_7_U18 ( .A(md1FF_state_gff_7_n33), .B(
        md1FF_state_gff_7_n66), .S(md1FF_state_gff_7_n65), .Z(
        md1FF_state_gff_7_n69) );
  NAND2_X1 md1FF_state_gff_7_U17 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[27]), .ZN(md1FF_state_gff_7_n66) );
  NAND2_X1 md1FF_state_gff_7_U16 ( .A1(md1FF_state_gff_7_n64), .A2(
        md1FF_state_gff_7_n63), .ZN(md1FF_state_gff_7_n30) );
  NAND2_X1 md1FF_state_gff_7_U15 ( .A1(md1FF_state_gff_7_n67), .A2(
        md1FF_permOut[38]), .ZN(md1FF_state_gff_7_n63) );
  MUX2_X1 md1FF_state_gff_7_U14 ( .A(md1FF_state_gff_7_n34), .B(
        md1FF_state_gff_7_n62), .S(md1FF_state_gff_7_n65), .Z(
        md1FF_state_gff_7_n64) );
  NAND2_X1 md1FF_state_gff_7_U13 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[26]), .ZN(md1FF_state_gff_7_n62) );
  NAND2_X1 md1FF_state_gff_7_U12 ( .A1(md1FF_state_gff_7_n61), .A2(
        md1FF_state_gff_7_n60), .ZN(md1FF_state_gff_7_n31) );
  NAND2_X1 md1FF_state_gff_7_U11 ( .A1(md1FF_state_gff_7_n67), .A2(
        md1FF_permOut[22]), .ZN(md1FF_state_gff_7_n60) );
  MUX2_X1 md1FF_state_gff_7_U10 ( .A(md1FF_state_gff_7_n35), .B(
        md1FF_state_gff_7_n59), .S(md1FF_state_gff_7_n65), .Z(
        md1FF_state_gff_7_n61) );
  NAND2_X1 md1FF_state_gff_7_U9 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[25]), 
        .ZN(md1FF_state_gff_7_n59) );
  NAND2_X1 md1FF_state_gff_7_U8 ( .A1(md1FF_state_gff_7_n58), .A2(
        md1FF_state_gff_7_n57), .ZN(md1FF_state_gff_7_n32) );
  NAND2_X1 md1FF_state_gff_7_U7 ( .A1(md1FF_state_gff_7_n67), .A2(
        md1FF_permOut[6]), .ZN(md1FF_state_gff_7_n57) );
  NOR2_X1 md1FF_state_gff_7_U6 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_7_n56), .ZN(md1FF_state_gff_7_n67) );
  MUX2_X1 md1FF_state_gff_7_U5 ( .A(md1FF_state_gff_7_n36), .B(
        md1FF_state_gff_7_n55), .S(md1FF_state_gff_7_n65), .Z(
        md1FF_state_gff_7_n58) );
  INV_X1 md1FF_state_gff_7_U4 ( .A(md1FF_state_gff_7_n56), .ZN(
        md1FF_state_gff_7_n65) );
  INV_X1 md1FF_state_gff_7_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_7_n56)
         );
  NAND2_X1 md1FF_state_gff_7_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[24]), 
        .ZN(md1FF_state_gff_7_n55) );
  DFF_X1 md1FF_state_gff_7_s_current_state_reg_0_ ( .D(md1FF_state_gff_7_n32), 
        .CK(clk), .Q(md1FF_permOut[7]), .QN(md1FF_state_gff_7_n36) );
  DFF_X1 md1FF_state_gff_7_s_current_state_reg_1_ ( .D(md1FF_state_gff_7_n31), 
        .CK(clk), .Q(md1FF_permOut[23]), .QN(md1FF_state_gff_7_n35) );
  DFF_X1 md1FF_state_gff_7_s_current_state_reg_2_ ( .D(md1FF_state_gff_7_n30), 
        .CK(clk), .Q(md1FF_permOut[39]), .QN(md1FF_state_gff_7_n34) );
  DFF_X1 md1FF_state_gff_7_s_current_state_reg_3_ ( .D(md1FF_state_gff_7_n29), 
        .CK(clk), .Q(md1FF_permOut[55]), .QN(md1FF_state_gff_7_n33) );
  NAND2_X1 md1FF_state_gff_8_U20 ( .A1(md1FF_state_gff_8_n69), .A2(
        md1FF_state_gff_8_n68), .ZN(md1FF_state_gff_8_n29) );
  NAND2_X1 md1FF_state_gff_8_U19 ( .A1(md1FF_state_gff_8_n67), .A2(
        md1FF_permOut[55]), .ZN(md1FF_state_gff_8_n68) );
  MUX2_X1 md1FF_state_gff_8_U18 ( .A(md1FF_state_gff_8_n33), .B(
        md1FF_state_gff_8_n66), .S(md1FF_state_gff_8_n65), .Z(
        md1FF_state_gff_8_n69) );
  NAND2_X1 md1FF_state_gff_8_U17 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[31]), .ZN(md1FF_state_gff_8_n66) );
  NAND2_X1 md1FF_state_gff_8_U16 ( .A1(md1FF_state_gff_8_n64), .A2(
        md1FF_state_gff_8_n63), .ZN(md1FF_state_gff_8_n30) );
  NAND2_X1 md1FF_state_gff_8_U15 ( .A1(md1FF_state_gff_8_n67), .A2(
        md1FF_permOut[39]), .ZN(md1FF_state_gff_8_n63) );
  MUX2_X1 md1FF_state_gff_8_U14 ( .A(md1FF_state_gff_8_n34), .B(
        md1FF_state_gff_8_n62), .S(md1FF_state_gff_8_n65), .Z(
        md1FF_state_gff_8_n64) );
  NAND2_X1 md1FF_state_gff_8_U13 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[30]), .ZN(md1FF_state_gff_8_n62) );
  NAND2_X1 md1FF_state_gff_8_U12 ( .A1(md1FF_state_gff_8_n61), .A2(
        md1FF_state_gff_8_n60), .ZN(md1FF_state_gff_8_n31) );
  NAND2_X1 md1FF_state_gff_8_U11 ( .A1(md1FF_state_gff_8_n67), .A2(
        md1FF_permOut[23]), .ZN(md1FF_state_gff_8_n60) );
  MUX2_X1 md1FF_state_gff_8_U10 ( .A(md1FF_state_gff_8_n35), .B(
        md1FF_state_gff_8_n59), .S(md1FF_state_gff_8_n65), .Z(
        md1FF_state_gff_8_n61) );
  NAND2_X1 md1FF_state_gff_8_U9 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[29]), .ZN(md1FF_state_gff_8_n59) );
  NAND2_X1 md1FF_state_gff_8_U8 ( .A1(md1FF_state_gff_8_n58), .A2(
        md1FF_state_gff_8_n57), .ZN(md1FF_state_gff_8_n32) );
  NAND2_X1 md1FF_state_gff_8_U7 ( .A1(md1FF_state_gff_8_n67), .A2(
        md1FF_permOut[7]), .ZN(md1FF_state_gff_8_n57) );
  NOR2_X1 md1FF_state_gff_8_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_8_n56), .ZN(md1FF_state_gff_8_n67) );
  MUX2_X1 md1FF_state_gff_8_U5 ( .A(md1FF_state_gff_8_n36), .B(
        md1FF_state_gff_8_n55), .S(md1FF_state_gff_8_n65), .Z(
        md1FF_state_gff_8_n58) );
  INV_X1 md1FF_state_gff_8_U4 ( .A(md1FF_state_gff_8_n56), .ZN(
        md1FF_state_gff_8_n65) );
  INV_X1 md1FF_state_gff_8_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_8_n56)
         );
  NAND2_X1 md1FF_state_gff_8_U2 ( .A1(md1FF_state_n10), .A2(md1FF_inputPar[28]), .ZN(md1FF_state_gff_8_n55) );
  DFF_X1 md1FF_state_gff_8_s_current_state_reg_0_ ( .D(md1FF_state_gff_8_n32), 
        .CK(clk), .Q(md1FF_permOut[8]), .QN(md1FF_state_gff_8_n36) );
  DFF_X1 md1FF_state_gff_8_s_current_state_reg_1_ ( .D(md1FF_state_gff_8_n31), 
        .CK(clk), .Q(md1FF_permOut[24]), .QN(md1FF_state_gff_8_n35) );
  DFF_X1 md1FF_state_gff_8_s_current_state_reg_2_ ( .D(md1FF_state_gff_8_n30), 
        .CK(clk), .Q(md1FF_permOut[40]), .QN(md1FF_state_gff_8_n34) );
  DFF_X1 md1FF_state_gff_8_s_current_state_reg_3_ ( .D(md1FF_state_gff_8_n29), 
        .CK(clk), .Q(md1FF_permOut[56]), .QN(md1FF_state_gff_8_n33) );
  NAND2_X1 md1FF_state_gff_9_U20 ( .A1(md1FF_state_gff_9_n69), .A2(
        md1FF_state_gff_9_n68), .ZN(md1FF_state_gff_9_n29) );
  NAND2_X1 md1FF_state_gff_9_U19 ( .A1(md1FF_state_gff_9_n67), .A2(
        md1FF_permOut[56]), .ZN(md1FF_state_gff_9_n68) );
  MUX2_X1 md1FF_state_gff_9_U18 ( .A(md1FF_state_gff_9_n33), .B(
        md1FF_state_gff_9_n66), .S(md1FF_state_gff_9_n65), .Z(
        md1FF_state_gff_9_n69) );
  NAND2_X1 md1FF_state_gff_9_U17 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[35]), .ZN(md1FF_state_gff_9_n66) );
  NAND2_X1 md1FF_state_gff_9_U16 ( .A1(md1FF_state_gff_9_n64), .A2(
        md1FF_state_gff_9_n63), .ZN(md1FF_state_gff_9_n30) );
  NAND2_X1 md1FF_state_gff_9_U15 ( .A1(md1FF_state_gff_9_n67), .A2(
        md1FF_permOut[40]), .ZN(md1FF_state_gff_9_n63) );
  MUX2_X1 md1FF_state_gff_9_U14 ( .A(md1FF_state_gff_9_n34), .B(
        md1FF_state_gff_9_n62), .S(md1FF_state_gff_9_n65), .Z(
        md1FF_state_gff_9_n64) );
  NAND2_X1 md1FF_state_gff_9_U13 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[34]), .ZN(md1FF_state_gff_9_n62) );
  NAND2_X1 md1FF_state_gff_9_U12 ( .A1(md1FF_state_gff_9_n61), .A2(
        md1FF_state_gff_9_n60), .ZN(md1FF_state_gff_9_n31) );
  NAND2_X1 md1FF_state_gff_9_U11 ( .A1(md1FF_state_gff_9_n67), .A2(
        md1FF_permOut[24]), .ZN(md1FF_state_gff_9_n60) );
  MUX2_X1 md1FF_state_gff_9_U10 ( .A(md1FF_state_gff_9_n35), .B(
        md1FF_state_gff_9_n59), .S(md1FF_state_gff_9_n65), .Z(
        md1FF_state_gff_9_n61) );
  NAND2_X1 md1FF_state_gff_9_U9 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[33]), 
        .ZN(md1FF_state_gff_9_n59) );
  NAND2_X1 md1FF_state_gff_9_U8 ( .A1(md1FF_state_gff_9_n58), .A2(
        md1FF_state_gff_9_n57), .ZN(md1FF_state_gff_9_n32) );
  NAND2_X1 md1FF_state_gff_9_U7 ( .A1(md1FF_state_gff_9_n67), .A2(
        md1FF_permOut[8]), .ZN(md1FF_state_gff_9_n57) );
  NOR2_X1 md1FF_state_gff_9_U6 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_9_n56), .ZN(md1FF_state_gff_9_n67) );
  MUX2_X1 md1FF_state_gff_9_U5 ( .A(md1FF_state_gff_9_n36), .B(
        md1FF_state_gff_9_n55), .S(md1FF_state_gff_9_n65), .Z(
        md1FF_state_gff_9_n58) );
  INV_X1 md1FF_state_gff_9_U4 ( .A(md1FF_state_gff_9_n56), .ZN(
        md1FF_state_gff_9_n65) );
  INV_X1 md1FF_state_gff_9_U3 ( .A(md1FF_state_n7), .ZN(md1FF_state_gff_9_n56)
         );
  NAND2_X1 md1FF_state_gff_9_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[32]), 
        .ZN(md1FF_state_gff_9_n55) );
  DFF_X1 md1FF_state_gff_9_s_current_state_reg_0_ ( .D(md1FF_state_gff_9_n32), 
        .CK(clk), .Q(md1FF_permOut[9]), .QN(md1FF_state_gff_9_n36) );
  DFF_X1 md1FF_state_gff_9_s_current_state_reg_1_ ( .D(md1FF_state_gff_9_n31), 
        .CK(clk), .Q(md1FF_permOut[25]), .QN(md1FF_state_gff_9_n35) );
  DFF_X1 md1FF_state_gff_9_s_current_state_reg_2_ ( .D(md1FF_state_gff_9_n30), 
        .CK(clk), .Q(md1FF_permOut[41]), .QN(md1FF_state_gff_9_n34) );
  DFF_X1 md1FF_state_gff_9_s_current_state_reg_3_ ( .D(md1FF_state_gff_9_n29), 
        .CK(clk), .Q(md1FF_permOut[57]), .QN(md1FF_state_gff_9_n33) );
  NAND2_X1 md1FF_state_gff_10_U20 ( .A1(md1FF_state_gff_10_n69), .A2(
        md1FF_state_gff_10_n68), .ZN(md1FF_state_gff_10_n29) );
  NAND2_X1 md1FF_state_gff_10_U19 ( .A1(md1FF_state_gff_10_n67), .A2(
        md1FF_permOut[57]), .ZN(md1FF_state_gff_10_n68) );
  MUX2_X1 md1FF_state_gff_10_U18 ( .A(md1FF_state_gff_10_n33), .B(
        md1FF_state_gff_10_n66), .S(md1FF_state_gff_10_n65), .Z(
        md1FF_state_gff_10_n69) );
  NAND2_X1 md1FF_state_gff_10_U17 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[39]), .ZN(md1FF_state_gff_10_n66) );
  NAND2_X1 md1FF_state_gff_10_U16 ( .A1(md1FF_state_gff_10_n64), .A2(
        md1FF_state_gff_10_n63), .ZN(md1FF_state_gff_10_n30) );
  NAND2_X1 md1FF_state_gff_10_U15 ( .A1(md1FF_state_gff_10_n67), .A2(
        md1FF_permOut[41]), .ZN(md1FF_state_gff_10_n63) );
  MUX2_X1 md1FF_state_gff_10_U14 ( .A(md1FF_state_gff_10_n34), .B(
        md1FF_state_gff_10_n62), .S(md1FF_state_gff_10_n65), .Z(
        md1FF_state_gff_10_n64) );
  NAND2_X1 md1FF_state_gff_10_U13 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[38]), .ZN(md1FF_state_gff_10_n62) );
  NAND2_X1 md1FF_state_gff_10_U12 ( .A1(md1FF_state_gff_10_n61), .A2(
        md1FF_state_gff_10_n60), .ZN(md1FF_state_gff_10_n31) );
  NAND2_X1 md1FF_state_gff_10_U11 ( .A1(md1FF_state_gff_10_n67), .A2(
        md1FF_permOut[25]), .ZN(md1FF_state_gff_10_n60) );
  MUX2_X1 md1FF_state_gff_10_U10 ( .A(md1FF_state_gff_10_n35), .B(
        md1FF_state_gff_10_n59), .S(md1FF_state_gff_10_n65), .Z(
        md1FF_state_gff_10_n61) );
  NAND2_X1 md1FF_state_gff_10_U9 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[37]), .ZN(md1FF_state_gff_10_n59) );
  NAND2_X1 md1FF_state_gff_10_U8 ( .A1(md1FF_state_gff_10_n58), .A2(
        md1FF_state_gff_10_n57), .ZN(md1FF_state_gff_10_n32) );
  NAND2_X1 md1FF_state_gff_10_U7 ( .A1(md1FF_state_gff_10_n67), .A2(
        md1FF_permOut[9]), .ZN(md1FF_state_gff_10_n57) );
  NOR2_X1 md1FF_state_gff_10_U6 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_10_n56), .ZN(md1FF_state_gff_10_n67) );
  MUX2_X1 md1FF_state_gff_10_U5 ( .A(md1FF_state_gff_10_n36), .B(
        md1FF_state_gff_10_n55), .S(md1FF_state_gff_10_n65), .Z(
        md1FF_state_gff_10_n58) );
  INV_X1 md1FF_state_gff_10_U4 ( .A(md1FF_state_gff_10_n56), .ZN(
        md1FF_state_gff_10_n65) );
  INV_X1 md1FF_state_gff_10_U3 ( .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_10_n56) );
  NAND2_X1 md1FF_state_gff_10_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[36]), .ZN(md1FF_state_gff_10_n55) );
DFF_X1 md1FF_state_gff_10_s_current_state_reg_0_ ( .D(md1FF_state_gff_10_n32), .CK(clk), .Q(md1FF_permOut[10]), .QN(md1FF_state_gff_10_n36) );
DFF_X1 md1FF_state_gff_10_s_current_state_reg_1_ ( .D(md1FF_state_gff_10_n31), .CK(clk), .Q(md1FF_permOut[26]), .QN(md1FF_state_gff_10_n35) );
DFF_X1 md1FF_state_gff_10_s_current_state_reg_2_ ( .D(md1FF_state_gff_10_n30), .CK(clk), .Q(md1FF_permOut[42]), .QN(md1FF_state_gff_10_n34) );
DFF_X1 md1FF_state_gff_10_s_current_state_reg_3_ ( .D(md1FF_state_gff_10_n29), .CK(clk), .Q(md1FF_permOut[58]), .QN(md1FF_state_gff_10_n33) );
  NAND2_X1 md1FF_state_gff_11_U20 ( .A1(md1FF_state_gff_11_n69), .A2(
        md1FF_state_gff_11_n68), .ZN(md1FF_state_gff_11_n29) );
  NAND2_X1 md1FF_state_gff_11_U19 ( .A1(md1FF_state_gff_11_n67), .A2(
        md1FF_permOut[58]), .ZN(md1FF_state_gff_11_n68) );
  MUX2_X1 md1FF_state_gff_11_U18 ( .A(md1FF_state_gff_11_n33), .B(
        md1FF_state_gff_11_n66), .S(md1FF_state_gff_11_n65), .Z(
        md1FF_state_gff_11_n69) );
  NAND2_X1 md1FF_state_gff_11_U17 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[43]), .ZN(md1FF_state_gff_11_n66) );
  NAND2_X1 md1FF_state_gff_11_U16 ( .A1(md1FF_state_gff_11_n64), .A2(
        md1FF_state_gff_11_n63), .ZN(md1FF_state_gff_11_n30) );
  NAND2_X1 md1FF_state_gff_11_U15 ( .A1(md1FF_state_gff_11_n67), .A2(
        md1FF_permOut[42]), .ZN(md1FF_state_gff_11_n63) );
  MUX2_X1 md1FF_state_gff_11_U14 ( .A(md1FF_state_gff_11_n34), .B(
        md1FF_state_gff_11_n62), .S(md1FF_state_gff_11_n65), .Z(
        md1FF_state_gff_11_n64) );
  NAND2_X1 md1FF_state_gff_11_U13 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[42]), .ZN(md1FF_state_gff_11_n62) );
  NAND2_X1 md1FF_state_gff_11_U12 ( .A1(md1FF_state_gff_11_n61), .A2(
        md1FF_state_gff_11_n60), .ZN(md1FF_state_gff_11_n31) );
  NAND2_X1 md1FF_state_gff_11_U11 ( .A1(md1FF_state_gff_11_n67), .A2(
        md1FF_permOut[26]), .ZN(md1FF_state_gff_11_n60) );
  MUX2_X1 md1FF_state_gff_11_U10 ( .A(md1FF_state_gff_11_n35), .B(
        md1FF_state_gff_11_n59), .S(md1FF_state_gff_11_n65), .Z(
        md1FF_state_gff_11_n61) );
  NAND2_X1 md1FF_state_gff_11_U9 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[41]), .ZN(md1FF_state_gff_11_n59) );
  NAND2_X1 md1FF_state_gff_11_U8 ( .A1(md1FF_state_gff_11_n58), .A2(
        md1FF_state_gff_11_n57), .ZN(md1FF_state_gff_11_n32) );
  NAND2_X1 md1FF_state_gff_11_U7 ( .A1(md1FF_state_gff_11_n67), .A2(
        md1FF_permOut[10]), .ZN(md1FF_state_gff_11_n57) );
  NOR2_X1 md1FF_state_gff_11_U6 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_11_n56), .ZN(md1FF_state_gff_11_n67) );
  MUX2_X1 md1FF_state_gff_11_U5 ( .A(md1FF_state_gff_11_n36), .B(
        md1FF_state_gff_11_n55), .S(md1FF_state_gff_11_n65), .Z(
        md1FF_state_gff_11_n58) );
  INV_X1 md1FF_state_gff_11_U4 ( .A(md1FF_state_gff_11_n56), .ZN(
        md1FF_state_gff_11_n65) );
  INV_X1 md1FF_state_gff_11_U3 ( .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_11_n56) );
  NAND2_X1 md1FF_state_gff_11_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[40]), .ZN(md1FF_state_gff_11_n55) );
DFF_X1 md1FF_state_gff_11_s_current_state_reg_0_ ( .D(md1FF_state_gff_11_n32), .CK(clk), .Q(md1FF_permOut[11]), .QN(md1FF_state_gff_11_n36) );
DFF_X1 md1FF_state_gff_11_s_current_state_reg_1_ ( .D(md1FF_state_gff_11_n31), .CK(clk), .Q(md1FF_permOut[27]), .QN(md1FF_state_gff_11_n35) );
DFF_X1 md1FF_state_gff_11_s_current_state_reg_2_ ( .D(md1FF_state_gff_11_n30), .CK(clk), .Q(md1FF_permOut[43]), .QN(md1FF_state_gff_11_n34) );
DFF_X1 md1FF_state_gff_11_s_current_state_reg_3_ ( .D(md1FF_state_gff_11_n29), .CK(clk), .Q(md1FF_permOut[59]), .QN(md1FF_state_gff_11_n33) );
  NAND2_X1 md1FF_state_gff_12_U20 ( .A1(md1FF_state_gff_12_n69), .A2(
        md1FF_state_gff_12_n68), .ZN(md1FF_state_gff_12_n29) );
  NAND2_X1 md1FF_state_gff_12_U19 ( .A1(md1FF_state_gff_12_n67), .A2(
        md1FF_permOut[59]), .ZN(md1FF_state_gff_12_n68) );
  MUX2_X1 md1FF_state_gff_12_U18 ( .A(md1FF_state_gff_12_n33), .B(
        md1FF_state_gff_12_n66), .S(md1FF_state_gff_12_n65), .Z(
        md1FF_state_gff_12_n69) );
  NAND2_X1 md1FF_state_gff_12_U17 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[47]), .ZN(md1FF_state_gff_12_n66) );
  NAND2_X1 md1FF_state_gff_12_U16 ( .A1(md1FF_state_gff_12_n64), .A2(
        md1FF_state_gff_12_n63), .ZN(md1FF_state_gff_12_n30) );
  NAND2_X1 md1FF_state_gff_12_U15 ( .A1(md1FF_state_gff_12_n67), .A2(
        md1FF_permOut[43]), .ZN(md1FF_state_gff_12_n63) );
  MUX2_X1 md1FF_state_gff_12_U14 ( .A(md1FF_state_gff_12_n34), .B(
        md1FF_state_gff_12_n62), .S(md1FF_state_gff_12_n65), .Z(
        md1FF_state_gff_12_n64) );
  NAND2_X1 md1FF_state_gff_12_U13 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[46]), .ZN(md1FF_state_gff_12_n62) );
  NAND2_X1 md1FF_state_gff_12_U12 ( .A1(md1FF_state_gff_12_n61), .A2(
        md1FF_state_gff_12_n60), .ZN(md1FF_state_gff_12_n31) );
  NAND2_X1 md1FF_state_gff_12_U11 ( .A1(md1FF_state_gff_12_n67), .A2(
        md1FF_permOut[27]), .ZN(md1FF_state_gff_12_n60) );
  MUX2_X1 md1FF_state_gff_12_U10 ( .A(md1FF_state_gff_12_n35), .B(
        md1FF_state_gff_12_n59), .S(md1FF_state_gff_12_n65), .Z(
        md1FF_state_gff_12_n61) );
  NAND2_X1 md1FF_state_gff_12_U9 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[45]), .ZN(md1FF_state_gff_12_n59) );
  NAND2_X1 md1FF_state_gff_12_U8 ( .A1(md1FF_state_gff_12_n58), .A2(
        md1FF_state_gff_12_n57), .ZN(md1FF_state_gff_12_n32) );
  NAND2_X1 md1FF_state_gff_12_U7 ( .A1(md1FF_state_gff_12_n67), .A2(
        md1FF_permOut[11]), .ZN(md1FF_state_gff_12_n57) );
  NOR2_X1 md1FF_state_gff_12_U6 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_12_n56), .ZN(md1FF_state_gff_12_n67) );
  MUX2_X1 md1FF_state_gff_12_U5 ( .A(md1FF_state_gff_12_n36), .B(
        md1FF_state_gff_12_n55), .S(md1FF_state_gff_12_n65), .Z(
        md1FF_state_gff_12_n58) );
  INV_X1 md1FF_state_gff_12_U4 ( .A(md1FF_state_gff_12_n56), .ZN(
        md1FF_state_gff_12_n65) );
  INV_X1 md1FF_state_gff_12_U3 ( .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_12_n56) );
  NAND2_X1 md1FF_state_gff_12_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[44]), .ZN(md1FF_state_gff_12_n55) );
DFF_X1 md1FF_state_gff_12_s_current_state_reg_0_ ( .D(md1FF_state_gff_12_n32), .CK(clk), .Q(md1FF_permOut[12]), .QN(md1FF_state_gff_12_n36) );
DFF_X1 md1FF_state_gff_12_s_current_state_reg_1_ ( .D(md1FF_state_gff_12_n31), .CK(clk), .Q(md1FF_permOut[28]), .QN(md1FF_state_gff_12_n35) );
DFF_X1 md1FF_state_gff_12_s_current_state_reg_2_ ( .D(md1FF_state_gff_12_n30), .CK(clk), .Q(md1FF_permOut[44]), .QN(md1FF_state_gff_12_n34) );
DFF_X1 md1FF_state_gff_12_s_current_state_reg_3_ ( .D(md1FF_state_gff_12_n29), .CK(clk), .Q(md1FF_permOut[60]), .QN(md1FF_state_gff_12_n33) );
  NAND2_X1 md1FF_state_gff_13_U20 ( .A1(md1FF_state_gff_13_n69), .A2(
        md1FF_state_gff_13_n68), .ZN(md1FF_state_gff_13_n29) );
  NAND2_X1 md1FF_state_gff_13_U19 ( .A1(md1FF_state_gff_13_n67), .A2(
        md1FF_permOut[60]), .ZN(md1FF_state_gff_13_n68) );
  MUX2_X1 md1FF_state_gff_13_U18 ( .A(md1FF_state_gff_13_n33), .B(
        md1FF_state_gff_13_n66), .S(md1FF_state_gff_13_n65), .Z(
        md1FF_state_gff_13_n69) );
  NAND2_X1 md1FF_state_gff_13_U17 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[51]), .ZN(md1FF_state_gff_13_n66) );
  NAND2_X1 md1FF_state_gff_13_U16 ( .A1(md1FF_state_gff_13_n64), .A2(
        md1FF_state_gff_13_n63), .ZN(md1FF_state_gff_13_n30) );
  NAND2_X1 md1FF_state_gff_13_U15 ( .A1(md1FF_state_gff_13_n67), .A2(
        md1FF_permOut[44]), .ZN(md1FF_state_gff_13_n63) );
  MUX2_X1 md1FF_state_gff_13_U14 ( .A(md1FF_state_gff_13_n34), .B(
        md1FF_state_gff_13_n62), .S(md1FF_state_gff_13_n65), .Z(
        md1FF_state_gff_13_n64) );
  NAND2_X1 md1FF_state_gff_13_U13 ( .A1(md1FF_state_n9), .A2(
        md1FF_inputPar[50]), .ZN(md1FF_state_gff_13_n62) );
  NAND2_X1 md1FF_state_gff_13_U12 ( .A1(md1FF_state_gff_13_n61), .A2(
        md1FF_state_gff_13_n60), .ZN(md1FF_state_gff_13_n31) );
  NAND2_X1 md1FF_state_gff_13_U11 ( .A1(md1FF_state_gff_13_n67), .A2(
        md1FF_permOut[28]), .ZN(md1FF_state_gff_13_n60) );
  MUX2_X1 md1FF_state_gff_13_U10 ( .A(md1FF_state_gff_13_n35), .B(
        md1FF_state_gff_13_n59), .S(md1FF_state_gff_13_n65), .Z(
        md1FF_state_gff_13_n61) );
  NAND2_X1 md1FF_state_gff_13_U9 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[49]), .ZN(md1FF_state_gff_13_n59) );
  NAND2_X1 md1FF_state_gff_13_U8 ( .A1(md1FF_state_gff_13_n58), .A2(
        md1FF_state_gff_13_n57), .ZN(md1FF_state_gff_13_n32) );
  NAND2_X1 md1FF_state_gff_13_U7 ( .A1(md1FF_state_gff_13_n67), .A2(
        md1FF_permOut[12]), .ZN(md1FF_state_gff_13_n57) );
  NOR2_X1 md1FF_state_gff_13_U6 ( .A1(md1FF_state_n9), .A2(
        md1FF_state_gff_13_n56), .ZN(md1FF_state_gff_13_n67) );
  MUX2_X1 md1FF_state_gff_13_U5 ( .A(md1FF_state_gff_13_n36), .B(
        md1FF_state_gff_13_n55), .S(md1FF_state_gff_13_n65), .Z(
        md1FF_state_gff_13_n58) );
  INV_X1 md1FF_state_gff_13_U4 ( .A(md1FF_state_gff_13_n56), .ZN(
        md1FF_state_gff_13_n65) );
  INV_X1 md1FF_state_gff_13_U3 ( .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_13_n56) );
  NAND2_X1 md1FF_state_gff_13_U2 ( .A1(md1FF_state_n9), .A2(md1FF_inputPar[48]), .ZN(md1FF_state_gff_13_n55) );
DFF_X1 md1FF_state_gff_13_s_current_state_reg_0_ ( .D(md1FF_state_gff_13_n32), .CK(clk), .Q(md1FF_permOut[13]), .QN(md1FF_state_gff_13_n36) );
DFF_X1 md1FF_state_gff_13_s_current_state_reg_1_ ( .D(md1FF_state_gff_13_n31), .CK(clk), .Q(md1FF_permOut[29]), .QN(md1FF_state_gff_13_n35) );
DFF_X1 md1FF_state_gff_13_s_current_state_reg_2_ ( .D(md1FF_state_gff_13_n30), .CK(clk), .Q(md1FF_permOut[45]), .QN(md1FF_state_gff_13_n34) );
DFF_X1 md1FF_state_gff_13_s_current_state_reg_3_ ( .D(md1FF_state_gff_13_n29), .CK(clk), .Q(md1FF_permOut[61]), .QN(md1FF_state_gff_13_n33) );
  NAND2_X1 md1FF_state_gff_14_U20 ( .A1(md1FF_state_gff_14_n69), .A2(
        md1FF_state_gff_14_n68), .ZN(md1FF_state_gff_14_n29) );
  NAND2_X1 md1FF_state_gff_14_U19 ( .A1(md1FF_state_gff_14_n67), .A2(
        md1FF_permOut[61]), .ZN(md1FF_state_gff_14_n68) );
  MUX2_X1 md1FF_state_gff_14_U18 ( .A(md1FF_state_gff_14_n33), .B(
        md1FF_state_gff_14_n66), .S(md1FF_state_gff_14_n65), .Z(
        md1FF_state_gff_14_n69) );
  NAND2_X1 md1FF_state_gff_14_U17 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[55]), .ZN(md1FF_state_gff_14_n66) );
  NAND2_X1 md1FF_state_gff_14_U16 ( .A1(md1FF_state_gff_14_n64), .A2(
        md1FF_state_gff_14_n63), .ZN(md1FF_state_gff_14_n30) );
  NAND2_X1 md1FF_state_gff_14_U15 ( .A1(md1FF_state_gff_14_n67), .A2(
        md1FF_permOut[45]), .ZN(md1FF_state_gff_14_n63) );
  MUX2_X1 md1FF_state_gff_14_U14 ( .A(md1FF_state_gff_14_n34), .B(
        md1FF_state_gff_14_n62), .S(md1FF_state_gff_14_n65), .Z(
        md1FF_state_gff_14_n64) );
  NAND2_X1 md1FF_state_gff_14_U13 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[54]), .ZN(md1FF_state_gff_14_n62) );
  NAND2_X1 md1FF_state_gff_14_U12 ( .A1(md1FF_state_gff_14_n61), .A2(
        md1FF_state_gff_14_n60), .ZN(md1FF_state_gff_14_n31) );
  NAND2_X1 md1FF_state_gff_14_U11 ( .A1(md1FF_state_gff_14_n67), .A2(
        md1FF_permOut[29]), .ZN(md1FF_state_gff_14_n60) );
  MUX2_X1 md1FF_state_gff_14_U10 ( .A(md1FF_state_gff_14_n35), .B(
        md1FF_state_gff_14_n59), .S(md1FF_state_gff_14_n65), .Z(
        md1FF_state_gff_14_n61) );
  NAND2_X1 md1FF_state_gff_14_U9 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[53]), .ZN(md1FF_state_gff_14_n59) );
  NAND2_X1 md1FF_state_gff_14_U8 ( .A1(md1FF_state_gff_14_n58), .A2(
        md1FF_state_gff_14_n57), .ZN(md1FF_state_gff_14_n32) );
  NAND2_X1 md1FF_state_gff_14_U7 ( .A1(md1FF_state_gff_14_n67), .A2(
        md1FF_permOut[13]), .ZN(md1FF_state_gff_14_n57) );
  NOR2_X1 md1FF_state_gff_14_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_14_n56), .ZN(md1FF_state_gff_14_n67) );
  MUX2_X1 md1FF_state_gff_14_U5 ( .A(md1FF_state_gff_14_n36), .B(
        md1FF_state_gff_14_n55), .S(md1FF_state_gff_14_n65), .Z(
        md1FF_state_gff_14_n58) );
  INV_X1 md1FF_state_gff_14_U4 ( .A(md1FF_state_gff_14_n56), .ZN(
        md1FF_state_gff_14_n65) );
  INV_X1 md1FF_state_gff_14_U3 ( .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_14_n56) );
  NAND2_X1 md1FF_state_gff_14_U2 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[52]), .ZN(md1FF_state_gff_14_n55) );
DFF_X1 md1FF_state_gff_14_s_current_state_reg_0_ ( .D(md1FF_state_gff_14_n32), .CK(clk), .Q(md1FF_permOut[14]), .QN(md1FF_state_gff_14_n36) );
DFF_X1 md1FF_state_gff_14_s_current_state_reg_1_ ( .D(md1FF_state_gff_14_n31), .CK(clk), .Q(md1FF_permOut[30]), .QN(md1FF_state_gff_14_n35) );
DFF_X1 md1FF_state_gff_14_s_current_state_reg_2_ ( .D(md1FF_state_gff_14_n30), .CK(clk), .Q(md1FF_permOut[46]), .QN(md1FF_state_gff_14_n34) );
DFF_X1 md1FF_state_gff_14_s_current_state_reg_3_ ( .D(md1FF_state_gff_14_n29), .CK(clk), .Q(md1FF_permOut[62]), .QN(md1FF_state_gff_14_n33) );
  NAND2_X1 md1FF_state_gff_15_U20 ( .A1(md1FF_state_gff_15_n68), .A2(
        md1FF_state_gff_15_n67), .ZN(md1FF_state_gff_15_n28) );
  NAND2_X1 md1FF_state_gff_15_U19 ( .A1(md1FF_state_gff_15_n66), .A2(
        md1FF_permOut[62]), .ZN(md1FF_state_gff_15_n67) );
  MUX2_X1 md1FF_state_gff_15_U18 ( .A(md1FF_state_gff_15_n32), .B(
        md1FF_state_gff_15_n65), .S(md1FF_state_gff_15_n64), .Z(
        md1FF_state_gff_15_n68) );
  NAND2_X1 md1FF_state_gff_15_U17 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[59]), .ZN(md1FF_state_gff_15_n65) );
  NAND2_X1 md1FF_state_gff_15_U16 ( .A1(md1FF_state_gff_15_n63), .A2(
        md1FF_state_gff_15_n62), .ZN(md1FF_state_gff_15_n29) );
  NAND2_X1 md1FF_state_gff_15_U15 ( .A1(md1FF_state_gff_15_n66), .A2(
        md1FF_permOut[46]), .ZN(md1FF_state_gff_15_n62) );
  MUX2_X1 md1FF_state_gff_15_U14 ( .A(md1FF_state_gff_15_n33), .B(
        md1FF_state_gff_15_n61), .S(md1FF_state_gff_15_n64), .Z(
        md1FF_state_gff_15_n63) );
  NAND2_X1 md1FF_state_gff_15_U13 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[58]), .ZN(md1FF_state_gff_15_n61) );
  NAND2_X1 md1FF_state_gff_15_U12 ( .A1(md1FF_state_gff_15_n60), .A2(
        md1FF_state_gff_15_n59), .ZN(md1FF_state_gff_15_n30) );
  NAND2_X1 md1FF_state_gff_15_U11 ( .A1(md1FF_state_gff_15_n66), .A2(
        md1FF_permOut[30]), .ZN(md1FF_state_gff_15_n59) );
  MUX2_X1 md1FF_state_gff_15_U10 ( .A(md1FF_state_gff_15_n34), .B(
        md1FF_state_gff_15_n58), .S(md1FF_state_gff_15_n64), .Z(
        md1FF_state_gff_15_n60) );
  NAND2_X1 md1FF_state_gff_15_U9 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[57]), .ZN(md1FF_state_gff_15_n58) );
  NAND2_X1 md1FF_state_gff_15_U8 ( .A1(md1FF_state_gff_15_n57), .A2(
        md1FF_state_gff_15_n56), .ZN(md1FF_state_gff_15_n31) );
  NAND2_X1 md1FF_state_gff_15_U7 ( .A1(md1FF_state_gff_15_n66), .A2(
        md1FF_permOut[14]), .ZN(md1FF_state_gff_15_n56) );
  NOR2_X1 md1FF_state_gff_15_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_15_n55), .ZN(md1FF_state_gff_15_n66) );
  MUX2_X1 md1FF_state_gff_15_U5 ( .A(md1FF_state_gff_15_n35), .B(
        md1FF_state_gff_15_n54), .S(md1FF_state_gff_15_n64), .Z(
        md1FF_state_gff_15_n57) );
  INV_X1 md1FF_state_gff_15_U4 ( .A(md1FF_state_gff_15_n55), .ZN(
        md1FF_state_gff_15_n64) );
  INV_X1 md1FF_state_gff_15_U3 ( .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_15_n55) );
  NAND2_X1 md1FF_state_gff_15_U2 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[56]), .ZN(md1FF_state_gff_15_n54) );
DFF_X1 md1FF_state_gff_15_s_current_state_reg_0_ ( .D(md1FF_state_gff_15_n31), .CK(clk), .Q(md1FF_permOut[15]), .QN(md1FF_state_gff_15_n35) );
DFF_X1 md1FF_state_gff_15_s_current_state_reg_1_ ( .D(md1FF_state_gff_15_n30), .CK(clk), .Q(md1FF_permOut[31]), .QN(md1FF_state_gff_15_n34) );
DFF_X1 md1FF_state_gff_15_s_current_state_reg_2_ ( .D(md1FF_state_gff_15_n29), .CK(clk), .Q(md1FF_permOut[47]), .QN(md1FF_state_gff_15_n33) );
DFF_X1 md1FF_state_gff_15_s_current_state_reg_3_ ( .D(md1FF_state_gff_15_n28), .CK(clk), .Q(md1FF_permOut[63]), .QN(md1FF_state_gff_15_n32) );
  NAND2_X1 md1FF_state_gff_16_U20 ( .A1(md1FF_state_gff_16_n68), .A2(
        md1FF_state_gff_16_n67), .ZN(md1FF_state_gff_16_n28) );
  NAND2_X1 md1FF_state_gff_16_U19 ( .A1(md1FF_state_gff_16_n66), .A2(
        md1FF_permOut[63]), .ZN(md1FF_state_gff_16_n67) );
  MUX2_X1 md1FF_state_gff_16_U18 ( .A(md1FF_state_gff_16_n32), .B(
        md1FF_state_gff_16_n65), .S(md1FF_state_gff_16_n64), .Z(
        md1FF_state_gff_16_n68) );
  NAND2_X1 md1FF_state_gff_16_U17 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[63]), .ZN(md1FF_state_gff_16_n65) );
  NAND2_X1 md1FF_state_gff_16_U16 ( .A1(md1FF_state_gff_16_n63), .A2(
        md1FF_state_gff_16_n62), .ZN(md1FF_state_gff_16_n29) );
  NAND2_X1 md1FF_state_gff_16_U15 ( .A1(md1FF_state_gff_16_n66), .A2(
        md1FF_permOut[47]), .ZN(md1FF_state_gff_16_n62) );
  MUX2_X1 md1FF_state_gff_16_U14 ( .A(md1FF_state_gff_16_n33), .B(
        md1FF_state_gff_16_n61), .S(md1FF_state_gff_16_n64), .Z(
        md1FF_state_gff_16_n63) );
  NAND2_X1 md1FF_state_gff_16_U13 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[62]), .ZN(md1FF_state_gff_16_n61) );
  NAND2_X1 md1FF_state_gff_16_U12 ( .A1(md1FF_state_gff_16_n60), .A2(
        md1FF_state_gff_16_n59), .ZN(md1FF_state_gff_16_n30) );
  NAND2_X1 md1FF_state_gff_16_U11 ( .A1(md1FF_state_gff_16_n66), .A2(
        md1FF_permOut[31]), .ZN(md1FF_state_gff_16_n59) );
  MUX2_X1 md1FF_state_gff_16_U10 ( .A(md1FF_state_gff_16_n34), .B(
        md1FF_state_gff_16_n58), .S(md1FF_state_gff_16_n64), .Z(
        md1FF_state_gff_16_n60) );
  NAND2_X1 md1FF_state_gff_16_U9 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[61]), .ZN(md1FF_state_gff_16_n58) );
  NAND2_X1 md1FF_state_gff_16_U8 ( .A1(md1FF_state_gff_16_n57), .A2(
        md1FF_state_gff_16_n56), .ZN(md1FF_state_gff_16_n31) );
  NAND2_X1 md1FF_state_gff_16_U7 ( .A1(md1FF_state_gff_16_n66), .A2(
        md1FF_permOut[15]), .ZN(md1FF_state_gff_16_n56) );
  NOR2_X1 md1FF_state_gff_16_U6 ( .A1(md1FF_state_n10), .A2(
        md1FF_state_gff_16_n55), .ZN(md1FF_state_gff_16_n66) );
  MUX2_X1 md1FF_state_gff_16_U5 ( .A(md1FF_state_gff_16_n35), .B(
        md1FF_state_gff_16_n54), .S(md1FF_state_gff_16_n64), .Z(
        md1FF_state_gff_16_n57) );
  INV_X1 md1FF_state_gff_16_U4 ( .A(md1FF_state_gff_16_n55), .ZN(
        md1FF_state_gff_16_n64) );
  INV_X1 md1FF_state_gff_16_U3 ( .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_16_n55) );
  NAND2_X1 md1FF_state_gff_16_U2 ( .A1(md1FF_state_n10), .A2(
        md1FF_inputPar[60]), .ZN(md1FF_state_gff_16_n54) );
DFF_X1 md1FF_state_gff_16_s_current_state_reg_0_ ( .D(md1FF_state_gff_16_n31), .CK(clk), .Q(md1Reg[0]), .QN(md1FF_state_gff_16_n35) );
DFF_X1 md1FF_state_gff_16_s_current_state_reg_1_ ( .D(md1FF_state_gff_16_n30), .CK(clk), .Q(md1Reg[1]), .QN(md1FF_state_gff_16_n34) );
DFF_X1 md1FF_state_gff_16_s_current_state_reg_2_ ( .D(md1FF_state_gff_16_n29), .CK(clk), .Q(md1Reg[2]), .QN(md1FF_state_gff_16_n33) );
DFF_X1 md1FF_state_gff_16_s_current_state_reg_3_ ( .D(md1FF_state_gff_16_n28), .CK(clk), .Q(md1Reg[3]), .QN(md1FF_state_gff_16_n32) );
  MUX2_X1 md2FF_U70 ( .A(md2FF_permOut[9]), .B(data_in3[9]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[9]) );
  MUX2_X1 md2FF_U69 ( .A(md2FF_permOut[8]), .B(data_in3[8]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[8]) );
  MUX2_X1 md2FF_U68 ( .A(md2FF_permOut[7]), .B(data_in3[7]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[7]) );
  MUX2_X1 md2FF_U67 ( .A(md2FF_permOut[6]), .B(data_in3[6]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[6]) );
  MUX2_X1 md2FF_U66 ( .A(md2FF_permOut[5]), .B(data_in3[5]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[5]) );
  MUX2_X1 md2FF_U65 ( .A(md2FF_permOut[4]), .B(data_in3[4]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[4]) );
  MUX2_X1 md2FF_U64 ( .A(md2FF_permOut[63]), .B(data_in3[63]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[63]) );
  MUX2_X1 md2FF_U63 ( .A(md2FF_permOut[62]), .B(data_in3[62]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[62]) );
  MUX2_X1 md2FF_U62 ( .A(md2FF_permOut[61]), .B(data_in3[61]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[61]) );
  MUX2_X1 md2FF_U61 ( .A(md2FF_permOut[60]), .B(data_in3[60]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[60]) );
  MUX2_X1 md2FF_U60 ( .A(md2FF_permOut[59]), .B(data_in3[59]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[59]) );
  MUX2_X1 md2FF_U59 ( .A(md2FF_permOut[58]), .B(data_in3[58]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[58]) );
  MUX2_X1 md2FF_U58 ( .A(md2FF_permOut[57]), .B(data_in3[57]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[57]) );
  MUX2_X1 md2FF_U57 ( .A(md2FF_permOut[56]), .B(data_in3[56]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[56]) );
  MUX2_X1 md2FF_U56 ( .A(md2FF_permOut[55]), .B(data_in3[55]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[55]) );
  MUX2_X1 md2FF_U55 ( .A(md2FF_permOut[54]), .B(data_in3[54]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[54]) );
  MUX2_X1 md2FF_U54 ( .A(md2FF_permOut[53]), .B(data_in3[53]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[53]) );
  MUX2_X1 md2FF_U53 ( .A(md2FF_permOut[52]), .B(data_in3[52]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[52]) );
  MUX2_X1 md2FF_U52 ( .A(md2FF_permOut[51]), .B(data_in3[51]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[51]) );
  MUX2_X1 md2FF_U51 ( .A(md2FF_permOut[50]), .B(data_in3[50]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[50]) );
  MUX2_X1 md2FF_U50 ( .A(md2FF_permOut[49]), .B(data_in3[49]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[49]) );
  MUX2_X1 md2FF_U49 ( .A(md2FF_permOut[48]), .B(data_in3[48]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[48]) );
  MUX2_X1 md2FF_U48 ( .A(md2FF_permOut[47]), .B(data_in3[47]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[47]) );
  MUX2_X1 md2FF_U47 ( .A(md2FF_permOut[46]), .B(data_in3[46]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[46]) );
  MUX2_X1 md2FF_U46 ( .A(md2FF_permOut[45]), .B(data_in3[45]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[45]) );
  MUX2_X1 md2FF_U45 ( .A(md2FF_permOut[44]), .B(data_in3[44]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[44]) );
  MUX2_X1 md2FF_U44 ( .A(md2FF_permOut[43]), .B(data_in3[43]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[43]) );
  MUX2_X1 md2FF_U43 ( .A(md2FF_permOut[42]), .B(data_in3[42]), .S(md2FF_n265), 
        .Z(md2FF_inputPar[42]) );
  INV_X1 md2FF_U42 ( .A(md2FF_n263), .ZN(md2FF_n265) );
  MUX2_X1 md2FF_U41 ( .A(md2FF_permOut[41]), .B(data_in3[41]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[41]) );
  MUX2_X1 md2FF_U40 ( .A(md2FF_permOut[40]), .B(data_in3[40]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[40]) );
  MUX2_X1 md2FF_U39 ( .A(md2FF_permOut[39]), .B(data_in3[39]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[39]) );
  MUX2_X1 md2FF_U38 ( .A(md2FF_permOut[38]), .B(data_in3[38]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[38]) );
  MUX2_X1 md2FF_U37 ( .A(md2FF_permOut[37]), .B(data_in3[37]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[37]) );
  MUX2_X1 md2FF_U36 ( .A(md2FF_permOut[36]), .B(data_in3[36]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[36]) );
  MUX2_X1 md2FF_U35 ( .A(md2FF_permOut[35]), .B(data_in3[35]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[35]) );
  MUX2_X1 md2FF_U34 ( .A(md2FF_permOut[34]), .B(data_in3[34]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[34]) );
  MUX2_X1 md2FF_U33 ( .A(md2FF_permOut[33]), .B(data_in3[33]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[33]) );
  MUX2_X1 md2FF_U32 ( .A(md2FF_permOut[32]), .B(data_in3[32]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[32]) );
  MUX2_X1 md2FF_U31 ( .A(md2FF_permOut[31]), .B(data_in3[31]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[31]) );
  MUX2_X1 md2FF_U30 ( .A(md2FF_permOut[30]), .B(data_in3[30]), .S(md2FF_n266), 
        .Z(md2FF_inputPar[30]) );
  INV_X1 md2FF_U29 ( .A(md2FF_n263), .ZN(md2FF_n266) );
  MUX2_X1 md2FF_U28 ( .A(md2FF_permOut[29]), .B(data_in3[29]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[29]) );
  MUX2_X1 md2FF_U27 ( .A(md2FF_permOut[28]), .B(data_in3[28]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[28]) );
  MUX2_X1 md2FF_U26 ( .A(md2FF_permOut[27]), .B(data_in3[27]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[27]) );
  MUX2_X1 md2FF_U25 ( .A(md2FF_permOut[26]), .B(data_in3[26]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[26]) );
  MUX2_X1 md2FF_U24 ( .A(md2FF_permOut[25]), .B(data_in3[25]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[25]) );
  MUX2_X1 md2FF_U23 ( .A(md2FF_permOut[24]), .B(data_in3[24]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[24]) );
  MUX2_X1 md2FF_U22 ( .A(md2FF_permOut[23]), .B(data_in3[23]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[23]) );
  MUX2_X1 md2FF_U21 ( .A(md2FF_permOut[22]), .B(data_in3[22]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[22]) );
  MUX2_X1 md2FF_U20 ( .A(md2FF_permOut[21]), .B(data_in3[21]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[21]) );
  MUX2_X1 md2FF_U19 ( .A(md2FF_permOut[20]), .B(data_in3[20]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[20]) );
  MUX2_X1 md2FF_U18 ( .A(md2FF_permOut[19]), .B(data_in3[19]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[19]) );
  MUX2_X1 md2FF_U17 ( .A(md2FF_permOut[18]), .B(data_in3[18]), .S(md2FF_n267), 
        .Z(md2FF_inputPar[18]) );
  INV_X1 md2FF_U16 ( .A(md2FF_n263), .ZN(md2FF_n267) );
  MUX2_X1 md2FF_U15 ( .A(md2FF_permOut[17]), .B(data_in3[17]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[17]) );
  MUX2_X1 md2FF_U14 ( .A(md2FF_permOut[16]), .B(data_in3[16]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[16]) );
  MUX2_X1 md2FF_U13 ( .A(md2FF_permOut[15]), .B(data_in3[15]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[15]) );
  MUX2_X1 md2FF_U12 ( .A(md2FF_permOut[14]), .B(data_in3[14]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[14]) );
  MUX2_X1 md2FF_U11 ( .A(md2FF_permOut[13]), .B(data_in3[13]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[13]) );
  MUX2_X1 md2FF_U10 ( .A(md2FF_permOut[12]), .B(data_in3[12]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[12]) );
  MUX2_X1 md2FF_U9 ( .A(md2FF_permOut[11]), .B(data_in3[11]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[11]) );
  MUX2_X1 md2FF_U8 ( .A(md2FF_permOut[10]), .B(data_in3[10]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[10]) );
  MUX2_X1 md2FF_U7 ( .A(md2FF_permOut[3]), .B(data_in3[3]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[3]) );
  MUX2_X1 md2FF_U6 ( .A(md2FF_permOut[2]), .B(data_in3[2]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[2]) );
  MUX2_X1 md2FF_U5 ( .A(md2FF_permOut[1]), .B(data_in3[1]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[1]) );
  MUX2_X1 md2FF_U4 ( .A(md2FF_permOut[0]), .B(data_in3[0]), .S(md2FF_n264), 
        .Z(md2FF_inputPar[0]) );
  INV_X1 md2FF_U3 ( .A(md2FF_n263), .ZN(md2FF_n264) );
  INV_X1 md2FF_U2 ( .A(ctrlData[2]), .ZN(md2FF_n263) );
  INV_X2 md2FF_state_U5 ( .A(md2FF_state_n11), .ZN(md2FF_state_n10) );
  INV_X2 md2FF_state_U4 ( .A(md2FF_state_n11), .ZN(md2FF_state_n9) );
  INV_X1 md2FF_state_U3 ( .A(ctrlData[0]), .ZN(md2FF_state_n11) );
  INV_X1 md2FF_state_U2 ( .A(md2FF_state_n8), .ZN(md2FF_state_n7) );
  INV_X1 md2FF_state_U1 ( .A(ctrlData[1]), .ZN(md2FF_state_n8) );
  NAND2_X1 md2FF_state_gff_1_U19 ( .A1(md2FF_state_gff_1_n67), .A2(
        md2FF_state_gff_1_n66), .ZN(md2FF_state_gff_1_n30) );
  NAND2_X1 md2FF_state_gff_1_U18 ( .A1(md2FF_state_gff_1_n65), .A2(
        md2FF_permOut[16]), .ZN(md2FF_state_gff_1_n66) );
  MUX2_X1 md2FF_state_gff_1_U17 ( .A(md2FF_state_gff_1_n34), .B(
        md2FF_state_gff_1_n64), .S(md2FF_state_n7), .Z(md2FF_state_gff_1_n67)
         );
  NAND2_X1 md2FF_state_gff_1_U16 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[1]), 
        .ZN(md2FF_state_gff_1_n64) );
  NAND2_X1 md2FF_state_gff_1_U15 ( .A1(md2FF_state_gff_1_n63), .A2(
        md2FF_state_gff_1_n62), .ZN(md2FF_state_gff_1_n28) );
  NAND2_X1 md2FF_state_gff_1_U14 ( .A1(md2FF_state_gff_1_n65), .A2(
        md2FF_permOut[48]), .ZN(md2FF_state_gff_1_n62) );
  MUX2_X1 md2FF_state_gff_1_U13 ( .A(md2FF_state_gff_1_n32), .B(
        md2FF_state_gff_1_n61), .S(md2FF_state_n7), .Z(md2FF_state_gff_1_n63)
         );
  NAND2_X1 md2FF_state_gff_1_U12 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[3]), 
        .ZN(md2FF_state_gff_1_n61) );
  NAND2_X1 md2FF_state_gff_1_U11 ( .A1(md2FF_state_gff_1_n60), .A2(
        md2FF_state_gff_1_n59), .ZN(md2FF_state_gff_1_n31) );
  NAND2_X1 md2FF_state_gff_1_U10 ( .A1(md2FF_state_gff_1_n65), .A2(
        md2FF_permOut[0]), .ZN(md2FF_state_gff_1_n59) );
  MUX2_X1 md2FF_state_gff_1_U9 ( .A(md2FF_state_gff_1_n35), .B(
        md2FF_state_gff_1_n58), .S(md2FF_state_n7), .Z(md2FF_state_gff_1_n60)
         );
  NAND2_X1 md2FF_state_gff_1_U8 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[0]), 
        .ZN(md2FF_state_gff_1_n58) );
  NAND2_X1 md2FF_state_gff_1_U7 ( .A1(md2FF_state_gff_1_n57), .A2(
        md2FF_state_gff_1_n56), .ZN(md2FF_state_gff_1_n29) );
  NAND2_X1 md2FF_state_gff_1_U6 ( .A1(md2FF_state_gff_1_n65), .A2(
        md2FF_permOut[32]), .ZN(md2FF_state_gff_1_n56) );
  NOR2_X1 md2FF_state_gff_1_U5 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_1_n55), .ZN(md2FF_state_gff_1_n65) );
  INV_X1 md2FF_state_gff_1_U4 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_1_n55)
         );
  MUX2_X1 md2FF_state_gff_1_U3 ( .A(md2FF_state_gff_1_n33), .B(
        md2FF_state_gff_1_n54), .S(md2FF_state_n7), .Z(md2FF_state_gff_1_n57)
         );
  NAND2_X1 md2FF_state_gff_1_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[2]), 
        .ZN(md2FF_state_gff_1_n54) );
  DFF_X1 md2FF_state_gff_1_s_current_state_reg_0_ ( .D(md2FF_state_gff_1_n31), 
        .CK(clk), .Q(md2FF_permOut[1]), .QN(md2FF_state_gff_1_n35) );
  DFF_X1 md2FF_state_gff_1_s_current_state_reg_1_ ( .D(md2FF_state_gff_1_n30), 
        .CK(clk), .Q(md2FF_permOut[17]), .QN(md2FF_state_gff_1_n34) );
  DFF_X1 md2FF_state_gff_1_s_current_state_reg_2_ ( .D(md2FF_state_gff_1_n29), 
        .CK(clk), .Q(md2FF_permOut[33]), .QN(md2FF_state_gff_1_n33) );
  DFF_X1 md2FF_state_gff_1_s_current_state_reg_3_ ( .D(md2FF_state_gff_1_n28), 
        .CK(clk), .Q(md2FF_permOut[49]), .QN(md2FF_state_gff_1_n32) );
  NAND2_X1 md2FF_state_gff_2_U20 ( .A1(md2FF_state_gff_2_n68), .A2(
        md2FF_state_gff_2_n67), .ZN(md2FF_state_gff_2_n28) );
  NAND2_X1 md2FF_state_gff_2_U19 ( .A1(md2FF_state_gff_2_n66), .A2(
        md2FF_permOut[49]), .ZN(md2FF_state_gff_2_n67) );
  MUX2_X1 md2FF_state_gff_2_U18 ( .A(md2FF_state_gff_2_n32), .B(
        md2FF_state_gff_2_n65), .S(md2FF_state_gff_2_n64), .Z(
        md2FF_state_gff_2_n68) );
  NAND2_X1 md2FF_state_gff_2_U17 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[7]), 
        .ZN(md2FF_state_gff_2_n65) );
  NAND2_X1 md2FF_state_gff_2_U16 ( .A1(md2FF_state_gff_2_n63), .A2(
        md2FF_state_gff_2_n62), .ZN(md2FF_state_gff_2_n29) );
  NAND2_X1 md2FF_state_gff_2_U15 ( .A1(md2FF_state_gff_2_n66), .A2(
        md2FF_permOut[33]), .ZN(md2FF_state_gff_2_n62) );
  MUX2_X1 md2FF_state_gff_2_U14 ( .A(md2FF_state_gff_2_n33), .B(
        md2FF_state_gff_2_n61), .S(md2FF_state_gff_2_n64), .Z(
        md2FF_state_gff_2_n63) );
  NAND2_X1 md2FF_state_gff_2_U13 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[6]), 
        .ZN(md2FF_state_gff_2_n61) );
  NAND2_X1 md2FF_state_gff_2_U12 ( .A1(md2FF_state_gff_2_n60), .A2(
        md2FF_state_gff_2_n59), .ZN(md2FF_state_gff_2_n30) );
  NAND2_X1 md2FF_state_gff_2_U11 ( .A1(md2FF_state_gff_2_n66), .A2(
        md2FF_permOut[17]), .ZN(md2FF_state_gff_2_n59) );
  MUX2_X1 md2FF_state_gff_2_U10 ( .A(md2FF_state_gff_2_n34), .B(
        md2FF_state_gff_2_n58), .S(md2FF_state_gff_2_n64), .Z(
        md2FF_state_gff_2_n60) );
  NAND2_X1 md2FF_state_gff_2_U9 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[5]), 
        .ZN(md2FF_state_gff_2_n58) );
  NAND2_X1 md2FF_state_gff_2_U8 ( .A1(md2FF_state_gff_2_n57), .A2(
        md2FF_state_gff_2_n56), .ZN(md2FF_state_gff_2_n31) );
  NAND2_X1 md2FF_state_gff_2_U7 ( .A1(md2FF_state_gff_2_n66), .A2(
        md2FF_permOut[1]), .ZN(md2FF_state_gff_2_n56) );
  NOR2_X1 md2FF_state_gff_2_U6 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_2_n55), .ZN(md2FF_state_gff_2_n66) );
  MUX2_X1 md2FF_state_gff_2_U5 ( .A(md2FF_state_gff_2_n35), .B(
        md2FF_state_gff_2_n54), .S(md2FF_state_gff_2_n64), .Z(
        md2FF_state_gff_2_n57) );
  INV_X1 md2FF_state_gff_2_U4 ( .A(md2FF_state_gff_2_n55), .ZN(
        md2FF_state_gff_2_n64) );
  INV_X1 md2FF_state_gff_2_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_2_n55)
         );
  NAND2_X1 md2FF_state_gff_2_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[4]), 
        .ZN(md2FF_state_gff_2_n54) );
  DFF_X1 md2FF_state_gff_2_s_current_state_reg_0_ ( .D(md2FF_state_gff_2_n31), 
        .CK(clk), .Q(md2FF_permOut[2]), .QN(md2FF_state_gff_2_n35) );
  DFF_X1 md2FF_state_gff_2_s_current_state_reg_1_ ( .D(md2FF_state_gff_2_n30), 
        .CK(clk), .Q(md2FF_permOut[18]), .QN(md2FF_state_gff_2_n34) );
  DFF_X1 md2FF_state_gff_2_s_current_state_reg_2_ ( .D(md2FF_state_gff_2_n29), 
        .CK(clk), .Q(md2FF_permOut[34]), .QN(md2FF_state_gff_2_n33) );
  DFF_X1 md2FF_state_gff_2_s_current_state_reg_3_ ( .D(md2FF_state_gff_2_n28), 
        .CK(clk), .Q(md2FF_permOut[50]), .QN(md2FF_state_gff_2_n32) );
  NAND2_X1 md2FF_state_gff_3_U20 ( .A1(md2FF_state_gff_3_n68), .A2(
        md2FF_state_gff_3_n67), .ZN(md2FF_state_gff_3_n30) );
  NAND2_X1 md2FF_state_gff_3_U19 ( .A1(md2FF_state_gff_3_n66), .A2(
        md2FF_permOut[18]), .ZN(md2FF_state_gff_3_n67) );
  MUX2_X1 md2FF_state_gff_3_U18 ( .A(md2FF_state_gff_3_n34), .B(
        md2FF_state_gff_3_n65), .S(md2FF_state_gff_3_n64), .Z(
        md2FF_state_gff_3_n68) );
  NAND2_X1 md2FF_state_gff_3_U17 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[9]), .ZN(md2FF_state_gff_3_n65) );
  NAND2_X1 md2FF_state_gff_3_U16 ( .A1(md2FF_state_gff_3_n63), .A2(
        md2FF_state_gff_3_n62), .ZN(md2FF_state_gff_3_n31) );
  NAND2_X1 md2FF_state_gff_3_U15 ( .A1(md2FF_state_gff_3_n66), .A2(
        md2FF_permOut[2]), .ZN(md2FF_state_gff_3_n62) );
  MUX2_X1 md2FF_state_gff_3_U14 ( .A(md2FF_state_gff_3_n35), .B(
        md2FF_state_gff_3_n61), .S(md2FF_state_gff_3_n64), .Z(
        md2FF_state_gff_3_n63) );
  NAND2_X1 md2FF_state_gff_3_U13 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[8]), .ZN(md2FF_state_gff_3_n61) );
  NAND2_X1 md2FF_state_gff_3_U12 ( .A1(md2FF_state_gff_3_n60), .A2(
        md2FF_state_gff_3_n59), .ZN(md2FF_state_gff_3_n28) );
  NAND2_X1 md2FF_state_gff_3_U11 ( .A1(md2FF_state_gff_3_n66), .A2(
        md2FF_permOut[50]), .ZN(md2FF_state_gff_3_n59) );
  MUX2_X1 md2FF_state_gff_3_U10 ( .A(md2FF_state_gff_3_n32), .B(
        md2FF_state_gff_3_n58), .S(md2FF_state_gff_3_n64), .Z(
        md2FF_state_gff_3_n60) );
  NAND2_X1 md2FF_state_gff_3_U9 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[11]), .ZN(md2FF_state_gff_3_n58) );
  NAND2_X1 md2FF_state_gff_3_U8 ( .A1(md2FF_state_gff_3_n57), .A2(
        md2FF_state_gff_3_n56), .ZN(md2FF_state_gff_3_n29) );
  NAND2_X1 md2FF_state_gff_3_U7 ( .A1(md2FF_state_gff_3_n66), .A2(
        md2FF_permOut[34]), .ZN(md2FF_state_gff_3_n56) );
  NOR2_X1 md2FF_state_gff_3_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_3_n55), .ZN(md2FF_state_gff_3_n66) );
  MUX2_X1 md2FF_state_gff_3_U5 ( .A(md2FF_state_gff_3_n33), .B(
        md2FF_state_gff_3_n54), .S(md2FF_state_gff_3_n64), .Z(
        md2FF_state_gff_3_n57) );
  INV_X1 md2FF_state_gff_3_U4 ( .A(md2FF_state_gff_3_n55), .ZN(
        md2FF_state_gff_3_n64) );
  INV_X1 md2FF_state_gff_3_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_3_n55)
         );
  NAND2_X1 md2FF_state_gff_3_U2 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[10]), .ZN(md2FF_state_gff_3_n54) );
  DFF_X1 md2FF_state_gff_3_s_current_state_reg_0_ ( .D(md2FF_state_gff_3_n31), 
        .CK(clk), .Q(md2FF_permOut[3]), .QN(md2FF_state_gff_3_n35) );
  DFF_X1 md2FF_state_gff_3_s_current_state_reg_1_ ( .D(md2FF_state_gff_3_n30), 
        .CK(clk), .Q(md2FF_permOut[19]), .QN(md2FF_state_gff_3_n34) );
  DFF_X1 md2FF_state_gff_3_s_current_state_reg_2_ ( .D(md2FF_state_gff_3_n29), 
        .CK(clk), .Q(md2FF_permOut[35]), .QN(md2FF_state_gff_3_n33) );
  DFF_X1 md2FF_state_gff_3_s_current_state_reg_3_ ( .D(md2FF_state_gff_3_n28), 
        .CK(clk), .Q(md2FF_permOut[51]), .QN(md2FF_state_gff_3_n32) );
  NAND2_X1 md2FF_state_gff_4_U20 ( .A1(md2FF_state_gff_4_n68), .A2(
        md2FF_state_gff_4_n67), .ZN(md2FF_state_gff_4_n28) );
  NAND2_X1 md2FF_state_gff_4_U19 ( .A1(md2FF_state_gff_4_n66), .A2(
        md2FF_permOut[51]), .ZN(md2FF_state_gff_4_n67) );
  MUX2_X1 md2FF_state_gff_4_U18 ( .A(md2FF_state_gff_4_n32), .B(
        md2FF_state_gff_4_n65), .S(md2FF_state_gff_4_n64), .Z(
        md2FF_state_gff_4_n68) );
  NAND2_X1 md2FF_state_gff_4_U17 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[15]), .ZN(md2FF_state_gff_4_n65) );
  NAND2_X1 md2FF_state_gff_4_U16 ( .A1(md2FF_state_gff_4_n63), .A2(
        md2FF_state_gff_4_n62), .ZN(md2FF_state_gff_4_n29) );
  NAND2_X1 md2FF_state_gff_4_U15 ( .A1(md2FF_state_gff_4_n66), .A2(
        md2FF_permOut[35]), .ZN(md2FF_state_gff_4_n62) );
  MUX2_X1 md2FF_state_gff_4_U14 ( .A(md2FF_state_gff_4_n33), .B(
        md2FF_state_gff_4_n61), .S(md2FF_state_gff_4_n64), .Z(
        md2FF_state_gff_4_n63) );
  NAND2_X1 md2FF_state_gff_4_U13 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[14]), .ZN(md2FF_state_gff_4_n61) );
  NAND2_X1 md2FF_state_gff_4_U12 ( .A1(md2FF_state_gff_4_n60), .A2(
        md2FF_state_gff_4_n59), .ZN(md2FF_state_gff_4_n30) );
  NAND2_X1 md2FF_state_gff_4_U11 ( .A1(md2FF_state_gff_4_n66), .A2(
        md2FF_permOut[19]), .ZN(md2FF_state_gff_4_n59) );
  MUX2_X1 md2FF_state_gff_4_U10 ( .A(md2FF_state_gff_4_n34), .B(
        md2FF_state_gff_4_n58), .S(md2FF_state_gff_4_n64), .Z(
        md2FF_state_gff_4_n60) );
  NAND2_X1 md2FF_state_gff_4_U9 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[13]), 
        .ZN(md2FF_state_gff_4_n58) );
  NAND2_X1 md2FF_state_gff_4_U8 ( .A1(md2FF_state_gff_4_n57), .A2(
        md2FF_state_gff_4_n56), .ZN(md2FF_state_gff_4_n31) );
  NAND2_X1 md2FF_state_gff_4_U7 ( .A1(md2FF_state_gff_4_n66), .A2(
        md2FF_permOut[3]), .ZN(md2FF_state_gff_4_n56) );
  NOR2_X1 md2FF_state_gff_4_U6 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_4_n55), .ZN(md2FF_state_gff_4_n66) );
  MUX2_X1 md2FF_state_gff_4_U5 ( .A(md2FF_state_gff_4_n35), .B(
        md2FF_state_gff_4_n54), .S(md2FF_state_gff_4_n64), .Z(
        md2FF_state_gff_4_n57) );
  INV_X1 md2FF_state_gff_4_U4 ( .A(md2FF_state_gff_4_n55), .ZN(
        md2FF_state_gff_4_n64) );
  INV_X1 md2FF_state_gff_4_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_4_n55)
         );
  NAND2_X1 md2FF_state_gff_4_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[12]), 
        .ZN(md2FF_state_gff_4_n54) );
  DFF_X1 md2FF_state_gff_4_s_current_state_reg_0_ ( .D(md2FF_state_gff_4_n31), 
        .CK(clk), .Q(md2FF_permOut[4]), .QN(md2FF_state_gff_4_n35) );
  DFF_X1 md2FF_state_gff_4_s_current_state_reg_1_ ( .D(md2FF_state_gff_4_n30), 
        .CK(clk), .Q(md2FF_permOut[20]), .QN(md2FF_state_gff_4_n34) );
  DFF_X1 md2FF_state_gff_4_s_current_state_reg_2_ ( .D(md2FF_state_gff_4_n29), 
        .CK(clk), .Q(md2FF_permOut[36]), .QN(md2FF_state_gff_4_n33) );
  DFF_X1 md2FF_state_gff_4_s_current_state_reg_3_ ( .D(md2FF_state_gff_4_n28), 
        .CK(clk), .Q(md2FF_permOut[52]), .QN(md2FF_state_gff_4_n32) );
  NAND2_X1 md2FF_state_gff_5_U20 ( .A1(md2FF_state_gff_5_n69), .A2(
        md2FF_state_gff_5_n68), .ZN(md2FF_state_gff_5_n29) );
  NAND2_X1 md2FF_state_gff_5_U19 ( .A1(md2FF_state_gff_5_n67), .A2(
        md2FF_permOut[52]), .ZN(md2FF_state_gff_5_n68) );
  MUX2_X1 md2FF_state_gff_5_U18 ( .A(md2FF_state_gff_5_n33), .B(
        md2FF_state_gff_5_n66), .S(md2FF_state_gff_5_n65), .Z(
        md2FF_state_gff_5_n69) );
  NAND2_X1 md2FF_state_gff_5_U17 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[19]), .ZN(md2FF_state_gff_5_n66) );
  NAND2_X1 md2FF_state_gff_5_U16 ( .A1(md2FF_state_gff_5_n64), .A2(
        md2FF_state_gff_5_n63), .ZN(md2FF_state_gff_5_n30) );
  NAND2_X1 md2FF_state_gff_5_U15 ( .A1(md2FF_state_gff_5_n67), .A2(
        md2FF_permOut[36]), .ZN(md2FF_state_gff_5_n63) );
  MUX2_X1 md2FF_state_gff_5_U14 ( .A(md2FF_state_gff_5_n34), .B(
        md2FF_state_gff_5_n62), .S(md2FF_state_gff_5_n65), .Z(
        md2FF_state_gff_5_n64) );
  NAND2_X1 md2FF_state_gff_5_U13 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[18]), .ZN(md2FF_state_gff_5_n62) );
  NAND2_X1 md2FF_state_gff_5_U12 ( .A1(md2FF_state_gff_5_n61), .A2(
        md2FF_state_gff_5_n60), .ZN(md2FF_state_gff_5_n31) );
  NAND2_X1 md2FF_state_gff_5_U11 ( .A1(md2FF_state_gff_5_n67), .A2(
        md2FF_permOut[20]), .ZN(md2FF_state_gff_5_n60) );
  MUX2_X1 md2FF_state_gff_5_U10 ( .A(md2FF_state_gff_5_n35), .B(
        md2FF_state_gff_5_n59), .S(md2FF_state_gff_5_n65), .Z(
        md2FF_state_gff_5_n61) );
  NAND2_X1 md2FF_state_gff_5_U9 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[17]), 
        .ZN(md2FF_state_gff_5_n59) );
  NAND2_X1 md2FF_state_gff_5_U8 ( .A1(md2FF_state_gff_5_n58), .A2(
        md2FF_state_gff_5_n57), .ZN(md2FF_state_gff_5_n32) );
  NAND2_X1 md2FF_state_gff_5_U7 ( .A1(md2FF_state_gff_5_n67), .A2(
        md2FF_permOut[4]), .ZN(md2FF_state_gff_5_n57) );
  NOR2_X1 md2FF_state_gff_5_U6 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_5_n56), .ZN(md2FF_state_gff_5_n67) );
  MUX2_X1 md2FF_state_gff_5_U5 ( .A(md2FF_state_gff_5_n36), .B(
        md2FF_state_gff_5_n55), .S(md2FF_state_gff_5_n65), .Z(
        md2FF_state_gff_5_n58) );
  INV_X1 md2FF_state_gff_5_U4 ( .A(md2FF_state_gff_5_n56), .ZN(
        md2FF_state_gff_5_n65) );
  INV_X1 md2FF_state_gff_5_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_5_n56)
         );
  NAND2_X1 md2FF_state_gff_5_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[16]), 
        .ZN(md2FF_state_gff_5_n55) );
  DFF_X1 md2FF_state_gff_5_s_current_state_reg_0_ ( .D(md2FF_state_gff_5_n32), 
        .CK(clk), .Q(md2FF_permOut[5]), .QN(md2FF_state_gff_5_n36) );
  DFF_X1 md2FF_state_gff_5_s_current_state_reg_1_ ( .D(md2FF_state_gff_5_n31), 
        .CK(clk), .Q(md2FF_permOut[21]), .QN(md2FF_state_gff_5_n35) );
  DFF_X1 md2FF_state_gff_5_s_current_state_reg_2_ ( .D(md2FF_state_gff_5_n30), 
        .CK(clk), .Q(md2FF_permOut[37]), .QN(md2FF_state_gff_5_n34) );
  DFF_X1 md2FF_state_gff_5_s_current_state_reg_3_ ( .D(md2FF_state_gff_5_n29), 
        .CK(clk), .Q(md2FF_permOut[53]), .QN(md2FF_state_gff_5_n33) );
  NAND2_X1 md2FF_state_gff_6_U20 ( .A1(md2FF_state_gff_6_n69), .A2(
        md2FF_state_gff_6_n68), .ZN(md2FF_state_gff_6_n29) );
  NAND2_X1 md2FF_state_gff_6_U19 ( .A1(md2FF_state_gff_6_n67), .A2(
        md2FF_permOut[53]), .ZN(md2FF_state_gff_6_n68) );
  MUX2_X1 md2FF_state_gff_6_U18 ( .A(md2FF_state_gff_6_n33), .B(
        md2FF_state_gff_6_n66), .S(md2FF_state_gff_6_n65), .Z(
        md2FF_state_gff_6_n69) );
  NAND2_X1 md2FF_state_gff_6_U17 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[23]), .ZN(md2FF_state_gff_6_n66) );
  NAND2_X1 md2FF_state_gff_6_U16 ( .A1(md2FF_state_gff_6_n64), .A2(
        md2FF_state_gff_6_n63), .ZN(md2FF_state_gff_6_n30) );
  NAND2_X1 md2FF_state_gff_6_U15 ( .A1(md2FF_state_gff_6_n67), .A2(
        md2FF_permOut[37]), .ZN(md2FF_state_gff_6_n63) );
  MUX2_X1 md2FF_state_gff_6_U14 ( .A(md2FF_state_gff_6_n34), .B(
        md2FF_state_gff_6_n62), .S(md2FF_state_gff_6_n65), .Z(
        md2FF_state_gff_6_n64) );
  NAND2_X1 md2FF_state_gff_6_U13 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[22]), .ZN(md2FF_state_gff_6_n62) );
  NAND2_X1 md2FF_state_gff_6_U12 ( .A1(md2FF_state_gff_6_n61), .A2(
        md2FF_state_gff_6_n60), .ZN(md2FF_state_gff_6_n31) );
  NAND2_X1 md2FF_state_gff_6_U11 ( .A1(md2FF_state_gff_6_n67), .A2(
        md2FF_permOut[21]), .ZN(md2FF_state_gff_6_n60) );
  MUX2_X1 md2FF_state_gff_6_U10 ( .A(md2FF_state_gff_6_n35), .B(
        md2FF_state_gff_6_n59), .S(md2FF_state_gff_6_n65), .Z(
        md2FF_state_gff_6_n61) );
  NAND2_X1 md2FF_state_gff_6_U9 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[21]), .ZN(md2FF_state_gff_6_n59) );
  NAND2_X1 md2FF_state_gff_6_U8 ( .A1(md2FF_state_gff_6_n58), .A2(
        md2FF_state_gff_6_n57), .ZN(md2FF_state_gff_6_n32) );
  NAND2_X1 md2FF_state_gff_6_U7 ( .A1(md2FF_state_gff_6_n67), .A2(
        md2FF_permOut[5]), .ZN(md2FF_state_gff_6_n57) );
  NOR2_X1 md2FF_state_gff_6_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_6_n56), .ZN(md2FF_state_gff_6_n67) );
  MUX2_X1 md2FF_state_gff_6_U5 ( .A(md2FF_state_gff_6_n36), .B(
        md2FF_state_gff_6_n55), .S(md2FF_state_gff_6_n65), .Z(
        md2FF_state_gff_6_n58) );
  INV_X1 md2FF_state_gff_6_U4 ( .A(md2FF_state_gff_6_n56), .ZN(
        md2FF_state_gff_6_n65) );
  INV_X1 md2FF_state_gff_6_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_6_n56)
         );
  NAND2_X1 md2FF_state_gff_6_U2 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[20]), .ZN(md2FF_state_gff_6_n55) );
  DFF_X1 md2FF_state_gff_6_s_current_state_reg_0_ ( .D(md2FF_state_gff_6_n32), 
        .CK(clk), .Q(md2FF_permOut[6]), .QN(md2FF_state_gff_6_n36) );
  DFF_X1 md2FF_state_gff_6_s_current_state_reg_1_ ( .D(md2FF_state_gff_6_n31), 
        .CK(clk), .Q(md2FF_permOut[22]), .QN(md2FF_state_gff_6_n35) );
  DFF_X1 md2FF_state_gff_6_s_current_state_reg_2_ ( .D(md2FF_state_gff_6_n30), 
        .CK(clk), .Q(md2FF_permOut[38]), .QN(md2FF_state_gff_6_n34) );
  DFF_X1 md2FF_state_gff_6_s_current_state_reg_3_ ( .D(md2FF_state_gff_6_n29), 
        .CK(clk), .Q(md2FF_permOut[54]), .QN(md2FF_state_gff_6_n33) );
  NAND2_X1 md2FF_state_gff_7_U20 ( .A1(md2FF_state_gff_7_n69), .A2(
        md2FF_state_gff_7_n68), .ZN(md2FF_state_gff_7_n29) );
  NAND2_X1 md2FF_state_gff_7_U19 ( .A1(md2FF_state_gff_7_n67), .A2(
        md2FF_permOut[54]), .ZN(md2FF_state_gff_7_n68) );
  MUX2_X1 md2FF_state_gff_7_U18 ( .A(md2FF_state_gff_7_n33), .B(
        md2FF_state_gff_7_n66), .S(md2FF_state_gff_7_n65), .Z(
        md2FF_state_gff_7_n69) );
  NAND2_X1 md2FF_state_gff_7_U17 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[27]), .ZN(md2FF_state_gff_7_n66) );
  NAND2_X1 md2FF_state_gff_7_U16 ( .A1(md2FF_state_gff_7_n64), .A2(
        md2FF_state_gff_7_n63), .ZN(md2FF_state_gff_7_n30) );
  NAND2_X1 md2FF_state_gff_7_U15 ( .A1(md2FF_state_gff_7_n67), .A2(
        md2FF_permOut[38]), .ZN(md2FF_state_gff_7_n63) );
  MUX2_X1 md2FF_state_gff_7_U14 ( .A(md2FF_state_gff_7_n34), .B(
        md2FF_state_gff_7_n62), .S(md2FF_state_gff_7_n65), .Z(
        md2FF_state_gff_7_n64) );
  NAND2_X1 md2FF_state_gff_7_U13 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[26]), .ZN(md2FF_state_gff_7_n62) );
  NAND2_X1 md2FF_state_gff_7_U12 ( .A1(md2FF_state_gff_7_n61), .A2(
        md2FF_state_gff_7_n60), .ZN(md2FF_state_gff_7_n31) );
  NAND2_X1 md2FF_state_gff_7_U11 ( .A1(md2FF_state_gff_7_n67), .A2(
        md2FF_permOut[22]), .ZN(md2FF_state_gff_7_n60) );
  MUX2_X1 md2FF_state_gff_7_U10 ( .A(md2FF_state_gff_7_n35), .B(
        md2FF_state_gff_7_n59), .S(md2FF_state_gff_7_n65), .Z(
        md2FF_state_gff_7_n61) );
  NAND2_X1 md2FF_state_gff_7_U9 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[25]), 
        .ZN(md2FF_state_gff_7_n59) );
  NAND2_X1 md2FF_state_gff_7_U8 ( .A1(md2FF_state_gff_7_n58), .A2(
        md2FF_state_gff_7_n57), .ZN(md2FF_state_gff_7_n32) );
  NAND2_X1 md2FF_state_gff_7_U7 ( .A1(md2FF_state_gff_7_n67), .A2(
        md2FF_permOut[6]), .ZN(md2FF_state_gff_7_n57) );
  NOR2_X1 md2FF_state_gff_7_U6 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_7_n56), .ZN(md2FF_state_gff_7_n67) );
  MUX2_X1 md2FF_state_gff_7_U5 ( .A(md2FF_state_gff_7_n36), .B(
        md2FF_state_gff_7_n55), .S(md2FF_state_gff_7_n65), .Z(
        md2FF_state_gff_7_n58) );
  INV_X1 md2FF_state_gff_7_U4 ( .A(md2FF_state_gff_7_n56), .ZN(
        md2FF_state_gff_7_n65) );
  INV_X1 md2FF_state_gff_7_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_7_n56)
         );
  NAND2_X1 md2FF_state_gff_7_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[24]), 
        .ZN(md2FF_state_gff_7_n55) );
  DFF_X1 md2FF_state_gff_7_s_current_state_reg_0_ ( .D(md2FF_state_gff_7_n32), 
        .CK(clk), .Q(md2FF_permOut[7]), .QN(md2FF_state_gff_7_n36) );
  DFF_X1 md2FF_state_gff_7_s_current_state_reg_1_ ( .D(md2FF_state_gff_7_n31), 
        .CK(clk), .Q(md2FF_permOut[23]), .QN(md2FF_state_gff_7_n35) );
  DFF_X1 md2FF_state_gff_7_s_current_state_reg_2_ ( .D(md2FF_state_gff_7_n30), 
        .CK(clk), .Q(md2FF_permOut[39]), .QN(md2FF_state_gff_7_n34) );
  DFF_X1 md2FF_state_gff_7_s_current_state_reg_3_ ( .D(md2FF_state_gff_7_n29), 
        .CK(clk), .Q(md2FF_permOut[55]), .QN(md2FF_state_gff_7_n33) );
  NAND2_X1 md2FF_state_gff_8_U20 ( .A1(md2FF_state_gff_8_n69), .A2(
        md2FF_state_gff_8_n68), .ZN(md2FF_state_gff_8_n29) );
  NAND2_X1 md2FF_state_gff_8_U19 ( .A1(md2FF_state_gff_8_n67), .A2(
        md2FF_permOut[55]), .ZN(md2FF_state_gff_8_n68) );
  MUX2_X1 md2FF_state_gff_8_U18 ( .A(md2FF_state_gff_8_n33), .B(
        md2FF_state_gff_8_n66), .S(md2FF_state_gff_8_n65), .Z(
        md2FF_state_gff_8_n69) );
  NAND2_X1 md2FF_state_gff_8_U17 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[31]), .ZN(md2FF_state_gff_8_n66) );
  NAND2_X1 md2FF_state_gff_8_U16 ( .A1(md2FF_state_gff_8_n64), .A2(
        md2FF_state_gff_8_n63), .ZN(md2FF_state_gff_8_n30) );
  NAND2_X1 md2FF_state_gff_8_U15 ( .A1(md2FF_state_gff_8_n67), .A2(
        md2FF_permOut[39]), .ZN(md2FF_state_gff_8_n63) );
  MUX2_X1 md2FF_state_gff_8_U14 ( .A(md2FF_state_gff_8_n34), .B(
        md2FF_state_gff_8_n62), .S(md2FF_state_gff_8_n65), .Z(
        md2FF_state_gff_8_n64) );
  NAND2_X1 md2FF_state_gff_8_U13 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[30]), .ZN(md2FF_state_gff_8_n62) );
  NAND2_X1 md2FF_state_gff_8_U12 ( .A1(md2FF_state_gff_8_n61), .A2(
        md2FF_state_gff_8_n60), .ZN(md2FF_state_gff_8_n31) );
  NAND2_X1 md2FF_state_gff_8_U11 ( .A1(md2FF_state_gff_8_n67), .A2(
        md2FF_permOut[23]), .ZN(md2FF_state_gff_8_n60) );
  MUX2_X1 md2FF_state_gff_8_U10 ( .A(md2FF_state_gff_8_n35), .B(
        md2FF_state_gff_8_n59), .S(md2FF_state_gff_8_n65), .Z(
        md2FF_state_gff_8_n61) );
  NAND2_X1 md2FF_state_gff_8_U9 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[29]), .ZN(md2FF_state_gff_8_n59) );
  NAND2_X1 md2FF_state_gff_8_U8 ( .A1(md2FF_state_gff_8_n58), .A2(
        md2FF_state_gff_8_n57), .ZN(md2FF_state_gff_8_n32) );
  NAND2_X1 md2FF_state_gff_8_U7 ( .A1(md2FF_state_gff_8_n67), .A2(
        md2FF_permOut[7]), .ZN(md2FF_state_gff_8_n57) );
  NOR2_X1 md2FF_state_gff_8_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_8_n56), .ZN(md2FF_state_gff_8_n67) );
  MUX2_X1 md2FF_state_gff_8_U5 ( .A(md2FF_state_gff_8_n36), .B(
        md2FF_state_gff_8_n55), .S(md2FF_state_gff_8_n65), .Z(
        md2FF_state_gff_8_n58) );
  INV_X1 md2FF_state_gff_8_U4 ( .A(md2FF_state_gff_8_n56), .ZN(
        md2FF_state_gff_8_n65) );
  INV_X1 md2FF_state_gff_8_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_8_n56)
         );
  NAND2_X1 md2FF_state_gff_8_U2 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[28]), .ZN(md2FF_state_gff_8_n55) );
  DFF_X1 md2FF_state_gff_8_s_current_state_reg_0_ ( .D(md2FF_state_gff_8_n32), 
        .CK(clk), .Q(md2FF_permOut[8]), .QN(md2FF_state_gff_8_n36) );
  DFF_X1 md2FF_state_gff_8_s_current_state_reg_1_ ( .D(md2FF_state_gff_8_n31), 
        .CK(clk), .Q(md2FF_permOut[24]), .QN(md2FF_state_gff_8_n35) );
  DFF_X1 md2FF_state_gff_8_s_current_state_reg_2_ ( .D(md2FF_state_gff_8_n30), 
        .CK(clk), .Q(md2FF_permOut[40]), .QN(md2FF_state_gff_8_n34) );
  DFF_X1 md2FF_state_gff_8_s_current_state_reg_3_ ( .D(md2FF_state_gff_8_n29), 
        .CK(clk), .Q(md2FF_permOut[56]), .QN(md2FF_state_gff_8_n33) );
  NAND2_X1 md2FF_state_gff_9_U20 ( .A1(md2FF_state_gff_9_n69), .A2(
        md2FF_state_gff_9_n68), .ZN(md2FF_state_gff_9_n29) );
  NAND2_X1 md2FF_state_gff_9_U19 ( .A1(md2FF_state_gff_9_n67), .A2(
        md2FF_permOut[56]), .ZN(md2FF_state_gff_9_n68) );
  MUX2_X1 md2FF_state_gff_9_U18 ( .A(md2FF_state_gff_9_n33), .B(
        md2FF_state_gff_9_n66), .S(md2FF_state_gff_9_n65), .Z(
        md2FF_state_gff_9_n69) );
  NAND2_X1 md2FF_state_gff_9_U17 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[35]), .ZN(md2FF_state_gff_9_n66) );
  NAND2_X1 md2FF_state_gff_9_U16 ( .A1(md2FF_state_gff_9_n64), .A2(
        md2FF_state_gff_9_n63), .ZN(md2FF_state_gff_9_n30) );
  NAND2_X1 md2FF_state_gff_9_U15 ( .A1(md2FF_state_gff_9_n67), .A2(
        md2FF_permOut[40]), .ZN(md2FF_state_gff_9_n63) );
  MUX2_X1 md2FF_state_gff_9_U14 ( .A(md2FF_state_gff_9_n34), .B(
        md2FF_state_gff_9_n62), .S(md2FF_state_gff_9_n65), .Z(
        md2FF_state_gff_9_n64) );
  NAND2_X1 md2FF_state_gff_9_U13 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[34]), .ZN(md2FF_state_gff_9_n62) );
  NAND2_X1 md2FF_state_gff_9_U12 ( .A1(md2FF_state_gff_9_n61), .A2(
        md2FF_state_gff_9_n60), .ZN(md2FF_state_gff_9_n31) );
  NAND2_X1 md2FF_state_gff_9_U11 ( .A1(md2FF_state_gff_9_n67), .A2(
        md2FF_permOut[24]), .ZN(md2FF_state_gff_9_n60) );
  MUX2_X1 md2FF_state_gff_9_U10 ( .A(md2FF_state_gff_9_n35), .B(
        md2FF_state_gff_9_n59), .S(md2FF_state_gff_9_n65), .Z(
        md2FF_state_gff_9_n61) );
  NAND2_X1 md2FF_state_gff_9_U9 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[33]), .ZN(md2FF_state_gff_9_n59) );
  NAND2_X1 md2FF_state_gff_9_U8 ( .A1(md2FF_state_gff_9_n58), .A2(
        md2FF_state_gff_9_n57), .ZN(md2FF_state_gff_9_n32) );
  NAND2_X1 md2FF_state_gff_9_U7 ( .A1(md2FF_state_gff_9_n67), .A2(
        md2FF_permOut[8]), .ZN(md2FF_state_gff_9_n57) );
  NOR2_X1 md2FF_state_gff_9_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_9_n56), .ZN(md2FF_state_gff_9_n67) );
  MUX2_X1 md2FF_state_gff_9_U5 ( .A(md2FF_state_gff_9_n36), .B(
        md2FF_state_gff_9_n55), .S(md2FF_state_gff_9_n65), .Z(
        md2FF_state_gff_9_n58) );
  INV_X1 md2FF_state_gff_9_U4 ( .A(md2FF_state_gff_9_n56), .ZN(
        md2FF_state_gff_9_n65) );
  INV_X1 md2FF_state_gff_9_U3 ( .A(md2FF_state_n7), .ZN(md2FF_state_gff_9_n56)
         );
  NAND2_X1 md2FF_state_gff_9_U2 ( .A1(md2FF_state_n10), .A2(md2FF_inputPar[32]), .ZN(md2FF_state_gff_9_n55) );
  DFF_X1 md2FF_state_gff_9_s_current_state_reg_0_ ( .D(md2FF_state_gff_9_n32), 
        .CK(clk), .Q(md2FF_permOut[9]), .QN(md2FF_state_gff_9_n36) );
  DFF_X1 md2FF_state_gff_9_s_current_state_reg_1_ ( .D(md2FF_state_gff_9_n31), 
        .CK(clk), .Q(md2FF_permOut[25]), .QN(md2FF_state_gff_9_n35) );
  DFF_X1 md2FF_state_gff_9_s_current_state_reg_2_ ( .D(md2FF_state_gff_9_n30), 
        .CK(clk), .Q(md2FF_permOut[41]), .QN(md2FF_state_gff_9_n34) );
  DFF_X1 md2FF_state_gff_9_s_current_state_reg_3_ ( .D(md2FF_state_gff_9_n29), 
        .CK(clk), .Q(md2FF_permOut[57]), .QN(md2FF_state_gff_9_n33) );
  NAND2_X1 md2FF_state_gff_10_U20 ( .A1(md2FF_state_gff_10_n69), .A2(
        md2FF_state_gff_10_n68), .ZN(md2FF_state_gff_10_n29) );
  NAND2_X1 md2FF_state_gff_10_U19 ( .A1(md2FF_state_gff_10_n67), .A2(
        md2FF_permOut[57]), .ZN(md2FF_state_gff_10_n68) );
  MUX2_X1 md2FF_state_gff_10_U18 ( .A(md2FF_state_gff_10_n33), .B(
        md2FF_state_gff_10_n66), .S(md2FF_state_gff_10_n65), .Z(
        md2FF_state_gff_10_n69) );
  NAND2_X1 md2FF_state_gff_10_U17 ( .A1(md2FF_state_n9), .A2(
        md2FF_inputPar[39]), .ZN(md2FF_state_gff_10_n66) );
  NAND2_X1 md2FF_state_gff_10_U16 ( .A1(md2FF_state_gff_10_n64), .A2(
        md2FF_state_gff_10_n63), .ZN(md2FF_state_gff_10_n30) );
  NAND2_X1 md2FF_state_gff_10_U15 ( .A1(md2FF_state_gff_10_n67), .A2(
        md2FF_permOut[41]), .ZN(md2FF_state_gff_10_n63) );
  MUX2_X1 md2FF_state_gff_10_U14 ( .A(md2FF_state_gff_10_n34), .B(
        md2FF_state_gff_10_n62), .S(md2FF_state_gff_10_n65), .Z(
        md2FF_state_gff_10_n64) );
  NAND2_X1 md2FF_state_gff_10_U13 ( .A1(md2FF_state_n9), .A2(
        md2FF_inputPar[38]), .ZN(md2FF_state_gff_10_n62) );
  NAND2_X1 md2FF_state_gff_10_U12 ( .A1(md2FF_state_gff_10_n61), .A2(
        md2FF_state_gff_10_n60), .ZN(md2FF_state_gff_10_n31) );
  NAND2_X1 md2FF_state_gff_10_U11 ( .A1(md2FF_state_gff_10_n67), .A2(
        md2FF_permOut[25]), .ZN(md2FF_state_gff_10_n60) );
  MUX2_X1 md2FF_state_gff_10_U10 ( .A(md2FF_state_gff_10_n35), .B(
        md2FF_state_gff_10_n59), .S(md2FF_state_gff_10_n65), .Z(
        md2FF_state_gff_10_n61) );
  NAND2_X1 md2FF_state_gff_10_U9 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[37]), .ZN(md2FF_state_gff_10_n59) );
  NAND2_X1 md2FF_state_gff_10_U8 ( .A1(md2FF_state_gff_10_n58), .A2(
        md2FF_state_gff_10_n57), .ZN(md2FF_state_gff_10_n32) );
  NAND2_X1 md2FF_state_gff_10_U7 ( .A1(md2FF_state_gff_10_n67), .A2(
        md2FF_permOut[9]), .ZN(md2FF_state_gff_10_n57) );
  NOR2_X1 md2FF_state_gff_10_U6 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_10_n56), .ZN(md2FF_state_gff_10_n67) );
  MUX2_X1 md2FF_state_gff_10_U5 ( .A(md2FF_state_gff_10_n36), .B(
        md2FF_state_gff_10_n55), .S(md2FF_state_gff_10_n65), .Z(
        md2FF_state_gff_10_n58) );
  INV_X1 md2FF_state_gff_10_U4 ( .A(md2FF_state_gff_10_n56), .ZN(
        md2FF_state_gff_10_n65) );
  INV_X1 md2FF_state_gff_10_U3 ( .A(md2FF_state_n7), .ZN(
        md2FF_state_gff_10_n56) );
  NAND2_X1 md2FF_state_gff_10_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[36]), .ZN(md2FF_state_gff_10_n55) );
DFF_X1 md2FF_state_gff_10_s_current_state_reg_0_ ( .D(md2FF_state_gff_10_n32), .CK(clk), .Q(md2FF_permOut[10]), .QN(md2FF_state_gff_10_n36) );
DFF_X1 md2FF_state_gff_10_s_current_state_reg_1_ ( .D(md2FF_state_gff_10_n31), .CK(clk), .Q(md2FF_permOut[26]), .QN(md2FF_state_gff_10_n35) );
DFF_X1 md2FF_state_gff_10_s_current_state_reg_2_ ( .D(md2FF_state_gff_10_n30), .CK(clk), .Q(md2FF_permOut[42]), .QN(md2FF_state_gff_10_n34) );
DFF_X1 md2FF_state_gff_10_s_current_state_reg_3_ ( .D(md2FF_state_gff_10_n29), .CK(clk), .Q(md2FF_permOut[58]), .QN(md2FF_state_gff_10_n33) );
  NAND2_X1 md2FF_state_gff_11_U20 ( .A1(md2FF_state_gff_11_n69), .A2(
        md2FF_state_gff_11_n68), .ZN(md2FF_state_gff_11_n29) );
  NAND2_X1 md2FF_state_gff_11_U19 ( .A1(md2FF_state_gff_11_n67), .A2(
        md2FF_permOut[58]), .ZN(md2FF_state_gff_11_n68) );
  MUX2_X1 md2FF_state_gff_11_U18 ( .A(md2FF_state_gff_11_n33), .B(
        md2FF_state_gff_11_n66), .S(md2FF_state_gff_11_n65), .Z(
        md2FF_state_gff_11_n69) );
  NAND2_X1 md2FF_state_gff_11_U17 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[43]), .ZN(md2FF_state_gff_11_n66) );
  NAND2_X1 md2FF_state_gff_11_U16 ( .A1(md2FF_state_gff_11_n64), .A2(
        md2FF_state_gff_11_n63), .ZN(md2FF_state_gff_11_n30) );
  NAND2_X1 md2FF_state_gff_11_U15 ( .A1(md2FF_state_gff_11_n67), .A2(
        md2FF_permOut[42]), .ZN(md2FF_state_gff_11_n63) );
  MUX2_X1 md2FF_state_gff_11_U14 ( .A(md2FF_state_gff_11_n34), .B(
        md2FF_state_gff_11_n62), .S(md2FF_state_gff_11_n65), .Z(
        md2FF_state_gff_11_n64) );
  NAND2_X1 md2FF_state_gff_11_U13 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[42]), .ZN(md2FF_state_gff_11_n62) );
  NAND2_X1 md2FF_state_gff_11_U12 ( .A1(md2FF_state_gff_11_n61), .A2(
        md2FF_state_gff_11_n60), .ZN(md2FF_state_gff_11_n31) );
  NAND2_X1 md2FF_state_gff_11_U11 ( .A1(md2FF_state_gff_11_n67), .A2(
        md2FF_permOut[26]), .ZN(md2FF_state_gff_11_n60) );
  MUX2_X1 md2FF_state_gff_11_U10 ( .A(md2FF_state_gff_11_n35), .B(
        md2FF_state_gff_11_n59), .S(md2FF_state_gff_11_n65), .Z(
        md2FF_state_gff_11_n61) );
  NAND2_X1 md2FF_state_gff_11_U9 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[41]), .ZN(md2FF_state_gff_11_n59) );
  NAND2_X1 md2FF_state_gff_11_U8 ( .A1(md2FF_state_gff_11_n58), .A2(
        md2FF_state_gff_11_n57), .ZN(md2FF_state_gff_11_n32) );
  NAND2_X1 md2FF_state_gff_11_U7 ( .A1(md2FF_state_gff_11_n67), .A2(
        md2FF_permOut[10]), .ZN(md2FF_state_gff_11_n57) );
  NOR2_X1 md2FF_state_gff_11_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_11_n56), .ZN(md2FF_state_gff_11_n67) );
  MUX2_X1 md2FF_state_gff_11_U5 ( .A(md2FF_state_gff_11_n36), .B(
        md2FF_state_gff_11_n55), .S(md2FF_state_gff_11_n65), .Z(
        md2FF_state_gff_11_n58) );
  INV_X1 md2FF_state_gff_11_U4 ( .A(md2FF_state_gff_11_n56), .ZN(
        md2FF_state_gff_11_n65) );
  INV_X1 md2FF_state_gff_11_U3 ( .A(md2FF_state_n7), .ZN(
        md2FF_state_gff_11_n56) );
  NAND2_X1 md2FF_state_gff_11_U2 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[40]), .ZN(md2FF_state_gff_11_n55) );
DFF_X1 md2FF_state_gff_11_s_current_state_reg_0_ ( .D(md2FF_state_gff_11_n32), .CK(clk), .Q(md2FF_permOut[11]), .QN(md2FF_state_gff_11_n36) );
DFF_X1 md2FF_state_gff_11_s_current_state_reg_1_ ( .D(md2FF_state_gff_11_n31), .CK(clk), .Q(md2FF_permOut[27]), .QN(md2FF_state_gff_11_n35) );
DFF_X1 md2FF_state_gff_11_s_current_state_reg_2_ ( .D(md2FF_state_gff_11_n30), .CK(clk), .Q(md2FF_permOut[43]), .QN(md2FF_state_gff_11_n34) );
DFF_X1 md2FF_state_gff_11_s_current_state_reg_3_ ( .D(md2FF_state_gff_11_n29), .CK(clk), .Q(md2FF_permOut[59]), .QN(md2FF_state_gff_11_n33) );
  NAND2_X1 md2FF_state_gff_12_U20 ( .A1(md2FF_state_gff_12_n69), .A2(
        md2FF_state_gff_12_n68), .ZN(md2FF_state_gff_12_n29) );
  NAND2_X1 md2FF_state_gff_12_U19 ( .A1(md2FF_state_gff_12_n67), .A2(
        md2FF_permOut[59]), .ZN(md2FF_state_gff_12_n68) );
  MUX2_X1 md2FF_state_gff_12_U18 ( .A(md2FF_state_gff_12_n33), .B(
        md2FF_state_gff_12_n66), .S(md2FF_state_gff_12_n65), .Z(
        md2FF_state_gff_12_n69) );
  NAND2_X1 md2FF_state_gff_12_U17 ( .A1(md2FF_state_n9), .A2(
        md2FF_inputPar[47]), .ZN(md2FF_state_gff_12_n66) );
  NAND2_X1 md2FF_state_gff_12_U16 ( .A1(md2FF_state_gff_12_n64), .A2(
        md2FF_state_gff_12_n63), .ZN(md2FF_state_gff_12_n30) );
  NAND2_X1 md2FF_state_gff_12_U15 ( .A1(md2FF_state_gff_12_n67), .A2(
        md2FF_permOut[43]), .ZN(md2FF_state_gff_12_n63) );
  MUX2_X1 md2FF_state_gff_12_U14 ( .A(md2FF_state_gff_12_n34), .B(
        md2FF_state_gff_12_n62), .S(md2FF_state_gff_12_n65), .Z(
        md2FF_state_gff_12_n64) );
  NAND2_X1 md2FF_state_gff_12_U13 ( .A1(md2FF_state_n9), .A2(
        md2FF_inputPar[46]), .ZN(md2FF_state_gff_12_n62) );
  NAND2_X1 md2FF_state_gff_12_U12 ( .A1(md2FF_state_gff_12_n61), .A2(
        md2FF_state_gff_12_n60), .ZN(md2FF_state_gff_12_n31) );
  NAND2_X1 md2FF_state_gff_12_U11 ( .A1(md2FF_state_gff_12_n67), .A2(
        md2FF_permOut[27]), .ZN(md2FF_state_gff_12_n60) );
  MUX2_X1 md2FF_state_gff_12_U10 ( .A(md2FF_state_gff_12_n35), .B(
        md2FF_state_gff_12_n59), .S(md2FF_state_gff_12_n65), .Z(
        md2FF_state_gff_12_n61) );
  NAND2_X1 md2FF_state_gff_12_U9 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[45]), .ZN(md2FF_state_gff_12_n59) );
  NAND2_X1 md2FF_state_gff_12_U8 ( .A1(md2FF_state_gff_12_n58), .A2(
        md2FF_state_gff_12_n57), .ZN(md2FF_state_gff_12_n32) );
  NAND2_X1 md2FF_state_gff_12_U7 ( .A1(md2FF_state_gff_12_n67), .A2(
        md2FF_permOut[11]), .ZN(md2FF_state_gff_12_n57) );
  NOR2_X1 md2FF_state_gff_12_U6 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_12_n56), .ZN(md2FF_state_gff_12_n67) );
  MUX2_X1 md2FF_state_gff_12_U5 ( .A(md2FF_state_gff_12_n36), .B(
        md2FF_state_gff_12_n55), .S(md2FF_state_gff_12_n65), .Z(
        md2FF_state_gff_12_n58) );
  INV_X1 md2FF_state_gff_12_U4 ( .A(md2FF_state_gff_12_n56), .ZN(
        md2FF_state_gff_12_n65) );
  INV_X1 md2FF_state_gff_12_U3 ( .A(md2FF_state_n7), .ZN(
        md2FF_state_gff_12_n56) );
  NAND2_X1 md2FF_state_gff_12_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[44]), .ZN(md2FF_state_gff_12_n55) );
DFF_X1 md2FF_state_gff_12_s_current_state_reg_0_ ( .D(md2FF_state_gff_12_n32), .CK(clk), .Q(md2FF_permOut[12]), .QN(md2FF_state_gff_12_n36) );
DFF_X1 md2FF_state_gff_12_s_current_state_reg_1_ ( .D(md2FF_state_gff_12_n31), .CK(clk), .Q(md2FF_permOut[28]), .QN(md2FF_state_gff_12_n35) );
DFF_X1 md2FF_state_gff_12_s_current_state_reg_2_ ( .D(md2FF_state_gff_12_n30), .CK(clk), .Q(md2FF_permOut[44]), .QN(md2FF_state_gff_12_n34) );
DFF_X1 md2FF_state_gff_12_s_current_state_reg_3_ ( .D(md2FF_state_gff_12_n29), .CK(clk), .Q(md2FF_permOut[60]), .QN(md2FF_state_gff_12_n33) );
  NAND2_X1 md2FF_state_gff_13_U20 ( .A1(md2FF_state_gff_13_n69), .A2(
        md2FF_state_gff_13_n68), .ZN(md2FF_state_gff_13_n29) );
  NAND2_X1 md2FF_state_gff_13_U19 ( .A1(md2FF_state_gff_13_n67), .A2(
        md2FF_permOut[60]), .ZN(md2FF_state_gff_13_n68) );
  MUX2_X1 md2FF_state_gff_13_U18 ( .A(md2FF_state_gff_13_n33), .B(
        md2FF_state_gff_13_n66), .S(md2FF_state_gff_13_n65), .Z(
        md2FF_state_gff_13_n69) );
  NAND2_X1 md2FF_state_gff_13_U17 ( .A1(md2FF_state_n9), .A2(
        md2FF_inputPar[51]), .ZN(md2FF_state_gff_13_n66) );
  NAND2_X1 md2FF_state_gff_13_U16 ( .A1(md2FF_state_gff_13_n64), .A2(
        md2FF_state_gff_13_n63), .ZN(md2FF_state_gff_13_n30) );
  NAND2_X1 md2FF_state_gff_13_U15 ( .A1(md2FF_state_gff_13_n67), .A2(
        md2FF_permOut[44]), .ZN(md2FF_state_gff_13_n63) );
  MUX2_X1 md2FF_state_gff_13_U14 ( .A(md2FF_state_gff_13_n34), .B(
        md2FF_state_gff_13_n62), .S(md2FF_state_gff_13_n65), .Z(
        md2FF_state_gff_13_n64) );
  NAND2_X1 md2FF_state_gff_13_U13 ( .A1(md2FF_state_n9), .A2(
        md2FF_inputPar[50]), .ZN(md2FF_state_gff_13_n62) );
  NAND2_X1 md2FF_state_gff_13_U12 ( .A1(md2FF_state_gff_13_n61), .A2(
        md2FF_state_gff_13_n60), .ZN(md2FF_state_gff_13_n31) );
  NAND2_X1 md2FF_state_gff_13_U11 ( .A1(md2FF_state_gff_13_n67), .A2(
        md2FF_permOut[28]), .ZN(md2FF_state_gff_13_n60) );
  MUX2_X1 md2FF_state_gff_13_U10 ( .A(md2FF_state_gff_13_n35), .B(
        md2FF_state_gff_13_n59), .S(md2FF_state_gff_13_n65), .Z(
        md2FF_state_gff_13_n61) );
  NAND2_X1 md2FF_state_gff_13_U9 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[49]), .ZN(md2FF_state_gff_13_n59) );
  NAND2_X1 md2FF_state_gff_13_U8 ( .A1(md2FF_state_gff_13_n58), .A2(
        md2FF_state_gff_13_n57), .ZN(md2FF_state_gff_13_n32) );
  NAND2_X1 md2FF_state_gff_13_U7 ( .A1(md2FF_state_gff_13_n67), .A2(
        md2FF_permOut[12]), .ZN(md2FF_state_gff_13_n57) );
  NOR2_X1 md2FF_state_gff_13_U6 ( .A1(md2FF_state_n9), .A2(
        md2FF_state_gff_13_n56), .ZN(md2FF_state_gff_13_n67) );
  MUX2_X1 md2FF_state_gff_13_U5 ( .A(md2FF_state_gff_13_n36), .B(
        md2FF_state_gff_13_n55), .S(md2FF_state_gff_13_n65), .Z(
        md2FF_state_gff_13_n58) );
  INV_X1 md2FF_state_gff_13_U4 ( .A(md2FF_state_gff_13_n56), .ZN(
        md2FF_state_gff_13_n65) );
  INV_X1 md2FF_state_gff_13_U3 ( .A(md2FF_state_n7), .ZN(
        md2FF_state_gff_13_n56) );
  NAND2_X1 md2FF_state_gff_13_U2 ( .A1(md2FF_state_n9), .A2(md2FF_inputPar[48]), .ZN(md2FF_state_gff_13_n55) );
DFF_X1 md2FF_state_gff_13_s_current_state_reg_0_ ( .D(md2FF_state_gff_13_n32), .CK(clk), .Q(md2FF_permOut[13]), .QN(md2FF_state_gff_13_n36) );
DFF_X1 md2FF_state_gff_13_s_current_state_reg_1_ ( .D(md2FF_state_gff_13_n31), .CK(clk), .Q(md2FF_permOut[29]), .QN(md2FF_state_gff_13_n35) );
DFF_X1 md2FF_state_gff_13_s_current_state_reg_2_ ( .D(md2FF_state_gff_13_n30), .CK(clk), .Q(md2FF_permOut[45]), .QN(md2FF_state_gff_13_n34) );
DFF_X1 md2FF_state_gff_13_s_current_state_reg_3_ ( .D(md2FF_state_gff_13_n29), .CK(clk), .Q(md2FF_permOut[61]), .QN(md2FF_state_gff_13_n33) );
  NAND2_X1 md2FF_state_gff_14_U20 ( .A1(md2FF_state_gff_14_n69), .A2(
        md2FF_state_gff_14_n68), .ZN(md2FF_state_gff_14_n29) );
  NAND2_X1 md2FF_state_gff_14_U19 ( .A1(md2FF_state_gff_14_n67), .A2(
        md2FF_permOut[61]), .ZN(md2FF_state_gff_14_n68) );
  MUX2_X1 md2FF_state_gff_14_U18 ( .A(md2FF_state_gff_14_n33), .B(
        md2FF_state_gff_14_n66), .S(md2FF_state_gff_14_n65), .Z(
        md2FF_state_gff_14_n69) );
  NAND2_X1 md2FF_state_gff_14_U17 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[55]), .ZN(md2FF_state_gff_14_n66) );
  NAND2_X1 md2FF_state_gff_14_U16 ( .A1(md2FF_state_gff_14_n64), .A2(
        md2FF_state_gff_14_n63), .ZN(md2FF_state_gff_14_n30) );
  NAND2_X1 md2FF_state_gff_14_U15 ( .A1(md2FF_state_gff_14_n67), .A2(
        md2FF_permOut[45]), .ZN(md2FF_state_gff_14_n63) );
  MUX2_X1 md2FF_state_gff_14_U14 ( .A(md2FF_state_gff_14_n34), .B(
        md2FF_state_gff_14_n62), .S(md2FF_state_gff_14_n65), .Z(
        md2FF_state_gff_14_n64) );
  NAND2_X1 md2FF_state_gff_14_U13 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[54]), .ZN(md2FF_state_gff_14_n62) );
  NAND2_X1 md2FF_state_gff_14_U12 ( .A1(md2FF_state_gff_14_n61), .A2(
        md2FF_state_gff_14_n60), .ZN(md2FF_state_gff_14_n31) );
  NAND2_X1 md2FF_state_gff_14_U11 ( .A1(md2FF_state_gff_14_n67), .A2(
        md2FF_permOut[29]), .ZN(md2FF_state_gff_14_n60) );
  MUX2_X1 md2FF_state_gff_14_U10 ( .A(md2FF_state_gff_14_n35), .B(
        md2FF_state_gff_14_n59), .S(md2FF_state_gff_14_n65), .Z(
        md2FF_state_gff_14_n61) );
  NAND2_X1 md2FF_state_gff_14_U9 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[53]), .ZN(md2FF_state_gff_14_n59) );
  NAND2_X1 md2FF_state_gff_14_U8 ( .A1(md2FF_state_gff_14_n58), .A2(
        md2FF_state_gff_14_n57), .ZN(md2FF_state_gff_14_n32) );
  NAND2_X1 md2FF_state_gff_14_U7 ( .A1(md2FF_state_gff_14_n67), .A2(
        md2FF_permOut[13]), .ZN(md2FF_state_gff_14_n57) );
  NOR2_X1 md2FF_state_gff_14_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_14_n56), .ZN(md2FF_state_gff_14_n67) );
  MUX2_X1 md2FF_state_gff_14_U5 ( .A(md2FF_state_gff_14_n36), .B(
        md2FF_state_gff_14_n55), .S(md2FF_state_gff_14_n65), .Z(
        md2FF_state_gff_14_n58) );
  INV_X1 md2FF_state_gff_14_U4 ( .A(md2FF_state_gff_14_n56), .ZN(
        md2FF_state_gff_14_n65) );
  INV_X1 md2FF_state_gff_14_U3 ( .A(md2FF_state_n7), .ZN(
        md2FF_state_gff_14_n56) );
  NAND2_X1 md2FF_state_gff_14_U2 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[52]), .ZN(md2FF_state_gff_14_n55) );
DFF_X1 md2FF_state_gff_14_s_current_state_reg_0_ ( .D(md2FF_state_gff_14_n32), .CK(clk), .Q(md2FF_permOut[14]), .QN(md2FF_state_gff_14_n36) );
DFF_X1 md2FF_state_gff_14_s_current_state_reg_1_ ( .D(md2FF_state_gff_14_n31), .CK(clk), .Q(md2FF_permOut[30]), .QN(md2FF_state_gff_14_n35) );
DFF_X1 md2FF_state_gff_14_s_current_state_reg_2_ ( .D(md2FF_state_gff_14_n30), .CK(clk), .Q(md2FF_permOut[46]), .QN(md2FF_state_gff_14_n34) );
DFF_X1 md2FF_state_gff_14_s_current_state_reg_3_ ( .D(md2FF_state_gff_14_n29), .CK(clk), .Q(md2FF_permOut[62]), .QN(md2FF_state_gff_14_n33) );
  NAND2_X1 md2FF_state_gff_15_U20 ( .A1(md2FF_state_gff_15_n68), .A2(
        md2FF_state_gff_15_n67), .ZN(md2FF_state_gff_15_n28) );
  NAND2_X1 md2FF_state_gff_15_U19 ( .A1(md2FF_state_gff_15_n66), .A2(
        md2FF_permOut[62]), .ZN(md2FF_state_gff_15_n67) );
  MUX2_X1 md2FF_state_gff_15_U18 ( .A(md2FF_state_gff_15_n32), .B(
        md2FF_state_gff_15_n65), .S(md2FF_state_gff_15_n64), .Z(
        md2FF_state_gff_15_n68) );
  NAND2_X1 md2FF_state_gff_15_U17 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[59]), .ZN(md2FF_state_gff_15_n65) );
  NAND2_X1 md2FF_state_gff_15_U16 ( .A1(md2FF_state_gff_15_n63), .A2(
        md2FF_state_gff_15_n62), .ZN(md2FF_state_gff_15_n29) );
  NAND2_X1 md2FF_state_gff_15_U15 ( .A1(md2FF_state_gff_15_n66), .A2(
        md2FF_permOut[46]), .ZN(md2FF_state_gff_15_n62) );
  MUX2_X1 md2FF_state_gff_15_U14 ( .A(md2FF_state_gff_15_n33), .B(
        md2FF_state_gff_15_n61), .S(md2FF_state_gff_15_n64), .Z(
        md2FF_state_gff_15_n63) );
  NAND2_X1 md2FF_state_gff_15_U13 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[58]), .ZN(md2FF_state_gff_15_n61) );
  NAND2_X1 md2FF_state_gff_15_U12 ( .A1(md2FF_state_gff_15_n60), .A2(
        md2FF_state_gff_15_n59), .ZN(md2FF_state_gff_15_n30) );
  NAND2_X1 md2FF_state_gff_15_U11 ( .A1(md2FF_state_gff_15_n66), .A2(
        md2FF_permOut[30]), .ZN(md2FF_state_gff_15_n59) );
  MUX2_X1 md2FF_state_gff_15_U10 ( .A(md2FF_state_gff_15_n34), .B(
        md2FF_state_gff_15_n58), .S(md2FF_state_gff_15_n64), .Z(
        md2FF_state_gff_15_n60) );
  NAND2_X1 md2FF_state_gff_15_U9 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[57]), .ZN(md2FF_state_gff_15_n58) );
  NAND2_X1 md2FF_state_gff_15_U8 ( .A1(md2FF_state_gff_15_n57), .A2(
        md2FF_state_gff_15_n56), .ZN(md2FF_state_gff_15_n31) );
  NAND2_X1 md2FF_state_gff_15_U7 ( .A1(md2FF_state_gff_15_n66), .A2(
        md2FF_permOut[14]), .ZN(md2FF_state_gff_15_n56) );
  NOR2_X1 md2FF_state_gff_15_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_15_n55), .ZN(md2FF_state_gff_15_n66) );
  MUX2_X1 md2FF_state_gff_15_U5 ( .A(md2FF_state_gff_15_n35), .B(
        md2FF_state_gff_15_n54), .S(md2FF_state_gff_15_n64), .Z(
        md2FF_state_gff_15_n57) );
  INV_X1 md2FF_state_gff_15_U4 ( .A(md2FF_state_gff_15_n55), .ZN(
        md2FF_state_gff_15_n64) );
  INV_X1 md2FF_state_gff_15_U3 ( .A(md2FF_state_n7), .ZN(
        md2FF_state_gff_15_n55) );
  NAND2_X1 md2FF_state_gff_15_U2 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[56]), .ZN(md2FF_state_gff_15_n54) );
DFF_X1 md2FF_state_gff_15_s_current_state_reg_0_ ( .D(md2FF_state_gff_15_n31), .CK(clk), .Q(md2FF_permOut[15]), .QN(md2FF_state_gff_15_n35) );
DFF_X1 md2FF_state_gff_15_s_current_state_reg_1_ ( .D(md2FF_state_gff_15_n30), .CK(clk), .Q(md2FF_permOut[31]), .QN(md2FF_state_gff_15_n34) );
DFF_X1 md2FF_state_gff_15_s_current_state_reg_2_ ( .D(md2FF_state_gff_15_n29), .CK(clk), .Q(md2FF_permOut[47]), .QN(md2FF_state_gff_15_n33) );
DFF_X1 md2FF_state_gff_15_s_current_state_reg_3_ ( .D(md2FF_state_gff_15_n28), .CK(clk), .Q(md2FF_permOut[63]), .QN(md2FF_state_gff_15_n32) );
  NAND2_X1 md2FF_state_gff_16_U20 ( .A1(md2FF_state_gff_16_n68), .A2(
        md2FF_state_gff_16_n67), .ZN(md2FF_state_gff_16_n28) );
  NAND2_X1 md2FF_state_gff_16_U19 ( .A1(md2FF_state_gff_16_n66), .A2(
        md2FF_permOut[63]), .ZN(md2FF_state_gff_16_n67) );
  MUX2_X1 md2FF_state_gff_16_U18 ( .A(md2FF_state_gff_16_n32), .B(
        md2FF_state_gff_16_n65), .S(md2FF_state_gff_16_n64), .Z(
        md2FF_state_gff_16_n68) );
  NAND2_X1 md2FF_state_gff_16_U17 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[63]), .ZN(md2FF_state_gff_16_n65) );
  NAND2_X1 md2FF_state_gff_16_U16 ( .A1(md2FF_state_gff_16_n63), .A2(
        md2FF_state_gff_16_n62), .ZN(md2FF_state_gff_16_n29) );
  NAND2_X1 md2FF_state_gff_16_U15 ( .A1(md2FF_state_gff_16_n66), .A2(
        md2FF_permOut[47]), .ZN(md2FF_state_gff_16_n62) );
  MUX2_X1 md2FF_state_gff_16_U14 ( .A(md2FF_state_gff_16_n33), .B(
        md2FF_state_gff_16_n61), .S(md2FF_state_gff_16_n64), .Z(
        md2FF_state_gff_16_n63) );
  NAND2_X1 md2FF_state_gff_16_U13 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[62]), .ZN(md2FF_state_gff_16_n61) );
  NAND2_X1 md2FF_state_gff_16_U12 ( .A1(md2FF_state_gff_16_n60), .A2(
        md2FF_state_gff_16_n59), .ZN(md2FF_state_gff_16_n30) );
  NAND2_X1 md2FF_state_gff_16_U11 ( .A1(md2FF_state_gff_16_n66), .A2(
        md2FF_permOut[31]), .ZN(md2FF_state_gff_16_n59) );
  MUX2_X1 md2FF_state_gff_16_U10 ( .A(md2FF_state_gff_16_n34), .B(
        md2FF_state_gff_16_n58), .S(md2FF_state_gff_16_n64), .Z(
        md2FF_state_gff_16_n60) );
  NAND2_X1 md2FF_state_gff_16_U9 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[61]), .ZN(md2FF_state_gff_16_n58) );
  NAND2_X1 md2FF_state_gff_16_U8 ( .A1(md2FF_state_gff_16_n57), .A2(
        md2FF_state_gff_16_n56), .ZN(md2FF_state_gff_16_n31) );
  NAND2_X1 md2FF_state_gff_16_U7 ( .A1(md2FF_state_gff_16_n66), .A2(
        md2FF_permOut[15]), .ZN(md2FF_state_gff_16_n56) );
  NOR2_X1 md2FF_state_gff_16_U6 ( .A1(md2FF_state_n10), .A2(
        md2FF_state_gff_16_n55), .ZN(md2FF_state_gff_16_n66) );
  MUX2_X1 md2FF_state_gff_16_U5 ( .A(md2FF_state_gff_16_n35), .B(
        md2FF_state_gff_16_n54), .S(md2FF_state_gff_16_n64), .Z(
        md2FF_state_gff_16_n57) );
  INV_X1 md2FF_state_gff_16_U4 ( .A(md2FF_state_gff_16_n55), .ZN(
        md2FF_state_gff_16_n64) );
  INV_X1 md2FF_state_gff_16_U3 ( .A(md2FF_state_n7), .ZN(
        md2FF_state_gff_16_n55) );
  NAND2_X1 md2FF_state_gff_16_U2 ( .A1(md2FF_state_n10), .A2(
        md2FF_inputPar[60]), .ZN(md2FF_state_gff_16_n54) );
DFF_X1 md2FF_state_gff_16_s_current_state_reg_0_ ( .D(md2FF_state_gff_16_n31), .CK(clk), .Q(md2Reg[0]), .QN(md2FF_state_gff_16_n35) );
DFF_X1 md2FF_state_gff_16_s_current_state_reg_1_ ( .D(md2FF_state_gff_16_n30), .CK(clk), .Q(md2Reg[1]), .QN(md2FF_state_gff_16_n34) );
DFF_X1 md2FF_state_gff_16_s_current_state_reg_2_ ( .D(md2FF_state_gff_16_n29), .CK(clk), .Q(md2Reg[2]), .QN(md2FF_state_gff_16_n33) );
DFF_X1 md2FF_state_gff_16_s_current_state_reg_3_ ( .D(md2FF_state_gff_16_n28), .CK(clk), .Q(md2Reg[3]), .QN(md2FF_state_gff_16_n32) );
  MUX2_X1 keyFF_U91 ( .A(sboxOut[3]), .B(key[79]), .S(ctrlData[2]), .Z(
        keyFF_inputPar[79]) );
  MUX2_X1 keyFF_U90 ( .A(sboxOut[2]), .B(key[78]), .S(ctrlData[2]), .Z(
        keyFF_inputPar[78]) );
  MUX2_X1 keyFF_U89 ( .A(sboxOut[1]), .B(key[77]), .S(ctrlData[2]), .Z(
        keyFF_inputPar[77]) );
  MUX2_X1 keyFF_U88 ( .A(sboxOut[0]), .B(key[76]), .S(keyFF_n183), .Z(
        keyFF_inputPar[76]) );
  MUX2_X1 keyFF_U87 ( .A(roundkey[2]), .B(key[75]), .S(keyFF_n182), .Z(
        keyFF_inputPar[75]) );
  MUX2_X1 keyFF_U86 ( .A(keyFF_outputPar[12]), .B(key[9]), .S(keyFF_n181), .Z(
        keyFF_inputPar[9]) );
  MUX2_X1 keyFF_U85 ( .A(keyFF_outputPar[11]), .B(key[8]), .S(keyFF_n180), .Z(
        keyFF_inputPar[8]) );
  MUX2_X1 keyFF_U84 ( .A(keyFF_outputPar[10]), .B(key[7]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[7]) );
  MUX2_X1 keyFF_U83 ( .A(roundkey[1]), .B(key[74]), .S(ctrlData[2]), .Z(
        keyFF_inputPar[74]) );
  MUX2_X1 keyFF_U82 ( .A(roundkey[0]), .B(key[73]), .S(ctrlData[2]), .Z(
        keyFF_inputPar[73]) );
  MUX2_X1 keyFF_U81 ( .A(keyFF_outputPar[75]), .B(key[72]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[72]) );
  MUX2_X1 keyFF_U80 ( .A(keyFF_outputPar[74]), .B(key[71]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[71]) );
  MUX2_X1 keyFF_U79 ( .A(keyFF_outputPar[73]), .B(key[70]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[70]) );
  MUX2_X1 keyFF_U78 ( .A(keyFF_outputPar[72]), .B(key[69]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[69]) );
  MUX2_X1 keyFF_U77 ( .A(keyFF_outputPar[71]), .B(key[68]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[68]) );
  MUX2_X1 keyFF_U76 ( .A(keyFF_outputPar[70]), .B(key[67]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[67]) );
  MUX2_X1 keyFF_U75 ( .A(keyFF_outputPar[69]), .B(key[66]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[66]) );
  MUX2_X1 keyFF_U74 ( .A(keyFF_outputPar[68]), .B(key[65]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[65]) );
  MUX2_X1 keyFF_U73 ( .A(keyFF_outputPar[67]), .B(key[64]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[64]) );
  MUX2_X1 keyFF_U72 ( .A(keyFF_outputPar[66]), .B(key[63]), .S(ctrlData[2]), 
        .Z(keyFF_inputPar[63]) );
  MUX2_X1 keyFF_U71 ( .A(keyFF_outputPar[65]), .B(key[62]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[62]) );
  MUX2_X1 keyFF_U70 ( .A(keyFF_outputPar[64]), .B(key[61]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[61]) );
  MUX2_X1 keyFF_U69 ( .A(keyFF_outputPar[63]), .B(key[60]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[60]) );
  MUX2_X1 keyFF_U68 ( .A(keyFF_outputPar[62]), .B(key[59]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[59]) );
  MUX2_X1 keyFF_U67 ( .A(keyFF_outputPar[61]), .B(key[58]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[58]) );
  MUX2_X1 keyFF_U66 ( .A(keyFF_outputPar[60]), .B(key[57]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[57]) );
  MUX2_X1 keyFF_U65 ( .A(keyFF_outputPar[59]), .B(key[56]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[56]) );
  MUX2_X1 keyFF_U64 ( .A(keyFF_outputPar[58]), .B(key[55]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[55]) );
  MUX2_X1 keyFF_U63 ( .A(keyFF_outputPar[57]), .B(key[54]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[54]) );
  MUX2_X1 keyFF_U62 ( .A(keyFF_outputPar[56]), .B(key[53]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[53]) );
  MUX2_X1 keyFF_U61 ( .A(keyFF_outputPar[55]), .B(key[52]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[52]) );
  MUX2_X1 keyFF_U60 ( .A(keyFF_outputPar[54]), .B(key[51]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[51]) );
  MUX2_X1 keyFF_U59 ( .A(keyFF_outputPar[53]), .B(key[50]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[50]) );
  MUX2_X1 keyFF_U58 ( .A(keyFF_outputPar[52]), .B(key[49]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[49]) );
  MUX2_X1 keyFF_U57 ( .A(keyFF_outputPar[51]), .B(key[48]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[48]) );
  MUX2_X1 keyFF_U56 ( .A(keyFF_outputPar[50]), .B(key[47]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[47]) );
  MUX2_X1 keyFF_U55 ( .A(keyFF_outputPar[49]), .B(key[46]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[46]) );
  MUX2_X1 keyFF_U54 ( .A(keyFF_outputPar[48]), .B(key[45]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[45]) );
  MUX2_X1 keyFF_U53 ( .A(keyFF_outputPar[47]), .B(key[44]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[44]) );
  MUX2_X1 keyFF_U52 ( .A(keyFF_outputPar[46]), .B(key[43]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[43]) );
  MUX2_X1 keyFF_U51 ( .A(keyFF_outputPar[45]), .B(key[42]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[42]) );
  MUX2_X1 keyFF_U50 ( .A(keyFF_outputPar[44]), .B(key[41]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[41]) );
  MUX2_X1 keyFF_U49 ( .A(keyFF_outputPar[43]), .B(key[40]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[40]) );
  MUX2_X1 keyFF_U48 ( .A(keyFF_outputPar[42]), .B(key[39]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[39]) );
  MUX2_X1 keyFF_U47 ( .A(keyFF_outputPar[41]), .B(key[38]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[38]) );
  MUX2_X1 keyFF_U46 ( .A(keyFF_outputPar[40]), .B(key[37]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[37]) );
  MUX2_X1 keyFF_U45 ( .A(keyFF_outputPar[39]), .B(key[36]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[36]) );
  MUX2_X1 keyFF_U44 ( .A(keyFF_outputPar[38]), .B(key[35]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[35]) );
  MUX2_X1 keyFF_U43 ( .A(keyFF_outputPar[37]), .B(key[34]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[34]) );
  MUX2_X1 keyFF_U42 ( .A(keyFF_outputPar[36]), .B(key[33]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[33]) );
  MUX2_X1 keyFF_U41 ( .A(keyFF_outputPar[35]), .B(key[32]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[32]) );
  MUX2_X1 keyFF_U40 ( .A(keyFF_outputPar[34]), .B(key[31]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[31]) );
  MUX2_X1 keyFF_U39 ( .A(keyFF_outputPar[33]), .B(key[30]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[30]) );
  MUX2_X1 keyFF_U38 ( .A(keyFF_outputPar[32]), .B(key[29]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[29]) );
  MUX2_X1 keyFF_U37 ( .A(keyFF_outputPar[31]), .B(key[28]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[28]) );
  MUX2_X1 keyFF_U36 ( .A(keyFF_outputPar[30]), .B(key[27]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[27]) );
  MUX2_X1 keyFF_U35 ( .A(keyFF_outputPar[29]), .B(key[26]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[26]) );
  MUX2_X1 keyFF_U34 ( .A(keyFF_outputPar[28]), .B(key[25]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[25]) );
  MUX2_X1 keyFF_U33 ( .A(keyFF_outputPar[27]), .B(key[24]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[24]) );
  MUX2_X1 keyFF_U32 ( .A(keyFF_outputPar[26]), .B(key[23]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[23]) );
  MUX2_X1 keyFF_U31 ( .A(keyFF_outputPar[25]), .B(key[22]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[22]) );
  MUX2_X1 keyFF_U30 ( .A(keyFF_outputPar[24]), .B(key[21]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[21]) );
  MUX2_X1 keyFF_U29 ( .A(keyFF_outputPar[23]), .B(key[20]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[20]) );
  MUX2_X1 keyFF_U28 ( .A(keyFF_n179), .B(key[19]), .S(keyFF_n183), .Z(
        keyFF_inputPar[19]) );
  XOR2_X1 keyFF_U27 ( .A(counter[4]), .B(keyFF_outputPar[22]), .Z(keyFF_n179)
         );
  MUX2_X1 keyFF_U26 ( .A(keyFF_n178), .B(key[18]), .S(keyFF_n183), .Z(
        keyFF_inputPar[18]) );
  XOR2_X1 keyFF_U25 ( .A(counter[3]), .B(keyFF_outputPar[21]), .Z(keyFF_n178)
         );
  MUX2_X1 keyFF_U24 ( .A(keyFF_n177), .B(key[17]), .S(keyFF_n183), .Z(
        keyFF_inputPar[17]) );
  XOR2_X1 keyFF_U23 ( .A(counter[2]), .B(keyFF_outputPar[20]), .Z(keyFF_n177)
         );
  MUX2_X1 keyFF_U22 ( .A(keyFF_n176), .B(key[16]), .S(keyFF_n183), .Z(
        keyFF_inputPar[16]) );
  XOR2_X1 keyFF_U21 ( .A(counter[1]), .B(keyFF_outputPar[19]), .Z(keyFF_n176)
         );
  MUX2_X1 keyFF_U20 ( .A(keyFF_n175), .B(key[15]), .S(keyFF_n183), .Z(
        keyFF_inputPar[15]) );
  XOR2_X1 keyFF_U19 ( .A(counter[0]), .B(keyFF_outputPar[18]), .Z(keyFF_n175)
         );
  MUX2_X1 keyFF_U18 ( .A(keyFF_outputPar[17]), .B(key[14]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[14]) );
  MUX2_X1 keyFF_U17 ( .A(keyFF_outputPar[16]), .B(key[13]), .S(keyFF_n182), 
        .Z(keyFF_inputPar[13]) );
  MUX2_X1 keyFF_U16 ( .A(keyFF_outputPar[15]), .B(key[12]), .S(keyFF_n181), 
        .Z(keyFF_inputPar[12]) );
  MUX2_X1 keyFF_U15 ( .A(keyFF_outputPar[14]), .B(key[11]), .S(keyFF_n180), 
        .Z(keyFF_inputPar[11]) );
  MUX2_X1 keyFF_U14 ( .A(keyFF_outputPar[13]), .B(key[10]), .S(keyFF_n183), 
        .Z(keyFF_inputPar[10]) );
  MUX2_X1 keyFF_U13 ( .A(keyFF_outputPar[9]), .B(key[6]), .S(keyFF_n182), .Z(
        keyFF_inputPar[6]) );
  MUX2_X1 keyFF_U12 ( .A(keyFF_outputPar[8]), .B(key[5]), .S(keyFF_n181), .Z(
        keyFF_inputPar[5]) );
  MUX2_X1 keyFF_U11 ( .A(keyFF_outputPar[7]), .B(key[4]), .S(keyFF_n180), .Z(
        keyFF_inputPar[4]) );
  MUX2_X1 keyFF_U10 ( .A(keyFF_outputPar[6]), .B(key[3]), .S(keyFF_n183), .Z(
        keyFF_inputPar[3]) );
  INV_X1 keyFF_U9 ( .A(keyFF_n174), .ZN(keyFF_n183) );
  MUX2_X1 keyFF_U8 ( .A(keyFF_outputPar[5]), .B(key[2]), .S(keyFF_n182), .Z(
        keyFF_inputPar[2]) );
  INV_X1 keyFF_U7 ( .A(keyFF_n174), .ZN(keyFF_n182) );
  MUX2_X1 keyFF_U6 ( .A(keyFF_outputPar[4]), .B(key[1]), .S(keyFF_n181), .Z(
        keyFF_inputPar[1]) );
  INV_X1 keyFF_U5 ( .A(keyFF_n174), .ZN(keyFF_n181) );
  MUX2_X1 keyFF_U4 ( .A(keyFF_outputPar[3]), .B(key[0]), .S(keyFF_n180), .Z(
        keyFF_inputPar[0]) );
  INV_X1 keyFF_U3 ( .A(keyFF_n174), .ZN(keyFF_n180) );
  INV_X1 keyFF_U2 ( .A(ctrlData[2]), .ZN(keyFF_n174) );
  INV_X2 keyFF_keystate_U3 ( .A(keyFF_keystate_n8), .ZN(keyFF_keystate_n7) );
  INV_X2 keyFF_keystate_U2 ( .A(keyFF_keystate_n8), .ZN(keyFF_keystate_n6) );
  INV_X1 keyFF_keystate_U1 ( .A(ctrlData[0]), .ZN(keyFF_keystate_n8) );
  NAND2_X1 keyFF_keystate_gff_1_U19 ( .A1(keyFF_keystate_gff_1_n68), .A2(
        keyFF_keystate_gff_1_n67), .ZN(keyFF_keystate_gff_1_n30) );
  NAND2_X1 keyFF_keystate_gff_1_U18 ( .A1(keyFF_keystate_gff_1_n66), .A2(
        roundkey[2]), .ZN(keyFF_keystate_gff_1_n67) );
  MUX2_X1 keyFF_keystate_gff_1_U17 ( .A(keyFF_keystate_gff_1_n34), .B(
        keyFF_keystate_gff_1_n65), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_1_n68) );
  NAND2_X1 keyFF_keystate_gff_1_U16 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[2]), 
        .ZN(keyFF_keystate_gff_1_n65) );
  NAND2_X1 keyFF_keystate_gff_1_U15 ( .A1(keyFF_keystate_gff_1_n64), .A2(
        keyFF_keystate_gff_1_n63), .ZN(keyFF_keystate_gff_1_n31) );
  NAND2_X1 keyFF_keystate_gff_1_U14 ( .A1(keyFF_keystate_gff_1_n66), .A2(
        roundkey[1]), .ZN(keyFF_keystate_gff_1_n63) );
  MUX2_X1 keyFF_keystate_gff_1_U13 ( .A(keyFF_keystate_gff_1_n35), .B(
        keyFF_keystate_gff_1_n62), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_1_n64) );
  NAND2_X1 keyFF_keystate_gff_1_U12 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[1]), 
        .ZN(keyFF_keystate_gff_1_n62) );
  NAND2_X1 keyFF_keystate_gff_1_U11 ( .A1(keyFF_keystate_gff_1_n61), .A2(
        keyFF_keystate_gff_1_n60), .ZN(keyFF_keystate_gff_1_n32) );
  NAND2_X1 keyFF_keystate_gff_1_U10 ( .A1(keyFF_keystate_gff_1_n66), .A2(
        roundkey[0]), .ZN(keyFF_keystate_gff_1_n60) );
  MUX2_X1 keyFF_keystate_gff_1_U9 ( .A(keyFF_keystate_gff_1_n36), .B(
        keyFF_keystate_gff_1_n59), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_1_n61) );
  NAND2_X1 keyFF_keystate_gff_1_U8 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[0]), 
        .ZN(keyFF_keystate_gff_1_n59) );
  NAND2_X1 keyFF_keystate_gff_1_U7 ( .A1(keyFF_keystate_gff_1_n58), .A2(
        keyFF_keystate_gff_1_n57), .ZN(keyFF_keystate_gff_1_n29) );
  NAND2_X1 keyFF_keystate_gff_1_U6 ( .A1(keyFF_keystate_gff_1_n66), .A2(
        roundkey[3]), .ZN(keyFF_keystate_gff_1_n57) );
  NOR2_X1 keyFF_keystate_gff_1_U5 ( .A1(ctrlData[0]), .A2(
        keyFF_keystate_gff_1_n56), .ZN(keyFF_keystate_gff_1_n66) );
  INV_X1 keyFF_keystate_gff_1_U4 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_1_n56) );
  MUX2_X1 keyFF_keystate_gff_1_U3 ( .A(keyFF_keystate_gff_1_n33), .B(
        keyFF_keystate_gff_1_n55), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_1_n58) );
  NAND2_X1 keyFF_keystate_gff_1_U2 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[3]), 
        .ZN(keyFF_keystate_gff_1_n55) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_1_n32), .CK(clk), .Q(keyRegKS[1]), .QN(
        keyFF_keystate_gff_1_n36) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_1_n31), .CK(clk), .Q(keyRegKS[2]), .QN(
        keyFF_keystate_gff_1_n35) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_1_n30), .CK(clk), .Q(keyRegKS[3]), .QN(
        keyFF_keystate_gff_1_n34) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_1_n29), .CK(clk), .Q(keyFF_outputPar[3]), .QN(
        keyFF_keystate_gff_1_n33) );
  NAND2_X1 keyFF_keystate_gff_2_U19 ( .A1(keyFF_keystate_gff_2_n68), .A2(
        keyFF_keystate_gff_2_n67), .ZN(keyFF_keystate_gff_2_n29) );
  NAND2_X1 keyFF_keystate_gff_2_U18 ( .A1(keyFF_keystate_gff_2_n66), .A2(
        keyFF_outputPar[3]), .ZN(keyFF_keystate_gff_2_n67) );
  MUX2_X1 keyFF_keystate_gff_2_U17 ( .A(keyFF_keystate_gff_2_n33), .B(
        keyFF_keystate_gff_2_n65), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_2_n68) );
  NAND2_X1 keyFF_keystate_gff_2_U16 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[7]), 
        .ZN(keyFF_keystate_gff_2_n65) );
  NAND2_X1 keyFF_keystate_gff_2_U15 ( .A1(keyFF_keystate_gff_2_n64), .A2(
        keyFF_keystate_gff_2_n63), .ZN(keyFF_keystate_gff_2_n32) );
  NAND2_X1 keyFF_keystate_gff_2_U14 ( .A1(keyFF_keystate_gff_2_n66), .A2(
        keyRegKS[1]), .ZN(keyFF_keystate_gff_2_n63) );
  MUX2_X1 keyFF_keystate_gff_2_U13 ( .A(keyFF_keystate_gff_2_n36), .B(
        keyFF_keystate_gff_2_n62), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_2_n64) );
  NAND2_X1 keyFF_keystate_gff_2_U12 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[4]), 
        .ZN(keyFF_keystate_gff_2_n62) );
  NAND2_X1 keyFF_keystate_gff_2_U11 ( .A1(keyFF_keystate_gff_2_n61), .A2(
        keyFF_keystate_gff_2_n60), .ZN(keyFF_keystate_gff_2_n31) );
  NAND2_X1 keyFF_keystate_gff_2_U10 ( .A1(keyFF_keystate_gff_2_n66), .A2(
        keyRegKS[2]), .ZN(keyFF_keystate_gff_2_n60) );
  MUX2_X1 keyFF_keystate_gff_2_U9 ( .A(keyFF_keystate_gff_2_n35), .B(
        keyFF_keystate_gff_2_n59), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_2_n61) );
  NAND2_X1 keyFF_keystate_gff_2_U8 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[5]), 
        .ZN(keyFF_keystate_gff_2_n59) );
  NAND2_X1 keyFF_keystate_gff_2_U7 ( .A1(keyFF_keystate_gff_2_n58), .A2(
        keyFF_keystate_gff_2_n57), .ZN(keyFF_keystate_gff_2_n30) );
  NAND2_X1 keyFF_keystate_gff_2_U6 ( .A1(keyFF_keystate_gff_2_n66), .A2(
        keyRegKS[3]), .ZN(keyFF_keystate_gff_2_n57) );
  NOR2_X1 keyFF_keystate_gff_2_U5 ( .A1(ctrlData[0]), .A2(
        keyFF_keystate_gff_2_n56), .ZN(keyFF_keystate_gff_2_n66) );
  INV_X1 keyFF_keystate_gff_2_U4 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_2_n56) );
  MUX2_X1 keyFF_keystate_gff_2_U3 ( .A(keyFF_keystate_gff_2_n34), .B(
        keyFF_keystate_gff_2_n55), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_2_n58) );
  NAND2_X1 keyFF_keystate_gff_2_U2 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[6]), 
        .ZN(keyFF_keystate_gff_2_n55) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_2_n32), .CK(clk), .Q(keyFF_outputPar[4]), .QN(
        keyFF_keystate_gff_2_n36) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_2_n31), .CK(clk), .Q(keyFF_outputPar[5]), .QN(
        keyFF_keystate_gff_2_n35) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_2_n30), .CK(clk), .Q(keyFF_outputPar[6]), .QN(
        keyFF_keystate_gff_2_n34) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_2_n29), .CK(clk), .Q(keyFF_outputPar[7]), .QN(
        keyFF_keystate_gff_2_n33) );
  NAND2_X1 keyFF_keystate_gff_3_U19 ( .A1(keyFF_keystate_gff_3_n68), .A2(
        keyFF_keystate_gff_3_n67), .ZN(keyFF_keystate_gff_3_n29) );
  NAND2_X1 keyFF_keystate_gff_3_U18 ( .A1(keyFF_keystate_gff_3_n66), .A2(
        keyFF_outputPar[7]), .ZN(keyFF_keystate_gff_3_n67) );
  MUX2_X1 keyFF_keystate_gff_3_U17 ( .A(keyFF_keystate_gff_3_n33), .B(
        keyFF_keystate_gff_3_n65), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_3_n68) );
  NAND2_X1 keyFF_keystate_gff_3_U16 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[11]), .ZN(keyFF_keystate_gff_3_n65) );
  NAND2_X1 keyFF_keystate_gff_3_U15 ( .A1(keyFF_keystate_gff_3_n64), .A2(
        keyFF_keystate_gff_3_n63), .ZN(keyFF_keystate_gff_3_n30) );
  NAND2_X1 keyFF_keystate_gff_3_U14 ( .A1(keyFF_keystate_gff_3_n66), .A2(
        keyFF_outputPar[6]), .ZN(keyFF_keystate_gff_3_n63) );
  MUX2_X1 keyFF_keystate_gff_3_U13 ( .A(keyFF_keystate_gff_3_n34), .B(
        keyFF_keystate_gff_3_n62), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_3_n64) );
  NAND2_X1 keyFF_keystate_gff_3_U12 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[10]), .ZN(keyFF_keystate_gff_3_n62) );
  NAND2_X1 keyFF_keystate_gff_3_U11 ( .A1(keyFF_keystate_gff_3_n61), .A2(
        keyFF_keystate_gff_3_n60), .ZN(keyFF_keystate_gff_3_n31) );
  NAND2_X1 keyFF_keystate_gff_3_U10 ( .A1(keyFF_keystate_gff_3_n66), .A2(
        keyFF_outputPar[5]), .ZN(keyFF_keystate_gff_3_n60) );
  MUX2_X1 keyFF_keystate_gff_3_U9 ( .A(keyFF_keystate_gff_3_n35), .B(
        keyFF_keystate_gff_3_n59), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_3_n61) );
  NAND2_X1 keyFF_keystate_gff_3_U8 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[9]), 
        .ZN(keyFF_keystate_gff_3_n59) );
  NAND2_X1 keyFF_keystate_gff_3_U7 ( .A1(keyFF_keystate_gff_3_n58), .A2(
        keyFF_keystate_gff_3_n57), .ZN(keyFF_keystate_gff_3_n32) );
  NAND2_X1 keyFF_keystate_gff_3_U6 ( .A1(keyFF_keystate_gff_3_n66), .A2(
        keyFF_outputPar[4]), .ZN(keyFF_keystate_gff_3_n57) );
  NOR2_X1 keyFF_keystate_gff_3_U5 ( .A1(ctrlData[0]), .A2(
        keyFF_keystate_gff_3_n56), .ZN(keyFF_keystate_gff_3_n66) );
  INV_X1 keyFF_keystate_gff_3_U4 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_3_n56) );
  MUX2_X1 keyFF_keystate_gff_3_U3 ( .A(keyFF_keystate_gff_3_n36), .B(
        keyFF_keystate_gff_3_n55), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_3_n58) );
  NAND2_X1 keyFF_keystate_gff_3_U2 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[8]), 
        .ZN(keyFF_keystate_gff_3_n55) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_3_n32), .CK(clk), .Q(keyFF_outputPar[8]), .QN(
        keyFF_keystate_gff_3_n36) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_3_n31), .CK(clk), .Q(keyFF_outputPar[9]), .QN(
        keyFF_keystate_gff_3_n35) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_3_n30), .CK(clk), .Q(keyFF_outputPar[10]), .QN(
        keyFF_keystate_gff_3_n34) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_3_n29), .CK(clk), .Q(keyFF_outputPar[11]), .QN(
        keyFF_keystate_gff_3_n33) );
  NAND2_X1 keyFF_keystate_gff_4_U19 ( .A1(keyFF_keystate_gff_4_n68), .A2(
        keyFF_keystate_gff_4_n67), .ZN(keyFF_keystate_gff_4_n29) );
  NAND2_X1 keyFF_keystate_gff_4_U18 ( .A1(keyFF_keystate_gff_4_n66), .A2(
        keyFF_outputPar[11]), .ZN(keyFF_keystate_gff_4_n67) );
  MUX2_X1 keyFF_keystate_gff_4_U17 ( .A(keyFF_keystate_gff_4_n33), .B(
        keyFF_keystate_gff_4_n65), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_4_n68) );
  NAND2_X1 keyFF_keystate_gff_4_U16 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[15]), .ZN(keyFF_keystate_gff_4_n65) );
  NAND2_X1 keyFF_keystate_gff_4_U15 ( .A1(keyFF_keystate_gff_4_n64), .A2(
        keyFF_keystate_gff_4_n63), .ZN(keyFF_keystate_gff_4_n30) );
  NAND2_X1 keyFF_keystate_gff_4_U14 ( .A1(keyFF_keystate_gff_4_n66), .A2(
        keyFF_outputPar[10]), .ZN(keyFF_keystate_gff_4_n63) );
  MUX2_X1 keyFF_keystate_gff_4_U13 ( .A(keyFF_keystate_gff_4_n34), .B(
        keyFF_keystate_gff_4_n62), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_4_n64) );
  NAND2_X1 keyFF_keystate_gff_4_U12 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[14]), .ZN(keyFF_keystate_gff_4_n62) );
  NAND2_X1 keyFF_keystate_gff_4_U11 ( .A1(keyFF_keystate_gff_4_n61), .A2(
        keyFF_keystate_gff_4_n60), .ZN(keyFF_keystate_gff_4_n31) );
  NAND2_X1 keyFF_keystate_gff_4_U10 ( .A1(keyFF_keystate_gff_4_n66), .A2(
        keyFF_outputPar[9]), .ZN(keyFF_keystate_gff_4_n60) );
  MUX2_X1 keyFF_keystate_gff_4_U9 ( .A(keyFF_keystate_gff_4_n35), .B(
        keyFF_keystate_gff_4_n59), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_4_n61) );
  NAND2_X1 keyFF_keystate_gff_4_U8 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[13]), 
        .ZN(keyFF_keystate_gff_4_n59) );
  NAND2_X1 keyFF_keystate_gff_4_U7 ( .A1(keyFF_keystate_gff_4_n58), .A2(
        keyFF_keystate_gff_4_n57), .ZN(keyFF_keystate_gff_4_n32) );
  NAND2_X1 keyFF_keystate_gff_4_U6 ( .A1(keyFF_keystate_gff_4_n66), .A2(
        keyFF_outputPar[8]), .ZN(keyFF_keystate_gff_4_n57) );
  NOR2_X1 keyFF_keystate_gff_4_U5 ( .A1(ctrlData[0]), .A2(
        keyFF_keystate_gff_4_n56), .ZN(keyFF_keystate_gff_4_n66) );
  INV_X1 keyFF_keystate_gff_4_U4 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_4_n56) );
  MUX2_X1 keyFF_keystate_gff_4_U3 ( .A(keyFF_keystate_gff_4_n36), .B(
        keyFF_keystate_gff_4_n55), .S(ctrlData[1]), .Z(
        keyFF_keystate_gff_4_n58) );
  NAND2_X1 keyFF_keystate_gff_4_U2 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[12]), 
        .ZN(keyFF_keystate_gff_4_n55) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_4_n32), .CK(clk), .Q(keyFF_outputPar[12]), .QN(
        keyFF_keystate_gff_4_n36) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_4_n31), .CK(clk), .Q(keyFF_outputPar[13]), .QN(
        keyFF_keystate_gff_4_n35) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_4_n30), .CK(clk), .Q(keyFF_outputPar[14]), .QN(
        keyFF_keystate_gff_4_n34) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_4_n29), .CK(clk), .Q(keyFF_outputPar[15]), .QN(
        keyFF_keystate_gff_4_n33) );
  NAND2_X1 keyFF_keystate_gff_5_U20 ( .A1(keyFF_keystate_gff_5_n69), .A2(
        keyFF_keystate_gff_5_n68), .ZN(keyFF_keystate_gff_5_n29) );
  NAND2_X1 keyFF_keystate_gff_5_U19 ( .A1(keyFF_keystate_gff_5_n67), .A2(
        keyFF_outputPar[15]), .ZN(keyFF_keystate_gff_5_n68) );
  MUX2_X1 keyFF_keystate_gff_5_U18 ( .A(keyFF_keystate_gff_5_n33), .B(
        keyFF_keystate_gff_5_n66), .S(keyFF_keystate_gff_5_n65), .Z(
        keyFF_keystate_gff_5_n69) );
  NAND2_X1 keyFF_keystate_gff_5_U17 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[19]), .ZN(keyFF_keystate_gff_5_n66) );
  NAND2_X1 keyFF_keystate_gff_5_U16 ( .A1(keyFF_keystate_gff_5_n64), .A2(
        keyFF_keystate_gff_5_n63), .ZN(keyFF_keystate_gff_5_n30) );
  NAND2_X1 keyFF_keystate_gff_5_U15 ( .A1(keyFF_keystate_gff_5_n67), .A2(
        keyFF_outputPar[14]), .ZN(keyFF_keystate_gff_5_n63) );
  MUX2_X1 keyFF_keystate_gff_5_U14 ( .A(keyFF_keystate_gff_5_n34), .B(
        keyFF_keystate_gff_5_n62), .S(keyFF_keystate_gff_5_n65), .Z(
        keyFF_keystate_gff_5_n64) );
  NAND2_X1 keyFF_keystate_gff_5_U13 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[18]), .ZN(keyFF_keystate_gff_5_n62) );
  NAND2_X1 keyFF_keystate_gff_5_U12 ( .A1(keyFF_keystate_gff_5_n61), .A2(
        keyFF_keystate_gff_5_n60), .ZN(keyFF_keystate_gff_5_n31) );
  NAND2_X1 keyFF_keystate_gff_5_U11 ( .A1(keyFF_keystate_gff_5_n67), .A2(
        keyFF_outputPar[13]), .ZN(keyFF_keystate_gff_5_n60) );
  MUX2_X1 keyFF_keystate_gff_5_U10 ( .A(keyFF_keystate_gff_5_n35), .B(
        keyFF_keystate_gff_5_n59), .S(keyFF_keystate_gff_5_n65), .Z(
        keyFF_keystate_gff_5_n61) );
  NAND2_X1 keyFF_keystate_gff_5_U9 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[17]), 
        .ZN(keyFF_keystate_gff_5_n59) );
  NAND2_X1 keyFF_keystate_gff_5_U8 ( .A1(keyFF_keystate_gff_5_n58), .A2(
        keyFF_keystate_gff_5_n57), .ZN(keyFF_keystate_gff_5_n32) );
  NAND2_X1 keyFF_keystate_gff_5_U7 ( .A1(keyFF_keystate_gff_5_n67), .A2(
        keyFF_outputPar[12]), .ZN(keyFF_keystate_gff_5_n57) );
  NOR2_X1 keyFF_keystate_gff_5_U6 ( .A1(ctrlData[0]), .A2(
        keyFF_keystate_gff_5_n56), .ZN(keyFF_keystate_gff_5_n67) );
  MUX2_X1 keyFF_keystate_gff_5_U5 ( .A(keyFF_keystate_gff_5_n36), .B(
        keyFF_keystate_gff_5_n55), .S(keyFF_keystate_gff_5_n65), .Z(
        keyFF_keystate_gff_5_n58) );
  INV_X1 keyFF_keystate_gff_5_U4 ( .A(keyFF_keystate_gff_5_n56), .ZN(
        keyFF_keystate_gff_5_n65) );
  INV_X1 keyFF_keystate_gff_5_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_5_n56) );
  NAND2_X1 keyFF_keystate_gff_5_U2 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[16]), 
        .ZN(keyFF_keystate_gff_5_n55) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_5_n32), .CK(clk), .Q(keyFF_outputPar[16]), .QN(
        keyFF_keystate_gff_5_n36) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_5_n31), .CK(clk), .Q(keyFF_outputPar[17]), .QN(
        keyFF_keystate_gff_5_n35) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_5_n30), .CK(clk), .Q(keyFF_outputPar[18]), .QN(
        keyFF_keystate_gff_5_n34) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_5_n29), .CK(clk), .Q(keyFF_outputPar[19]), .QN(
        keyFF_keystate_gff_5_n33) );
  NAND2_X1 keyFF_keystate_gff_6_U20 ( .A1(keyFF_keystate_gff_6_n68), .A2(
        keyFF_keystate_gff_6_n67), .ZN(keyFF_keystate_gff_6_n28) );
  NAND2_X1 keyFF_keystate_gff_6_U19 ( .A1(keyFF_keystate_gff_6_n66), .A2(
        keyFF_outputPar[19]), .ZN(keyFF_keystate_gff_6_n67) );
  MUX2_X1 keyFF_keystate_gff_6_U18 ( .A(keyFF_keystate_gff_6_n32), .B(
        keyFF_keystate_gff_6_n65), .S(keyFF_keystate_gff_6_n64), .Z(
        keyFF_keystate_gff_6_n68) );
  NAND2_X1 keyFF_keystate_gff_6_U17 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[23]), .ZN(keyFF_keystate_gff_6_n65) );
  NAND2_X1 keyFF_keystate_gff_6_U16 ( .A1(keyFF_keystate_gff_6_n63), .A2(
        keyFF_keystate_gff_6_n62), .ZN(keyFF_keystate_gff_6_n29) );
  NAND2_X1 keyFF_keystate_gff_6_U15 ( .A1(keyFF_keystate_gff_6_n66), .A2(
        keyFF_outputPar[18]), .ZN(keyFF_keystate_gff_6_n62) );
  MUX2_X1 keyFF_keystate_gff_6_U14 ( .A(keyFF_keystate_gff_6_n33), .B(
        keyFF_keystate_gff_6_n61), .S(keyFF_keystate_gff_6_n64), .Z(
        keyFF_keystate_gff_6_n63) );
  NAND2_X1 keyFF_keystate_gff_6_U13 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[22]), .ZN(keyFF_keystate_gff_6_n61) );
  NAND2_X1 keyFF_keystate_gff_6_U12 ( .A1(keyFF_keystate_gff_6_n60), .A2(
        keyFF_keystate_gff_6_n59), .ZN(keyFF_keystate_gff_6_n30) );
  NAND2_X1 keyFF_keystate_gff_6_U11 ( .A1(keyFF_keystate_gff_6_n66), .A2(
        keyFF_outputPar[17]), .ZN(keyFF_keystate_gff_6_n59) );
  MUX2_X1 keyFF_keystate_gff_6_U10 ( .A(keyFF_keystate_gff_6_n34), .B(
        keyFF_keystate_gff_6_n58), .S(keyFF_keystate_gff_6_n64), .Z(
        keyFF_keystate_gff_6_n60) );
  NAND2_X1 keyFF_keystate_gff_6_U9 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[21]), 
        .ZN(keyFF_keystate_gff_6_n58) );
  NAND2_X1 keyFF_keystate_gff_6_U8 ( .A1(keyFF_keystate_gff_6_n57), .A2(
        keyFF_keystate_gff_6_n56), .ZN(keyFF_keystate_gff_6_n31) );
  NAND2_X1 keyFF_keystate_gff_6_U7 ( .A1(keyFF_keystate_gff_6_n66), .A2(
        keyFF_outputPar[16]), .ZN(keyFF_keystate_gff_6_n56) );
  NOR2_X1 keyFF_keystate_gff_6_U6 ( .A1(ctrlData[0]), .A2(
        keyFF_keystate_gff_6_n55), .ZN(keyFF_keystate_gff_6_n66) );
  MUX2_X1 keyFF_keystate_gff_6_U5 ( .A(keyFF_keystate_gff_6_n35), .B(
        keyFF_keystate_gff_6_n54), .S(keyFF_keystate_gff_6_n64), .Z(
        keyFF_keystate_gff_6_n57) );
  INV_X1 keyFF_keystate_gff_6_U4 ( .A(keyFF_keystate_gff_6_n55), .ZN(
        keyFF_keystate_gff_6_n64) );
  INV_X1 keyFF_keystate_gff_6_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_6_n55) );
  NAND2_X1 keyFF_keystate_gff_6_U2 ( .A1(ctrlData[0]), .A2(keyFF_inputPar[20]), 
        .ZN(keyFF_keystate_gff_6_n54) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_6_n31), .CK(clk), .Q(keyFF_outputPar[20]), .QN(
        keyFF_keystate_gff_6_n35) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_6_n30), .CK(clk), .Q(keyFF_outputPar[21]), .QN(
        keyFF_keystate_gff_6_n34) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_6_n29), .CK(clk), .Q(keyFF_outputPar[22]), .QN(
        keyFF_keystate_gff_6_n33) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_6_n28), .CK(clk), .Q(keyFF_outputPar[23]), .QN(
        keyFF_keystate_gff_6_n32) );
  NAND2_X1 keyFF_keystate_gff_7_U20 ( .A1(keyFF_keystate_gff_7_n68), .A2(
        keyFF_keystate_gff_7_n67), .ZN(keyFF_keystate_gff_7_n28) );
  NAND2_X1 keyFF_keystate_gff_7_U19 ( .A1(keyFF_keystate_gff_7_n66), .A2(
        keyFF_outputPar[23]), .ZN(keyFF_keystate_gff_7_n67) );
  MUX2_X1 keyFF_keystate_gff_7_U18 ( .A(keyFF_keystate_gff_7_n32), .B(
        keyFF_keystate_gff_7_n65), .S(keyFF_keystate_gff_7_n64), .Z(
        keyFF_keystate_gff_7_n68) );
  NAND2_X1 keyFF_keystate_gff_7_U17 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[27]), .ZN(keyFF_keystate_gff_7_n65) );
  NAND2_X1 keyFF_keystate_gff_7_U16 ( .A1(keyFF_keystate_gff_7_n63), .A2(
        keyFF_keystate_gff_7_n62), .ZN(keyFF_keystate_gff_7_n29) );
  NAND2_X1 keyFF_keystate_gff_7_U15 ( .A1(keyFF_keystate_gff_7_n66), .A2(
        keyFF_outputPar[22]), .ZN(keyFF_keystate_gff_7_n62) );
  MUX2_X1 keyFF_keystate_gff_7_U14 ( .A(keyFF_keystate_gff_7_n33), .B(
        keyFF_keystate_gff_7_n61), .S(keyFF_keystate_gff_7_n64), .Z(
        keyFF_keystate_gff_7_n63) );
  NAND2_X1 keyFF_keystate_gff_7_U13 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[26]), .ZN(keyFF_keystate_gff_7_n61) );
  NAND2_X1 keyFF_keystate_gff_7_U12 ( .A1(keyFF_keystate_gff_7_n60), .A2(
        keyFF_keystate_gff_7_n59), .ZN(keyFF_keystate_gff_7_n30) );
  NAND2_X1 keyFF_keystate_gff_7_U11 ( .A1(keyFF_keystate_gff_7_n66), .A2(
        keyFF_outputPar[21]), .ZN(keyFF_keystate_gff_7_n59) );
  MUX2_X1 keyFF_keystate_gff_7_U10 ( .A(keyFF_keystate_gff_7_n34), .B(
        keyFF_keystate_gff_7_n58), .S(keyFF_keystate_gff_7_n64), .Z(
        keyFF_keystate_gff_7_n60) );
  NAND2_X1 keyFF_keystate_gff_7_U9 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[25]), .ZN(keyFF_keystate_gff_7_n58) );
  NAND2_X1 keyFF_keystate_gff_7_U8 ( .A1(keyFF_keystate_gff_7_n57), .A2(
        keyFF_keystate_gff_7_n56), .ZN(keyFF_keystate_gff_7_n31) );
  NAND2_X1 keyFF_keystate_gff_7_U7 ( .A1(keyFF_keystate_gff_7_n66), .A2(
        keyFF_outputPar[20]), .ZN(keyFF_keystate_gff_7_n56) );
  NOR2_X1 keyFF_keystate_gff_7_U6 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_keystate_gff_7_n55), .ZN(keyFF_keystate_gff_7_n66) );
  MUX2_X1 keyFF_keystate_gff_7_U5 ( .A(keyFF_keystate_gff_7_n35), .B(
        keyFF_keystate_gff_7_n54), .S(keyFF_keystate_gff_7_n64), .Z(
        keyFF_keystate_gff_7_n57) );
  INV_X1 keyFF_keystate_gff_7_U4 ( .A(keyFF_keystate_gff_7_n55), .ZN(
        keyFF_keystate_gff_7_n64) );
  INV_X1 keyFF_keystate_gff_7_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_7_n55) );
  NAND2_X1 keyFF_keystate_gff_7_U2 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[24]), .ZN(keyFF_keystate_gff_7_n54) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_7_n31), .CK(clk), .Q(keyFF_outputPar[24]), .QN(
        keyFF_keystate_gff_7_n35) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_7_n30), .CK(clk), .Q(keyFF_outputPar[25]), .QN(
        keyFF_keystate_gff_7_n34) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_7_n29), .CK(clk), .Q(keyFF_outputPar[26]), .QN(
        keyFF_keystate_gff_7_n33) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_7_n28), .CK(clk), .Q(keyFF_outputPar[27]), .QN(
        keyFF_keystate_gff_7_n32) );
  NAND2_X1 keyFF_keystate_gff_8_U20 ( .A1(keyFF_keystate_gff_8_n68), .A2(
        keyFF_keystate_gff_8_n67), .ZN(keyFF_keystate_gff_8_n28) );
  NAND2_X1 keyFF_keystate_gff_8_U19 ( .A1(keyFF_keystate_gff_8_n66), .A2(
        keyFF_outputPar[27]), .ZN(keyFF_keystate_gff_8_n67) );
  MUX2_X1 keyFF_keystate_gff_8_U18 ( .A(keyFF_keystate_gff_8_n32), .B(
        keyFF_keystate_gff_8_n65), .S(keyFF_keystate_gff_8_n64), .Z(
        keyFF_keystate_gff_8_n68) );
  NAND2_X1 keyFF_keystate_gff_8_U17 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[31]), .ZN(keyFF_keystate_gff_8_n65) );
  NAND2_X1 keyFF_keystate_gff_8_U16 ( .A1(keyFF_keystate_gff_8_n63), .A2(
        keyFF_keystate_gff_8_n62), .ZN(keyFF_keystate_gff_8_n29) );
  NAND2_X1 keyFF_keystate_gff_8_U15 ( .A1(keyFF_keystate_gff_8_n66), .A2(
        keyFF_outputPar[26]), .ZN(keyFF_keystate_gff_8_n62) );
  MUX2_X1 keyFF_keystate_gff_8_U14 ( .A(keyFF_keystate_gff_8_n33), .B(
        keyFF_keystate_gff_8_n61), .S(keyFF_keystate_gff_8_n64), .Z(
        keyFF_keystate_gff_8_n63) );
  NAND2_X1 keyFF_keystate_gff_8_U13 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[30]), .ZN(keyFF_keystate_gff_8_n61) );
  NAND2_X1 keyFF_keystate_gff_8_U12 ( .A1(keyFF_keystate_gff_8_n60), .A2(
        keyFF_keystate_gff_8_n59), .ZN(keyFF_keystate_gff_8_n30) );
  NAND2_X1 keyFF_keystate_gff_8_U11 ( .A1(keyFF_keystate_gff_8_n66), .A2(
        keyFF_outputPar[25]), .ZN(keyFF_keystate_gff_8_n59) );
  MUX2_X1 keyFF_keystate_gff_8_U10 ( .A(keyFF_keystate_gff_8_n34), .B(
        keyFF_keystate_gff_8_n58), .S(keyFF_keystate_gff_8_n64), .Z(
        keyFF_keystate_gff_8_n60) );
  NAND2_X1 keyFF_keystate_gff_8_U9 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[29]), .ZN(keyFF_keystate_gff_8_n58) );
  NAND2_X1 keyFF_keystate_gff_8_U8 ( .A1(keyFF_keystate_gff_8_n57), .A2(
        keyFF_keystate_gff_8_n56), .ZN(keyFF_keystate_gff_8_n31) );
  NAND2_X1 keyFF_keystate_gff_8_U7 ( .A1(keyFF_keystate_gff_8_n66), .A2(
        keyFF_outputPar[24]), .ZN(keyFF_keystate_gff_8_n56) );
  NOR2_X1 keyFF_keystate_gff_8_U6 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_keystate_gff_8_n55), .ZN(keyFF_keystate_gff_8_n66) );
  MUX2_X1 keyFF_keystate_gff_8_U5 ( .A(keyFF_keystate_gff_8_n35), .B(
        keyFF_keystate_gff_8_n54), .S(keyFF_keystate_gff_8_n64), .Z(
        keyFF_keystate_gff_8_n57) );
  INV_X1 keyFF_keystate_gff_8_U4 ( .A(keyFF_keystate_gff_8_n55), .ZN(
        keyFF_keystate_gff_8_n64) );
  INV_X1 keyFF_keystate_gff_8_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_8_n55) );
  NAND2_X1 keyFF_keystate_gff_8_U2 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[28]), .ZN(keyFF_keystate_gff_8_n54) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_8_n31), .CK(clk), .Q(keyFF_outputPar[28]), .QN(
        keyFF_keystate_gff_8_n35) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_8_n30), .CK(clk), .Q(keyFF_outputPar[29]), .QN(
        keyFF_keystate_gff_8_n34) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_8_n29), .CK(clk), .Q(keyFF_outputPar[30]), .QN(
        keyFF_keystate_gff_8_n33) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_8_n28), .CK(clk), .Q(keyFF_outputPar[31]), .QN(
        keyFF_keystate_gff_8_n32) );
  NAND2_X1 keyFF_keystate_gff_9_U20 ( .A1(keyFF_keystate_gff_9_n69), .A2(
        keyFF_keystate_gff_9_n68), .ZN(keyFF_keystate_gff_9_n29) );
  NAND2_X1 keyFF_keystate_gff_9_U19 ( .A1(keyFF_keystate_gff_9_n67), .A2(
        keyFF_outputPar[31]), .ZN(keyFF_keystate_gff_9_n68) );
  MUX2_X1 keyFF_keystate_gff_9_U18 ( .A(keyFF_keystate_gff_9_n33), .B(
        keyFF_keystate_gff_9_n66), .S(keyFF_keystate_gff_9_n65), .Z(
        keyFF_keystate_gff_9_n69) );
  NAND2_X1 keyFF_keystate_gff_9_U17 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[35]), .ZN(keyFF_keystate_gff_9_n66) );
  NAND2_X1 keyFF_keystate_gff_9_U16 ( .A1(keyFF_keystate_gff_9_n64), .A2(
        keyFF_keystate_gff_9_n63), .ZN(keyFF_keystate_gff_9_n30) );
  NAND2_X1 keyFF_keystate_gff_9_U15 ( .A1(keyFF_keystate_gff_9_n67), .A2(
        keyFF_outputPar[30]), .ZN(keyFF_keystate_gff_9_n63) );
  MUX2_X1 keyFF_keystate_gff_9_U14 ( .A(keyFF_keystate_gff_9_n34), .B(
        keyFF_keystate_gff_9_n62), .S(keyFF_keystate_gff_9_n65), .Z(
        keyFF_keystate_gff_9_n64) );
  NAND2_X1 keyFF_keystate_gff_9_U13 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[34]), .ZN(keyFF_keystate_gff_9_n62) );
  NAND2_X1 keyFF_keystate_gff_9_U12 ( .A1(keyFF_keystate_gff_9_n61), .A2(
        keyFF_keystate_gff_9_n60), .ZN(keyFF_keystate_gff_9_n31) );
  NAND2_X1 keyFF_keystate_gff_9_U11 ( .A1(keyFF_keystate_gff_9_n67), .A2(
        keyFF_outputPar[29]), .ZN(keyFF_keystate_gff_9_n60) );
  MUX2_X1 keyFF_keystate_gff_9_U10 ( .A(keyFF_keystate_gff_9_n35), .B(
        keyFF_keystate_gff_9_n59), .S(keyFF_keystate_gff_9_n65), .Z(
        keyFF_keystate_gff_9_n61) );
  NAND2_X1 keyFF_keystate_gff_9_U9 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[33]), .ZN(keyFF_keystate_gff_9_n59) );
  NAND2_X1 keyFF_keystate_gff_9_U8 ( .A1(keyFF_keystate_gff_9_n58), .A2(
        keyFF_keystate_gff_9_n57), .ZN(keyFF_keystate_gff_9_n32) );
  NAND2_X1 keyFF_keystate_gff_9_U7 ( .A1(keyFF_keystate_gff_9_n67), .A2(
        keyFF_outputPar[28]), .ZN(keyFF_keystate_gff_9_n57) );
  NOR2_X1 keyFF_keystate_gff_9_U6 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_keystate_gff_9_n56), .ZN(keyFF_keystate_gff_9_n67) );
  MUX2_X1 keyFF_keystate_gff_9_U5 ( .A(keyFF_keystate_gff_9_n36), .B(
        keyFF_keystate_gff_9_n55), .S(keyFF_keystate_gff_9_n65), .Z(
        keyFF_keystate_gff_9_n58) );
  INV_X1 keyFF_keystate_gff_9_U4 ( .A(keyFF_keystate_gff_9_n56), .ZN(
        keyFF_keystate_gff_9_n65) );
  INV_X1 keyFF_keystate_gff_9_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_9_n56) );
  NAND2_X1 keyFF_keystate_gff_9_U2 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[32]), .ZN(keyFF_keystate_gff_9_n55) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_9_n32), .CK(clk), .Q(keyFF_outputPar[32]), .QN(
        keyFF_keystate_gff_9_n36) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_9_n31), .CK(clk), .Q(keyFF_outputPar[33]), .QN(
        keyFF_keystate_gff_9_n35) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_9_n30), .CK(clk), .Q(keyFF_outputPar[34]), .QN(
        keyFF_keystate_gff_9_n34) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_9_n29), .CK(clk), .Q(keyFF_outputPar[35]), .QN(
        keyFF_keystate_gff_9_n33) );
  NAND2_X1 keyFF_keystate_gff_10_U20 ( .A1(keyFF_keystate_gff_10_n69), .A2(
        keyFF_keystate_gff_10_n68), .ZN(keyFF_keystate_gff_10_n29) );
  NAND2_X1 keyFF_keystate_gff_10_U19 ( .A1(keyFF_keystate_gff_10_n67), .A2(
        keyFF_outputPar[35]), .ZN(keyFF_keystate_gff_10_n68) );
  MUX2_X1 keyFF_keystate_gff_10_U18 ( .A(keyFF_keystate_gff_10_n33), .B(
        keyFF_keystate_gff_10_n66), .S(keyFF_keystate_gff_10_n65), .Z(
        keyFF_keystate_gff_10_n69) );
  NAND2_X1 keyFF_keystate_gff_10_U17 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[39]), .ZN(keyFF_keystate_gff_10_n66) );
  NAND2_X1 keyFF_keystate_gff_10_U16 ( .A1(keyFF_keystate_gff_10_n64), .A2(
        keyFF_keystate_gff_10_n63), .ZN(keyFF_keystate_gff_10_n30) );
  NAND2_X1 keyFF_keystate_gff_10_U15 ( .A1(keyFF_keystate_gff_10_n67), .A2(
        keyFF_outputPar[34]), .ZN(keyFF_keystate_gff_10_n63) );
  MUX2_X1 keyFF_keystate_gff_10_U14 ( .A(keyFF_keystate_gff_10_n34), .B(
        keyFF_keystate_gff_10_n62), .S(keyFF_keystate_gff_10_n65), .Z(
        keyFF_keystate_gff_10_n64) );
  NAND2_X1 keyFF_keystate_gff_10_U13 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[38]), .ZN(keyFF_keystate_gff_10_n62) );
  NAND2_X1 keyFF_keystate_gff_10_U12 ( .A1(keyFF_keystate_gff_10_n61), .A2(
        keyFF_keystate_gff_10_n60), .ZN(keyFF_keystate_gff_10_n31) );
  NAND2_X1 keyFF_keystate_gff_10_U11 ( .A1(keyFF_keystate_gff_10_n67), .A2(
        keyFF_outputPar[33]), .ZN(keyFF_keystate_gff_10_n60) );
  MUX2_X1 keyFF_keystate_gff_10_U10 ( .A(keyFF_keystate_gff_10_n35), .B(
        keyFF_keystate_gff_10_n59), .S(keyFF_keystate_gff_10_n65), .Z(
        keyFF_keystate_gff_10_n61) );
  NAND2_X1 keyFF_keystate_gff_10_U9 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[37]), .ZN(keyFF_keystate_gff_10_n59) );
  NAND2_X1 keyFF_keystate_gff_10_U8 ( .A1(keyFF_keystate_gff_10_n58), .A2(
        keyFF_keystate_gff_10_n57), .ZN(keyFF_keystate_gff_10_n32) );
  NAND2_X1 keyFF_keystate_gff_10_U7 ( .A1(keyFF_keystate_gff_10_n67), .A2(
        keyFF_outputPar[32]), .ZN(keyFF_keystate_gff_10_n57) );
  NOR2_X1 keyFF_keystate_gff_10_U6 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_keystate_gff_10_n56), .ZN(keyFF_keystate_gff_10_n67) );
  MUX2_X1 keyFF_keystate_gff_10_U5 ( .A(keyFF_keystate_gff_10_n36), .B(
        keyFF_keystate_gff_10_n55), .S(keyFF_keystate_gff_10_n65), .Z(
        keyFF_keystate_gff_10_n58) );
  INV_X1 keyFF_keystate_gff_10_U4 ( .A(keyFF_keystate_gff_10_n56), .ZN(
        keyFF_keystate_gff_10_n65) );
  INV_X1 keyFF_keystate_gff_10_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_10_n56) );
  NAND2_X1 keyFF_keystate_gff_10_U2 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[36]), .ZN(keyFF_keystate_gff_10_n55) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_10_n32), .CK(clk), .Q(keyFF_outputPar[36]), .QN(
        keyFF_keystate_gff_10_n36) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_10_n31), .CK(clk), .Q(keyFF_outputPar[37]), .QN(
        keyFF_keystate_gff_10_n35) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_10_n30), .CK(clk), .Q(keyFF_outputPar[38]), .QN(
        keyFF_keystate_gff_10_n34) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_10_n29), .CK(clk), .Q(keyFF_outputPar[39]), .QN(
        keyFF_keystate_gff_10_n33) );
  NAND2_X1 keyFF_keystate_gff_11_U20 ( .A1(keyFF_keystate_gff_11_n69), .A2(
        keyFF_keystate_gff_11_n68), .ZN(keyFF_keystate_gff_11_n29) );
  NAND2_X1 keyFF_keystate_gff_11_U19 ( .A1(keyFF_keystate_gff_11_n67), .A2(
        keyFF_outputPar[39]), .ZN(keyFF_keystate_gff_11_n68) );
  MUX2_X1 keyFF_keystate_gff_11_U18 ( .A(keyFF_keystate_gff_11_n33), .B(
        keyFF_keystate_gff_11_n66), .S(keyFF_keystate_gff_11_n65), .Z(
        keyFF_keystate_gff_11_n69) );
  NAND2_X1 keyFF_keystate_gff_11_U17 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[43]), .ZN(keyFF_keystate_gff_11_n66) );
  NAND2_X1 keyFF_keystate_gff_11_U16 ( .A1(keyFF_keystate_gff_11_n64), .A2(
        keyFF_keystate_gff_11_n63), .ZN(keyFF_keystate_gff_11_n30) );
  NAND2_X1 keyFF_keystate_gff_11_U15 ( .A1(keyFF_keystate_gff_11_n67), .A2(
        keyFF_outputPar[38]), .ZN(keyFF_keystate_gff_11_n63) );
  MUX2_X1 keyFF_keystate_gff_11_U14 ( .A(keyFF_keystate_gff_11_n34), .B(
        keyFF_keystate_gff_11_n62), .S(keyFF_keystate_gff_11_n65), .Z(
        keyFF_keystate_gff_11_n64) );
  NAND2_X1 keyFF_keystate_gff_11_U13 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[42]), .ZN(keyFF_keystate_gff_11_n62) );
  NAND2_X1 keyFF_keystate_gff_11_U12 ( .A1(keyFF_keystate_gff_11_n61), .A2(
        keyFF_keystate_gff_11_n60), .ZN(keyFF_keystate_gff_11_n31) );
  NAND2_X1 keyFF_keystate_gff_11_U11 ( .A1(keyFF_keystate_gff_11_n67), .A2(
        keyFF_outputPar[37]), .ZN(keyFF_keystate_gff_11_n60) );
  MUX2_X1 keyFF_keystate_gff_11_U10 ( .A(keyFF_keystate_gff_11_n35), .B(
        keyFF_keystate_gff_11_n59), .S(keyFF_keystate_gff_11_n65), .Z(
        keyFF_keystate_gff_11_n61) );
  NAND2_X1 keyFF_keystate_gff_11_U9 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[41]), .ZN(keyFF_keystate_gff_11_n59) );
  NAND2_X1 keyFF_keystate_gff_11_U8 ( .A1(keyFF_keystate_gff_11_n58), .A2(
        keyFF_keystate_gff_11_n57), .ZN(keyFF_keystate_gff_11_n32) );
  NAND2_X1 keyFF_keystate_gff_11_U7 ( .A1(keyFF_keystate_gff_11_n67), .A2(
        keyFF_outputPar[36]), .ZN(keyFF_keystate_gff_11_n57) );
  NOR2_X1 keyFF_keystate_gff_11_U6 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_keystate_gff_11_n56), .ZN(keyFF_keystate_gff_11_n67) );
  MUX2_X1 keyFF_keystate_gff_11_U5 ( .A(keyFF_keystate_gff_11_n36), .B(
        keyFF_keystate_gff_11_n55), .S(keyFF_keystate_gff_11_n65), .Z(
        keyFF_keystate_gff_11_n58) );
  INV_X1 keyFF_keystate_gff_11_U4 ( .A(keyFF_keystate_gff_11_n56), .ZN(
        keyFF_keystate_gff_11_n65) );
  INV_X1 keyFF_keystate_gff_11_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_11_n56) );
  NAND2_X1 keyFF_keystate_gff_11_U2 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[40]), .ZN(keyFF_keystate_gff_11_n55) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_11_n32), .CK(clk), .Q(keyFF_outputPar[40]), .QN(
        keyFF_keystate_gff_11_n36) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_11_n31), .CK(clk), .Q(keyFF_outputPar[41]), .QN(
        keyFF_keystate_gff_11_n35) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_11_n30), .CK(clk), .Q(keyFF_outputPar[42]), .QN(
        keyFF_keystate_gff_11_n34) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_11_n29), .CK(clk), .Q(keyFF_outputPar[43]), .QN(
        keyFF_keystate_gff_11_n33) );
  NAND2_X1 keyFF_keystate_gff_12_U20 ( .A1(keyFF_keystate_gff_12_n69), .A2(
        keyFF_keystate_gff_12_n68), .ZN(keyFF_keystate_gff_12_n29) );
  NAND2_X1 keyFF_keystate_gff_12_U19 ( .A1(keyFF_keystate_gff_12_n67), .A2(
        keyFF_outputPar[43]), .ZN(keyFF_keystate_gff_12_n68) );
  MUX2_X1 keyFF_keystate_gff_12_U18 ( .A(keyFF_keystate_gff_12_n33), .B(
        keyFF_keystate_gff_12_n66), .S(keyFF_keystate_gff_12_n65), .Z(
        keyFF_keystate_gff_12_n69) );
  NAND2_X1 keyFF_keystate_gff_12_U17 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[47]), .ZN(keyFF_keystate_gff_12_n66) );
  NAND2_X1 keyFF_keystate_gff_12_U16 ( .A1(keyFF_keystate_gff_12_n64), .A2(
        keyFF_keystate_gff_12_n63), .ZN(keyFF_keystate_gff_12_n30) );
  NAND2_X1 keyFF_keystate_gff_12_U15 ( .A1(keyFF_keystate_gff_12_n67), .A2(
        keyFF_outputPar[42]), .ZN(keyFF_keystate_gff_12_n63) );
  MUX2_X1 keyFF_keystate_gff_12_U14 ( .A(keyFF_keystate_gff_12_n34), .B(
        keyFF_keystate_gff_12_n62), .S(keyFF_keystate_gff_12_n65), .Z(
        keyFF_keystate_gff_12_n64) );
  NAND2_X1 keyFF_keystate_gff_12_U13 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[46]), .ZN(keyFF_keystate_gff_12_n62) );
  NAND2_X1 keyFF_keystate_gff_12_U12 ( .A1(keyFF_keystate_gff_12_n61), .A2(
        keyFF_keystate_gff_12_n60), .ZN(keyFF_keystate_gff_12_n31) );
  NAND2_X1 keyFF_keystate_gff_12_U11 ( .A1(keyFF_keystate_gff_12_n67), .A2(
        keyFF_outputPar[41]), .ZN(keyFF_keystate_gff_12_n60) );
  MUX2_X1 keyFF_keystate_gff_12_U10 ( .A(keyFF_keystate_gff_12_n35), .B(
        keyFF_keystate_gff_12_n59), .S(keyFF_keystate_gff_12_n65), .Z(
        keyFF_keystate_gff_12_n61) );
  NAND2_X1 keyFF_keystate_gff_12_U9 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[45]), .ZN(keyFF_keystate_gff_12_n59) );
  NAND2_X1 keyFF_keystate_gff_12_U8 ( .A1(keyFF_keystate_gff_12_n58), .A2(
        keyFF_keystate_gff_12_n57), .ZN(keyFF_keystate_gff_12_n32) );
  NAND2_X1 keyFF_keystate_gff_12_U7 ( .A1(keyFF_keystate_gff_12_n67), .A2(
        keyFF_outputPar[40]), .ZN(keyFF_keystate_gff_12_n57) );
  NOR2_X1 keyFF_keystate_gff_12_U6 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_keystate_gff_12_n56), .ZN(keyFF_keystate_gff_12_n67) );
  MUX2_X1 keyFF_keystate_gff_12_U5 ( .A(keyFF_keystate_gff_12_n36), .B(
        keyFF_keystate_gff_12_n55), .S(keyFF_keystate_gff_12_n65), .Z(
        keyFF_keystate_gff_12_n58) );
  INV_X1 keyFF_keystate_gff_12_U4 ( .A(keyFF_keystate_gff_12_n56), .ZN(
        keyFF_keystate_gff_12_n65) );
  INV_X1 keyFF_keystate_gff_12_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_12_n56) );
  NAND2_X1 keyFF_keystate_gff_12_U2 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[44]), .ZN(keyFF_keystate_gff_12_n55) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_12_n32), .CK(clk), .Q(keyFF_outputPar[44]), .QN(
        keyFF_keystate_gff_12_n36) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_12_n31), .CK(clk), .Q(keyFF_outputPar[45]), .QN(
        keyFF_keystate_gff_12_n35) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_12_n30), .CK(clk), .Q(keyFF_outputPar[46]), .QN(
        keyFF_keystate_gff_12_n34) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_12_n29), .CK(clk), .Q(keyFF_outputPar[47]), .QN(
        keyFF_keystate_gff_12_n33) );
  NAND2_X1 keyFF_keystate_gff_13_U20 ( .A1(keyFF_keystate_gff_13_n69), .A2(
        keyFF_keystate_gff_13_n68), .ZN(keyFF_keystate_gff_13_n29) );
  NAND2_X1 keyFF_keystate_gff_13_U19 ( .A1(keyFF_keystate_gff_13_n67), .A2(
        keyFF_outputPar[47]), .ZN(keyFF_keystate_gff_13_n68) );
  MUX2_X1 keyFF_keystate_gff_13_U18 ( .A(keyFF_keystate_gff_13_n33), .B(
        keyFF_keystate_gff_13_n66), .S(keyFF_keystate_gff_13_n65), .Z(
        keyFF_keystate_gff_13_n69) );
  NAND2_X1 keyFF_keystate_gff_13_U17 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[51]), .ZN(keyFF_keystate_gff_13_n66) );
  NAND2_X1 keyFF_keystate_gff_13_U16 ( .A1(keyFF_keystate_gff_13_n64), .A2(
        keyFF_keystate_gff_13_n63), .ZN(keyFF_keystate_gff_13_n30) );
  NAND2_X1 keyFF_keystate_gff_13_U15 ( .A1(keyFF_keystate_gff_13_n67), .A2(
        keyFF_outputPar[46]), .ZN(keyFF_keystate_gff_13_n63) );
  MUX2_X1 keyFF_keystate_gff_13_U14 ( .A(keyFF_keystate_gff_13_n34), .B(
        keyFF_keystate_gff_13_n62), .S(keyFF_keystate_gff_13_n65), .Z(
        keyFF_keystate_gff_13_n64) );
  NAND2_X1 keyFF_keystate_gff_13_U13 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[50]), .ZN(keyFF_keystate_gff_13_n62) );
  NAND2_X1 keyFF_keystate_gff_13_U12 ( .A1(keyFF_keystate_gff_13_n61), .A2(
        keyFF_keystate_gff_13_n60), .ZN(keyFF_keystate_gff_13_n31) );
  NAND2_X1 keyFF_keystate_gff_13_U11 ( .A1(keyFF_keystate_gff_13_n67), .A2(
        keyFF_outputPar[45]), .ZN(keyFF_keystate_gff_13_n60) );
  MUX2_X1 keyFF_keystate_gff_13_U10 ( .A(keyFF_keystate_gff_13_n35), .B(
        keyFF_keystate_gff_13_n59), .S(keyFF_keystate_gff_13_n65), .Z(
        keyFF_keystate_gff_13_n61) );
  NAND2_X1 keyFF_keystate_gff_13_U9 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[49]), .ZN(keyFF_keystate_gff_13_n59) );
  NAND2_X1 keyFF_keystate_gff_13_U8 ( .A1(keyFF_keystate_gff_13_n58), .A2(
        keyFF_keystate_gff_13_n57), .ZN(keyFF_keystate_gff_13_n32) );
  NAND2_X1 keyFF_keystate_gff_13_U7 ( .A1(keyFF_keystate_gff_13_n67), .A2(
        keyFF_outputPar[44]), .ZN(keyFF_keystate_gff_13_n57) );
  NOR2_X1 keyFF_keystate_gff_13_U6 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_keystate_gff_13_n56), .ZN(keyFF_keystate_gff_13_n67) );
  MUX2_X1 keyFF_keystate_gff_13_U5 ( .A(keyFF_keystate_gff_13_n36), .B(
        keyFF_keystate_gff_13_n55), .S(keyFF_keystate_gff_13_n65), .Z(
        keyFF_keystate_gff_13_n58) );
  INV_X1 keyFF_keystate_gff_13_U4 ( .A(keyFF_keystate_gff_13_n56), .ZN(
        keyFF_keystate_gff_13_n65) );
  INV_X1 keyFF_keystate_gff_13_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_13_n56) );
  NAND2_X1 keyFF_keystate_gff_13_U2 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[48]), .ZN(keyFF_keystate_gff_13_n55) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_13_n32), .CK(clk), .Q(keyFF_outputPar[48]), .QN(
        keyFF_keystate_gff_13_n36) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_13_n31), .CK(clk), .Q(keyFF_outputPar[49]), .QN(
        keyFF_keystate_gff_13_n35) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_13_n30), .CK(clk), .Q(keyFF_outputPar[50]), .QN(
        keyFF_keystate_gff_13_n34) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_13_n29), .CK(clk), .Q(keyFF_outputPar[51]), .QN(
        keyFF_keystate_gff_13_n33) );
  NAND2_X1 keyFF_keystate_gff_14_U20 ( .A1(keyFF_keystate_gff_14_n69), .A2(
        keyFF_keystate_gff_14_n68), .ZN(keyFF_keystate_gff_14_n29) );
  NAND2_X1 keyFF_keystate_gff_14_U19 ( .A1(keyFF_keystate_gff_14_n67), .A2(
        keyFF_outputPar[51]), .ZN(keyFF_keystate_gff_14_n68) );
  MUX2_X1 keyFF_keystate_gff_14_U18 ( .A(keyFF_keystate_gff_14_n33), .B(
        keyFF_keystate_gff_14_n66), .S(keyFF_keystate_gff_14_n65), .Z(
        keyFF_keystate_gff_14_n69) );
  NAND2_X1 keyFF_keystate_gff_14_U17 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[55]), .ZN(keyFF_keystate_gff_14_n66) );
  NAND2_X1 keyFF_keystate_gff_14_U16 ( .A1(keyFF_keystate_gff_14_n64), .A2(
        keyFF_keystate_gff_14_n63), .ZN(keyFF_keystate_gff_14_n30) );
  NAND2_X1 keyFF_keystate_gff_14_U15 ( .A1(keyFF_keystate_gff_14_n67), .A2(
        keyFF_outputPar[50]), .ZN(keyFF_keystate_gff_14_n63) );
  MUX2_X1 keyFF_keystate_gff_14_U14 ( .A(keyFF_keystate_gff_14_n34), .B(
        keyFF_keystate_gff_14_n62), .S(keyFF_keystate_gff_14_n65), .Z(
        keyFF_keystate_gff_14_n64) );
  NAND2_X1 keyFF_keystate_gff_14_U13 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[54]), .ZN(keyFF_keystate_gff_14_n62) );
  NAND2_X1 keyFF_keystate_gff_14_U12 ( .A1(keyFF_keystate_gff_14_n61), .A2(
        keyFF_keystate_gff_14_n60), .ZN(keyFF_keystate_gff_14_n31) );
  NAND2_X1 keyFF_keystate_gff_14_U11 ( .A1(keyFF_keystate_gff_14_n67), .A2(
        keyFF_outputPar[49]), .ZN(keyFF_keystate_gff_14_n60) );
  MUX2_X1 keyFF_keystate_gff_14_U10 ( .A(keyFF_keystate_gff_14_n35), .B(
        keyFF_keystate_gff_14_n59), .S(keyFF_keystate_gff_14_n65), .Z(
        keyFF_keystate_gff_14_n61) );
  NAND2_X1 keyFF_keystate_gff_14_U9 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[53]), .ZN(keyFF_keystate_gff_14_n59) );
  NAND2_X1 keyFF_keystate_gff_14_U8 ( .A1(keyFF_keystate_gff_14_n58), .A2(
        keyFF_keystate_gff_14_n57), .ZN(keyFF_keystate_gff_14_n32) );
  NAND2_X1 keyFF_keystate_gff_14_U7 ( .A1(keyFF_keystate_gff_14_n67), .A2(
        keyFF_outputPar[48]), .ZN(keyFF_keystate_gff_14_n57) );
  NOR2_X1 keyFF_keystate_gff_14_U6 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_keystate_gff_14_n56), .ZN(keyFF_keystate_gff_14_n67) );
  MUX2_X1 keyFF_keystate_gff_14_U5 ( .A(keyFF_keystate_gff_14_n36), .B(
        keyFF_keystate_gff_14_n55), .S(keyFF_keystate_gff_14_n65), .Z(
        keyFF_keystate_gff_14_n58) );
  INV_X1 keyFF_keystate_gff_14_U4 ( .A(keyFF_keystate_gff_14_n56), .ZN(
        keyFF_keystate_gff_14_n65) );
  INV_X1 keyFF_keystate_gff_14_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_14_n56) );
  NAND2_X1 keyFF_keystate_gff_14_U2 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[52]), .ZN(keyFF_keystate_gff_14_n55) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_14_n32), .CK(clk), .Q(keyFF_outputPar[52]), .QN(
        keyFF_keystate_gff_14_n36) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_14_n31), .CK(clk), .Q(keyFF_outputPar[53]), .QN(
        keyFF_keystate_gff_14_n35) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_14_n30), .CK(clk), .Q(keyFF_outputPar[54]), .QN(
        keyFF_keystate_gff_14_n34) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_14_n29), .CK(clk), .Q(keyFF_outputPar[55]), .QN(
        keyFF_keystate_gff_14_n33) );
  NAND2_X1 keyFF_keystate_gff_15_U20 ( .A1(keyFF_keystate_gff_15_n69), .A2(
        keyFF_keystate_gff_15_n68), .ZN(keyFF_keystate_gff_15_n29) );
  NAND2_X1 keyFF_keystate_gff_15_U19 ( .A1(keyFF_keystate_gff_15_n67), .A2(
        keyFF_outputPar[55]), .ZN(keyFF_keystate_gff_15_n68) );
  MUX2_X1 keyFF_keystate_gff_15_U18 ( .A(keyFF_keystate_gff_15_n33), .B(
        keyFF_keystate_gff_15_n66), .S(keyFF_keystate_gff_15_n65), .Z(
        keyFF_keystate_gff_15_n69) );
  NAND2_X1 keyFF_keystate_gff_15_U17 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[59]), .ZN(keyFF_keystate_gff_15_n66) );
  NAND2_X1 keyFF_keystate_gff_15_U16 ( .A1(keyFF_keystate_gff_15_n64), .A2(
        keyFF_keystate_gff_15_n63), .ZN(keyFF_keystate_gff_15_n30) );
  NAND2_X1 keyFF_keystate_gff_15_U15 ( .A1(keyFF_keystate_gff_15_n67), .A2(
        keyFF_outputPar[54]), .ZN(keyFF_keystate_gff_15_n63) );
  MUX2_X1 keyFF_keystate_gff_15_U14 ( .A(keyFF_keystate_gff_15_n34), .B(
        keyFF_keystate_gff_15_n62), .S(keyFF_keystate_gff_15_n65), .Z(
        keyFF_keystate_gff_15_n64) );
  NAND2_X1 keyFF_keystate_gff_15_U13 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[58]), .ZN(keyFF_keystate_gff_15_n62) );
  NAND2_X1 keyFF_keystate_gff_15_U12 ( .A1(keyFF_keystate_gff_15_n61), .A2(
        keyFF_keystate_gff_15_n60), .ZN(keyFF_keystate_gff_15_n31) );
  NAND2_X1 keyFF_keystate_gff_15_U11 ( .A1(keyFF_keystate_gff_15_n67), .A2(
        keyFF_outputPar[53]), .ZN(keyFF_keystate_gff_15_n60) );
  MUX2_X1 keyFF_keystate_gff_15_U10 ( .A(keyFF_keystate_gff_15_n35), .B(
        keyFF_keystate_gff_15_n59), .S(keyFF_keystate_gff_15_n65), .Z(
        keyFF_keystate_gff_15_n61) );
  NAND2_X1 keyFF_keystate_gff_15_U9 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[57]), .ZN(keyFF_keystate_gff_15_n59) );
  NAND2_X1 keyFF_keystate_gff_15_U8 ( .A1(keyFF_keystate_gff_15_n58), .A2(
        keyFF_keystate_gff_15_n57), .ZN(keyFF_keystate_gff_15_n32) );
  NAND2_X1 keyFF_keystate_gff_15_U7 ( .A1(keyFF_keystate_gff_15_n67), .A2(
        keyFF_outputPar[52]), .ZN(keyFF_keystate_gff_15_n57) );
  NOR2_X1 keyFF_keystate_gff_15_U6 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_keystate_gff_15_n56), .ZN(keyFF_keystate_gff_15_n67) );
  MUX2_X1 keyFF_keystate_gff_15_U5 ( .A(keyFF_keystate_gff_15_n36), .B(
        keyFF_keystate_gff_15_n55), .S(keyFF_keystate_gff_15_n65), .Z(
        keyFF_keystate_gff_15_n58) );
  INV_X1 keyFF_keystate_gff_15_U4 ( .A(keyFF_keystate_gff_15_n56), .ZN(
        keyFF_keystate_gff_15_n65) );
  INV_X1 keyFF_keystate_gff_15_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_15_n56) );
  NAND2_X1 keyFF_keystate_gff_15_U2 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[56]), .ZN(keyFF_keystate_gff_15_n55) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_15_n32), .CK(clk), .Q(keyFF_outputPar[56]), .QN(
        keyFF_keystate_gff_15_n36) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_15_n31), .CK(clk), .Q(keyFF_outputPar[57]), .QN(
        keyFF_keystate_gff_15_n35) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_15_n30), .CK(clk), .Q(keyFF_outputPar[58]), .QN(
        keyFF_keystate_gff_15_n34) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_15_n29), .CK(clk), .Q(keyFF_outputPar[59]), .QN(
        keyFF_keystate_gff_15_n33) );
  NAND2_X1 keyFF_keystate_gff_16_U20 ( .A1(keyFF_keystate_gff_16_n69), .A2(
        keyFF_keystate_gff_16_n68), .ZN(keyFF_keystate_gff_16_n29) );
  NAND2_X1 keyFF_keystate_gff_16_U19 ( .A1(keyFF_keystate_gff_16_n67), .A2(
        keyFF_outputPar[59]), .ZN(keyFF_keystate_gff_16_n68) );
  MUX2_X1 keyFF_keystate_gff_16_U18 ( .A(keyFF_keystate_gff_16_n33), .B(
        keyFF_keystate_gff_16_n66), .S(keyFF_keystate_gff_16_n65), .Z(
        keyFF_keystate_gff_16_n69) );
  NAND2_X1 keyFF_keystate_gff_16_U17 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[63]), .ZN(keyFF_keystate_gff_16_n66) );
  NAND2_X1 keyFF_keystate_gff_16_U16 ( .A1(keyFF_keystate_gff_16_n64), .A2(
        keyFF_keystate_gff_16_n63), .ZN(keyFF_keystate_gff_16_n30) );
  NAND2_X1 keyFF_keystate_gff_16_U15 ( .A1(keyFF_keystate_gff_16_n67), .A2(
        keyFF_outputPar[58]), .ZN(keyFF_keystate_gff_16_n63) );
  MUX2_X1 keyFF_keystate_gff_16_U14 ( .A(keyFF_keystate_gff_16_n34), .B(
        keyFF_keystate_gff_16_n62), .S(keyFF_keystate_gff_16_n65), .Z(
        keyFF_keystate_gff_16_n64) );
  NAND2_X1 keyFF_keystate_gff_16_U13 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[62]), .ZN(keyFF_keystate_gff_16_n62) );
  NAND2_X1 keyFF_keystate_gff_16_U12 ( .A1(keyFF_keystate_gff_16_n61), .A2(
        keyFF_keystate_gff_16_n60), .ZN(keyFF_keystate_gff_16_n31) );
  NAND2_X1 keyFF_keystate_gff_16_U11 ( .A1(keyFF_keystate_gff_16_n67), .A2(
        keyFF_outputPar[57]), .ZN(keyFF_keystate_gff_16_n60) );
  MUX2_X1 keyFF_keystate_gff_16_U10 ( .A(keyFF_keystate_gff_16_n35), .B(
        keyFF_keystate_gff_16_n59), .S(keyFF_keystate_gff_16_n65), .Z(
        keyFF_keystate_gff_16_n61) );
  NAND2_X1 keyFF_keystate_gff_16_U9 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[61]), .ZN(keyFF_keystate_gff_16_n59) );
  NAND2_X1 keyFF_keystate_gff_16_U8 ( .A1(keyFF_keystate_gff_16_n58), .A2(
        keyFF_keystate_gff_16_n57), .ZN(keyFF_keystate_gff_16_n32) );
  NAND2_X1 keyFF_keystate_gff_16_U7 ( .A1(keyFF_keystate_gff_16_n67), .A2(
        keyFF_outputPar[56]), .ZN(keyFF_keystate_gff_16_n57) );
  NOR2_X1 keyFF_keystate_gff_16_U6 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_keystate_gff_16_n56), .ZN(keyFF_keystate_gff_16_n67) );
  MUX2_X1 keyFF_keystate_gff_16_U5 ( .A(keyFF_keystate_gff_16_n36), .B(
        keyFF_keystate_gff_16_n55), .S(keyFF_keystate_gff_16_n65), .Z(
        keyFF_keystate_gff_16_n58) );
  INV_X1 keyFF_keystate_gff_16_U4 ( .A(keyFF_keystate_gff_16_n56), .ZN(
        keyFF_keystate_gff_16_n65) );
  INV_X1 keyFF_keystate_gff_16_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_16_n56) );
  NAND2_X1 keyFF_keystate_gff_16_U2 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[60]), .ZN(keyFF_keystate_gff_16_n55) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_16_n32), .CK(clk), .Q(keyFF_outputPar[60]), .QN(
        keyFF_keystate_gff_16_n36) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_16_n31), .CK(clk), .Q(keyFF_outputPar[61]), .QN(
        keyFF_keystate_gff_16_n35) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_16_n30), .CK(clk), .Q(keyFF_outputPar[62]), .QN(
        keyFF_keystate_gff_16_n34) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_16_n29), .CK(clk), .Q(keyFF_outputPar[63]), .QN(
        keyFF_keystate_gff_16_n33) );
  NAND2_X1 keyFF_keystate_gff_17_U20 ( .A1(keyFF_keystate_gff_17_n69), .A2(
        keyFF_keystate_gff_17_n68), .ZN(keyFF_keystate_gff_17_n29) );
  NAND2_X1 keyFF_keystate_gff_17_U19 ( .A1(keyFF_keystate_gff_17_n67), .A2(
        keyFF_outputPar[63]), .ZN(keyFF_keystate_gff_17_n68) );
  MUX2_X1 keyFF_keystate_gff_17_U18 ( .A(keyFF_keystate_gff_17_n33), .B(
        keyFF_keystate_gff_17_n66), .S(keyFF_keystate_gff_17_n65), .Z(
        keyFF_keystate_gff_17_n69) );
  NAND2_X1 keyFF_keystate_gff_17_U17 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[67]), .ZN(keyFF_keystate_gff_17_n66) );
  NAND2_X1 keyFF_keystate_gff_17_U16 ( .A1(keyFF_keystate_gff_17_n64), .A2(
        keyFF_keystate_gff_17_n63), .ZN(keyFF_keystate_gff_17_n30) );
  NAND2_X1 keyFF_keystate_gff_17_U15 ( .A1(keyFF_keystate_gff_17_n67), .A2(
        keyFF_outputPar[62]), .ZN(keyFF_keystate_gff_17_n63) );
  MUX2_X1 keyFF_keystate_gff_17_U14 ( .A(keyFF_keystate_gff_17_n34), .B(
        keyFF_keystate_gff_17_n62), .S(keyFF_keystate_gff_17_n65), .Z(
        keyFF_keystate_gff_17_n64) );
  NAND2_X1 keyFF_keystate_gff_17_U13 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[66]), .ZN(keyFF_keystate_gff_17_n62) );
  NAND2_X1 keyFF_keystate_gff_17_U12 ( .A1(keyFF_keystate_gff_17_n61), .A2(
        keyFF_keystate_gff_17_n60), .ZN(keyFF_keystate_gff_17_n31) );
  NAND2_X1 keyFF_keystate_gff_17_U11 ( .A1(keyFF_keystate_gff_17_n67), .A2(
        keyFF_outputPar[61]), .ZN(keyFF_keystate_gff_17_n60) );
  MUX2_X1 keyFF_keystate_gff_17_U10 ( .A(keyFF_keystate_gff_17_n35), .B(
        keyFF_keystate_gff_17_n59), .S(keyFF_keystate_gff_17_n65), .Z(
        keyFF_keystate_gff_17_n61) );
  NAND2_X1 keyFF_keystate_gff_17_U9 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[65]), .ZN(keyFF_keystate_gff_17_n59) );
  NAND2_X1 keyFF_keystate_gff_17_U8 ( .A1(keyFF_keystate_gff_17_n58), .A2(
        keyFF_keystate_gff_17_n57), .ZN(keyFF_keystate_gff_17_n32) );
  NAND2_X1 keyFF_keystate_gff_17_U7 ( .A1(keyFF_keystate_gff_17_n67), .A2(
        keyFF_outputPar[60]), .ZN(keyFF_keystate_gff_17_n57) );
  NOR2_X1 keyFF_keystate_gff_17_U6 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_keystate_gff_17_n56), .ZN(keyFF_keystate_gff_17_n67) );
  MUX2_X1 keyFF_keystate_gff_17_U5 ( .A(keyFF_keystate_gff_17_n36), .B(
        keyFF_keystate_gff_17_n55), .S(keyFF_keystate_gff_17_n65), .Z(
        keyFF_keystate_gff_17_n58) );
  INV_X1 keyFF_keystate_gff_17_U4 ( .A(keyFF_keystate_gff_17_n56), .ZN(
        keyFF_keystate_gff_17_n65) );
  INV_X1 keyFF_keystate_gff_17_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_17_n56) );
  NAND2_X1 keyFF_keystate_gff_17_U2 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[64]), .ZN(keyFF_keystate_gff_17_n55) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_17_n32), .CK(clk), .Q(keyFF_outputPar[64]), .QN(
        keyFF_keystate_gff_17_n36) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_17_n31), .CK(clk), .Q(keyFF_outputPar[65]), .QN(
        keyFF_keystate_gff_17_n35) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_17_n30), .CK(clk), .Q(keyFF_outputPar[66]), .QN(
        keyFF_keystate_gff_17_n34) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_17_n29), .CK(clk), .Q(keyFF_outputPar[67]), .QN(
        keyFF_keystate_gff_17_n33) );
  NAND2_X1 keyFF_keystate_gff_18_U20 ( .A1(keyFF_keystate_gff_18_n69), .A2(
        keyFF_keystate_gff_18_n68), .ZN(keyFF_keystate_gff_18_n29) );
  NAND2_X1 keyFF_keystate_gff_18_U19 ( .A1(keyFF_keystate_gff_18_n67), .A2(
        keyFF_outputPar[67]), .ZN(keyFF_keystate_gff_18_n68) );
  MUX2_X1 keyFF_keystate_gff_18_U18 ( .A(keyFF_keystate_gff_18_n33), .B(
        keyFF_keystate_gff_18_n66), .S(keyFF_keystate_gff_18_n65), .Z(
        keyFF_keystate_gff_18_n69) );
  NAND2_X1 keyFF_keystate_gff_18_U17 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[71]), .ZN(keyFF_keystate_gff_18_n66) );
  NAND2_X1 keyFF_keystate_gff_18_U16 ( .A1(keyFF_keystate_gff_18_n64), .A2(
        keyFF_keystate_gff_18_n63), .ZN(keyFF_keystate_gff_18_n30) );
  NAND2_X1 keyFF_keystate_gff_18_U15 ( .A1(keyFF_keystate_gff_18_n67), .A2(
        keyFF_outputPar[66]), .ZN(keyFF_keystate_gff_18_n63) );
  MUX2_X1 keyFF_keystate_gff_18_U14 ( .A(keyFF_keystate_gff_18_n34), .B(
        keyFF_keystate_gff_18_n62), .S(keyFF_keystate_gff_18_n65), .Z(
        keyFF_keystate_gff_18_n64) );
  NAND2_X1 keyFF_keystate_gff_18_U13 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[70]), .ZN(keyFF_keystate_gff_18_n62) );
  NAND2_X1 keyFF_keystate_gff_18_U12 ( .A1(keyFF_keystate_gff_18_n61), .A2(
        keyFF_keystate_gff_18_n60), .ZN(keyFF_keystate_gff_18_n31) );
  NAND2_X1 keyFF_keystate_gff_18_U11 ( .A1(keyFF_keystate_gff_18_n67), .A2(
        keyFF_outputPar[65]), .ZN(keyFF_keystate_gff_18_n60) );
  MUX2_X1 keyFF_keystate_gff_18_U10 ( .A(keyFF_keystate_gff_18_n35), .B(
        keyFF_keystate_gff_18_n59), .S(keyFF_keystate_gff_18_n65), .Z(
        keyFF_keystate_gff_18_n61) );
  NAND2_X1 keyFF_keystate_gff_18_U9 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[69]), .ZN(keyFF_keystate_gff_18_n59) );
  NAND2_X1 keyFF_keystate_gff_18_U8 ( .A1(keyFF_keystate_gff_18_n58), .A2(
        keyFF_keystate_gff_18_n57), .ZN(keyFF_keystate_gff_18_n32) );
  NAND2_X1 keyFF_keystate_gff_18_U7 ( .A1(keyFF_keystate_gff_18_n67), .A2(
        keyFF_outputPar[64]), .ZN(keyFF_keystate_gff_18_n57) );
  NOR2_X1 keyFF_keystate_gff_18_U6 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_keystate_gff_18_n56), .ZN(keyFF_keystate_gff_18_n67) );
  MUX2_X1 keyFF_keystate_gff_18_U5 ( .A(keyFF_keystate_gff_18_n36), .B(
        keyFF_keystate_gff_18_n55), .S(keyFF_keystate_gff_18_n65), .Z(
        keyFF_keystate_gff_18_n58) );
  INV_X1 keyFF_keystate_gff_18_U4 ( .A(keyFF_keystate_gff_18_n56), .ZN(
        keyFF_keystate_gff_18_n65) );
  INV_X1 keyFF_keystate_gff_18_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_18_n56) );
  NAND2_X1 keyFF_keystate_gff_18_U2 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[68]), .ZN(keyFF_keystate_gff_18_n55) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_18_n32), .CK(clk), .Q(keyFF_outputPar[68]), .QN(
        keyFF_keystate_gff_18_n36) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_18_n31), .CK(clk), .Q(keyFF_outputPar[69]), .QN(
        keyFF_keystate_gff_18_n35) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_18_n30), .CK(clk), .Q(keyFF_outputPar[70]), .QN(
        keyFF_keystate_gff_18_n34) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_18_n29), .CK(clk), .Q(keyFF_outputPar[71]), .QN(
        keyFF_keystate_gff_18_n33) );
  NAND2_X1 keyFF_keystate_gff_19_U20 ( .A1(keyFF_keystate_gff_19_n68), .A2(
        keyFF_keystate_gff_19_n67), .ZN(keyFF_keystate_gff_19_n28) );
  NAND2_X1 keyFF_keystate_gff_19_U19 ( .A1(keyFF_keystate_gff_19_n66), .A2(
        keyFF_outputPar[71]), .ZN(keyFF_keystate_gff_19_n67) );
  MUX2_X1 keyFF_keystate_gff_19_U18 ( .A(keyFF_keystate_gff_19_n32), .B(
        keyFF_keystate_gff_19_n65), .S(keyFF_keystate_gff_19_n64), .Z(
        keyFF_keystate_gff_19_n68) );
  NAND2_X1 keyFF_keystate_gff_19_U17 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[75]), .ZN(keyFF_keystate_gff_19_n65) );
  NAND2_X1 keyFF_keystate_gff_19_U16 ( .A1(keyFF_keystate_gff_19_n63), .A2(
        keyFF_keystate_gff_19_n62), .ZN(keyFF_keystate_gff_19_n29) );
  NAND2_X1 keyFF_keystate_gff_19_U15 ( .A1(keyFF_keystate_gff_19_n66), .A2(
        keyFF_outputPar[70]), .ZN(keyFF_keystate_gff_19_n62) );
  MUX2_X1 keyFF_keystate_gff_19_U14 ( .A(keyFF_keystate_gff_19_n33), .B(
        keyFF_keystate_gff_19_n61), .S(keyFF_keystate_gff_19_n64), .Z(
        keyFF_keystate_gff_19_n63) );
  NAND2_X1 keyFF_keystate_gff_19_U13 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[74]), .ZN(keyFF_keystate_gff_19_n61) );
  NAND2_X1 keyFF_keystate_gff_19_U12 ( .A1(keyFF_keystate_gff_19_n60), .A2(
        keyFF_keystate_gff_19_n59), .ZN(keyFF_keystate_gff_19_n30) );
  NAND2_X1 keyFF_keystate_gff_19_U11 ( .A1(keyFF_keystate_gff_19_n66), .A2(
        keyFF_outputPar[69]), .ZN(keyFF_keystate_gff_19_n59) );
  MUX2_X1 keyFF_keystate_gff_19_U10 ( .A(keyFF_keystate_gff_19_n34), .B(
        keyFF_keystate_gff_19_n58), .S(keyFF_keystate_gff_19_n64), .Z(
        keyFF_keystate_gff_19_n60) );
  NAND2_X1 keyFF_keystate_gff_19_U9 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[73]), .ZN(keyFF_keystate_gff_19_n58) );
  NAND2_X1 keyFF_keystate_gff_19_U8 ( .A1(keyFF_keystate_gff_19_n57), .A2(
        keyFF_keystate_gff_19_n56), .ZN(keyFF_keystate_gff_19_n31) );
  NAND2_X1 keyFF_keystate_gff_19_U7 ( .A1(keyFF_keystate_gff_19_n66), .A2(
        keyFF_outputPar[68]), .ZN(keyFF_keystate_gff_19_n56) );
  NOR2_X1 keyFF_keystate_gff_19_U6 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_keystate_gff_19_n55), .ZN(keyFF_keystate_gff_19_n66) );
  MUX2_X1 keyFF_keystate_gff_19_U5 ( .A(keyFF_keystate_gff_19_n35), .B(
        keyFF_keystate_gff_19_n54), .S(keyFF_keystate_gff_19_n64), .Z(
        keyFF_keystate_gff_19_n57) );
  INV_X1 keyFF_keystate_gff_19_U4 ( .A(keyFF_keystate_gff_19_n55), .ZN(
        keyFF_keystate_gff_19_n64) );
  INV_X1 keyFF_keystate_gff_19_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_19_n55) );
  NAND2_X1 keyFF_keystate_gff_19_U2 ( .A1(keyFF_keystate_n7), .A2(
        keyFF_inputPar[72]), .ZN(keyFF_keystate_gff_19_n54) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_19_n31), .CK(clk), .Q(keyFF_outputPar[72]), .QN(
        keyFF_keystate_gff_19_n35) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_19_n30), .CK(clk), .Q(keyFF_outputPar[73]), .QN(
        keyFF_keystate_gff_19_n34) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_19_n29), .CK(clk), .Q(keyFF_outputPar[74]), .QN(
        keyFF_keystate_gff_19_n33) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_19_n28), .CK(clk), .Q(keyFF_outputPar[75]), .QN(
        keyFF_keystate_gff_19_n32) );
  NAND2_X1 keyFF_keystate_gff_20_U20 ( .A1(keyFF_keystate_gff_20_n68), .A2(
        keyFF_keystate_gff_20_n67), .ZN(keyFF_keystate_gff_20_n28) );
  NAND2_X1 keyFF_keystate_gff_20_U19 ( .A1(keyFF_keystate_gff_20_n66), .A2(
        keyFF_outputPar[75]), .ZN(keyFF_keystate_gff_20_n67) );
  MUX2_X1 keyFF_keystate_gff_20_U18 ( .A(keyFF_keystate_gff_20_n32), .B(
        keyFF_keystate_gff_20_n65), .S(keyFF_keystate_gff_20_n64), .Z(
        keyFF_keystate_gff_20_n68) );
  NAND2_X1 keyFF_keystate_gff_20_U17 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[79]), .ZN(keyFF_keystate_gff_20_n65) );
  NAND2_X1 keyFF_keystate_gff_20_U16 ( .A1(keyFF_keystate_gff_20_n63), .A2(
        keyFF_keystate_gff_20_n62), .ZN(keyFF_keystate_gff_20_n29) );
  NAND2_X1 keyFF_keystate_gff_20_U15 ( .A1(keyFF_keystate_gff_20_n66), .A2(
        keyFF_outputPar[74]), .ZN(keyFF_keystate_gff_20_n62) );
  MUX2_X1 keyFF_keystate_gff_20_U14 ( .A(keyFF_keystate_gff_20_n33), .B(
        keyFF_keystate_gff_20_n61), .S(keyFF_keystate_gff_20_n64), .Z(
        keyFF_keystate_gff_20_n63) );
  NAND2_X1 keyFF_keystate_gff_20_U13 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[78]), .ZN(keyFF_keystate_gff_20_n61) );
  NAND2_X1 keyFF_keystate_gff_20_U12 ( .A1(keyFF_keystate_gff_20_n60), .A2(
        keyFF_keystate_gff_20_n59), .ZN(keyFF_keystate_gff_20_n30) );
  NAND2_X1 keyFF_keystate_gff_20_U11 ( .A1(keyFF_keystate_gff_20_n66), .A2(
        keyFF_outputPar[73]), .ZN(keyFF_keystate_gff_20_n59) );
  MUX2_X1 keyFF_keystate_gff_20_U10 ( .A(keyFF_keystate_gff_20_n34), .B(
        keyFF_keystate_gff_20_n58), .S(keyFF_keystate_gff_20_n64), .Z(
        keyFF_keystate_gff_20_n60) );
  NAND2_X1 keyFF_keystate_gff_20_U9 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[77]), .ZN(keyFF_keystate_gff_20_n58) );
  NAND2_X1 keyFF_keystate_gff_20_U8 ( .A1(keyFF_keystate_gff_20_n57), .A2(
        keyFF_keystate_gff_20_n56), .ZN(keyFF_keystate_gff_20_n31) );
  NAND2_X1 keyFF_keystate_gff_20_U7 ( .A1(keyFF_keystate_gff_20_n66), .A2(
        keyFF_outputPar[72]), .ZN(keyFF_keystate_gff_20_n56) );
  NOR2_X1 keyFF_keystate_gff_20_U6 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_keystate_gff_20_n55), .ZN(keyFF_keystate_gff_20_n66) );
  MUX2_X1 keyFF_keystate_gff_20_U5 ( .A(keyFF_keystate_gff_20_n35), .B(
        keyFF_keystate_gff_20_n54), .S(keyFF_keystate_gff_20_n64), .Z(
        keyFF_keystate_gff_20_n57) );
  INV_X1 keyFF_keystate_gff_20_U4 ( .A(keyFF_keystate_gff_20_n55), .ZN(
        keyFF_keystate_gff_20_n64) );
  INV_X1 keyFF_keystate_gff_20_U3 ( .A(ctrlData[1]), .ZN(
        keyFF_keystate_gff_20_n55) );
  NAND2_X1 keyFF_keystate_gff_20_U2 ( .A1(keyFF_keystate_n6), .A2(
        keyFF_inputPar[76]), .ZN(keyFF_keystate_gff_20_n54) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_0_ ( .D(
        keyFF_keystate_gff_20_n31), .CK(clk), .Q(roundkey[0]), .QN(
        keyFF_keystate_gff_20_n35) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_1_ ( .D(
        keyFF_keystate_gff_20_n30), .CK(clk), .Q(roundkey[1]), .QN(
        keyFF_keystate_gff_20_n34) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_2_ ( .D(
        keyFF_keystate_gff_20_n29), .CK(clk), .Q(roundkey[2]), .QN(
        keyFF_keystate_gff_20_n33) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_3_ ( .D(
        keyFF_keystate_gff_20_n28), .CK(clk), .Q(roundkey[3]), .QN(
        keyFF_keystate_gff_20_n32) );
  NAND2_X1 sboxInst_U22 ( .A1(sboxInst_n25), .A2(sboxInst_n24), .ZN(sboxOut[2]) );
  NAND2_X1 sboxInst_U21 ( .A1(sboxInst_n23), .A2(sboxInst_n22), .ZN(
        sboxInst_n24) );
  NAND2_X1 sboxInst_U20 ( .A1(sboxInst_n21), .A2(sboxInst_n20), .ZN(
        sboxInst_n25) );
  NOR2_X1 sboxInst_U19 ( .A1(keyRegKS[2]), .A2(sboxInst_n19), .ZN(sboxInst_n21) );
  NOR2_X1 sboxInst_U18 ( .A1(sboxInst_n19), .A2(sboxInst_n18), .ZN(sboxOut[3])
         );
  MUX2_X1 sboxInst_U17 ( .A(keyRegKS[2]), .B(sboxInst_n17), .S(sboxInst_n16), 
        .Z(sboxInst_n18) );
  AND2_X1 sboxInst_U16 ( .A1(sboxInst_n20), .A2(sboxInst_n15), .ZN(
        sboxInst_n17) );
  NOR2_X1 sboxInst_U15 ( .A1(sboxInst_n16), .A2(sboxInst_n15), .ZN(
        sboxInst_n19) );
  OR2_X1 sboxInst_U14 ( .A1(keyRegKS[1]), .A2(roundkey[3]), .ZN(sboxInst_n15)
         );
  MUX2_X1 sboxInst_U13 ( .A(sboxInst_n23), .B(sboxInst_n14), .S(sboxInst_n22), 
        .Z(sboxOut[1]) );
  NOR2_X1 sboxInst_U12 ( .A1(sboxInst_n13), .A2(sboxInst_n12), .ZN(
        sboxInst_n22) );
  MUX2_X1 sboxInst_U11 ( .A(sboxInst_n20), .B(keyRegKS[1]), .S(sboxInst_n16), 
        .Z(sboxInst_n23) );
  NAND2_X1 sboxInst_U10 ( .A1(keyRegKS[1]), .A2(sboxInst_n11), .ZN(
        sboxInst_n20) );
  NAND2_X1 sboxInst_U9 ( .A1(sboxInst_n10), .A2(sboxInst_n12), .ZN(
        sboxInst_n11) );
  XOR2_X1 sboxInst_U8 ( .A(sboxInst_n9), .B(sboxInst_n8), .Z(sboxOut[0]) );
  NOR2_X1 sboxInst_U7 ( .A1(sboxInst_n12), .A2(keyRegKS[1]), .ZN(sboxInst_n8)
         );
  INV_X1 sboxInst_U6 ( .A(keyRegKS[2]), .ZN(sboxInst_n12) );
  NOR2_X1 sboxInst_U5 ( .A1(sboxInst_n13), .A2(sboxInst_n14), .ZN(sboxInst_n9)
         );
  NOR2_X1 sboxInst_U4 ( .A1(sboxInst_n16), .A2(sboxInst_n10), .ZN(sboxInst_n14) );
  INV_X1 sboxInst_U3 ( .A(roundkey[3]), .ZN(sboxInst_n10) );
  INV_X1 sboxInst_U2 ( .A(keyRegKS[3]), .ZN(sboxInst_n16) );
  NOR2_X1 sboxInst_U1 ( .A1(keyRegKS[3]), .A2(roundkey[3]), .ZN(sboxInst_n13)
         );
  XOR2_X1 sboxTI_f1_U17 ( .A(sboxTI_g2Reg[0]), .B(stateFF_permOut[16]), .Z(
        stateFF_permOut[48]) );
  XNOR2_X1 sboxTI_f1_U16 ( .A(sboxTI_f1_n13), .B(sboxTI_f1_n12), .ZN(
        stateFF_permOut[16]) );
  XNOR2_X1 sboxTI_f1_U15 ( .A(sboxTI_f1_n11), .B(sboxTI_f1_n10), .ZN(
        sboxTI_f1_n12) );
  NAND2_X1 sboxTI_f1_U14 ( .A1(sboxTI_g3Reg[0]), .A2(sboxTI_g2Reg[3]), .ZN(
        sboxTI_f1_n10) );
  XOR2_X1 sboxTI_f1_U13 ( .A(sboxTI_g2Reg[1]), .B(sboxTI_g2Reg[2]), .Z(
        sboxTI_f1_n11) );
  NAND2_X1 sboxTI_f1_U12 ( .A1(sboxTI_f1_n9), .A2(sboxTI_g2Reg[0]), .ZN(
        sboxTI_f1_n13) );
  XOR2_X1 sboxTI_f1_U11 ( .A(sboxTI_g3Reg[3]), .B(sboxTI_g2Reg[3]), .Z(
        sboxTI_f1_n9) );
  XNOR2_X1 sboxTI_f1_U10 ( .A(sboxTI_g2Reg[1]), .B(sboxTI_f1_n8), .ZN(
        stateFF_permOut[0]) );
  XNOR2_X1 sboxTI_f1_U9 ( .A(sboxTI_f1_n7), .B(sboxTI_f1_n6), .ZN(sboxTI_f1_n8) );
  NAND2_X1 sboxTI_f1_U8 ( .A1(sboxTI_f1_n5), .A2(sboxTI_g2Reg[0]), .ZN(
        sboxTI_f1_n6) );
  XOR2_X1 sboxTI_f1_U7 ( .A(sboxTI_g2Reg[2]), .B(sboxTI_g3Reg[2]), .Z(
        sboxTI_f1_n5) );
  NAND2_X1 sboxTI_f1_U6 ( .A1(sboxTI_g2Reg[2]), .A2(sboxTI_g3Reg[0]), .ZN(
        sboxTI_f1_n7) );
  XNOR2_X1 sboxTI_f1_U5 ( .A(sboxTI_g2Reg[3]), .B(sboxTI_f1_n4), .ZN(
        stateFF_permOut[32]) );
  XNOR2_X1 sboxTI_f1_U4 ( .A(sboxTI_f1_n3), .B(sboxTI_f1_n2), .ZN(sboxTI_f1_n4) );
  NAND2_X1 sboxTI_f1_U3 ( .A1(sboxTI_g3Reg[1]), .A2(sboxTI_g2Reg[0]), .ZN(
        sboxTI_f1_n2) );
  NAND2_X1 sboxTI_f1_U2 ( .A1(sboxTI_g2Reg[1]), .A2(sboxTI_f1_n1), .ZN(
        sboxTI_f1_n3) );
  XOR2_X1 sboxTI_f1_U1 ( .A(sboxTI_g2Reg[0]), .B(sboxTI_g3Reg[0]), .Z(
        sboxTI_f1_n1) );
  XOR2_X1 sboxTI_f2_U15 ( .A(sboxTI_g3Reg[0]), .B(md1FF_permOut[16]), .Z(
        md1FF_permOut[48]) );
  XNOR2_X1 sboxTI_f2_U14 ( .A(sboxTI_f2_n11), .B(sboxTI_f2_n10), .ZN(
        md1FF_permOut[16]) );
  XNOR2_X1 sboxTI_f2_U13 ( .A(sboxTI_f2_n9), .B(sboxTI_f2_n8), .ZN(
        sboxTI_f2_n10) );
  NAND2_X1 sboxTI_f2_U12 ( .A1(sboxTI_g3Reg[3]), .A2(sboxTI_f2_n7), .ZN(
        sboxTI_f2_n8) );
  XOR2_X1 sboxTI_f2_U11 ( .A(sboxTI_g3Reg[2]), .B(sboxTI_g3Reg[1]), .Z(
        sboxTI_f2_n9) );
  NAND2_X1 sboxTI_f2_U10 ( .A1(sboxTI_g1Reg[3]), .A2(sboxTI_g3Reg[0]), .ZN(
        sboxTI_f2_n11) );
  XNOR2_X1 sboxTI_f2_U9 ( .A(sboxTI_g3Reg[1]), .B(sboxTI_f2_n6), .ZN(
        md1FF_permOut[0]) );
  XNOR2_X1 sboxTI_f2_U8 ( .A(sboxTI_f2_n5), .B(sboxTI_f2_n4), .ZN(sboxTI_f2_n6) );
  NAND2_X1 sboxTI_f2_U7 ( .A1(sboxTI_g1Reg[2]), .A2(sboxTI_g3Reg[0]), .ZN(
        sboxTI_f2_n4) );
  NAND2_X1 sboxTI_f2_U6 ( .A1(sboxTI_f2_n7), .A2(sboxTI_g3Reg[2]), .ZN(
        sboxTI_f2_n5) );
  XNOR2_X1 sboxTI_f2_U5 ( .A(sboxTI_g3Reg[3]), .B(sboxTI_f2_n3), .ZN(
        md1FF_permOut[32]) );
  XNOR2_X1 sboxTI_f2_U4 ( .A(sboxTI_f2_n2), .B(sboxTI_f2_n1), .ZN(sboxTI_f2_n3) );
  NAND2_X1 sboxTI_f2_U3 ( .A1(sboxTI_g1Reg[1]), .A2(sboxTI_g3Reg[0]), .ZN(
        sboxTI_f2_n1) );
  NAND2_X1 sboxTI_f2_U2 ( .A1(sboxTI_f2_n7), .A2(sboxTI_g3Reg[1]), .ZN(
        sboxTI_f2_n2) );
  XOR2_X1 sboxTI_f2_U1 ( .A(sboxTI_g3Reg[0]), .B(sboxTI_g1Reg[0]), .Z(
        sboxTI_f2_n7) );
  XOR2_X1 sboxTI_f3_U17 ( .A(sboxTI_g1Reg[0]), .B(md2FF_permOut[16]), .Z(
        md2FF_permOut[48]) );
  XNOR2_X1 sboxTI_f3_U16 ( .A(sboxTI_f3_n13), .B(sboxTI_f3_n12), .ZN(
        md2FF_permOut[16]) );
  XNOR2_X1 sboxTI_f3_U15 ( .A(sboxTI_f3_n11), .B(sboxTI_f3_n10), .ZN(
        sboxTI_f3_n12) );
  NAND2_X1 sboxTI_f3_U14 ( .A1(sboxTI_g2Reg[0]), .A2(sboxTI_g1Reg[3]), .ZN(
        sboxTI_f3_n10) );
  XOR2_X1 sboxTI_f3_U13 ( .A(sboxTI_g1Reg[1]), .B(sboxTI_g1Reg[2]), .Z(
        sboxTI_f3_n11) );
  NAND2_X1 sboxTI_f3_U12 ( .A1(sboxTI_f3_n9), .A2(sboxTI_g1Reg[0]), .ZN(
        sboxTI_f3_n13) );
  XOR2_X1 sboxTI_f3_U11 ( .A(sboxTI_g2Reg[3]), .B(sboxTI_g1Reg[3]), .Z(
        sboxTI_f3_n9) );
  XNOR2_X1 sboxTI_f3_U10 ( .A(sboxTI_g1Reg[1]), .B(sboxTI_f3_n8), .ZN(
        md2FF_permOut[0]) );
  XNOR2_X1 sboxTI_f3_U9 ( .A(sboxTI_f3_n7), .B(sboxTI_f3_n6), .ZN(sboxTI_f3_n8) );
  NAND2_X1 sboxTI_f3_U8 ( .A1(sboxTI_f3_n5), .A2(sboxTI_g1Reg[0]), .ZN(
        sboxTI_f3_n6) );
  XOR2_X1 sboxTI_f3_U7 ( .A(sboxTI_g1Reg[2]), .B(sboxTI_g2Reg[2]), .Z(
        sboxTI_f3_n5) );
  NAND2_X1 sboxTI_f3_U6 ( .A1(sboxTI_g1Reg[2]), .A2(sboxTI_g2Reg[0]), .ZN(
        sboxTI_f3_n7) );
  XNOR2_X1 sboxTI_f3_U5 ( .A(sboxTI_g1Reg[3]), .B(sboxTI_f3_n4), .ZN(
        md2FF_permOut[32]) );
  XNOR2_X1 sboxTI_f3_U4 ( .A(sboxTI_f3_n3), .B(sboxTI_f3_n2), .ZN(sboxTI_f3_n4) );
  NAND2_X1 sboxTI_f3_U3 ( .A1(sboxTI_g2Reg[1]), .A2(sboxTI_g1Reg[0]), .ZN(
        sboxTI_f3_n2) );
  NAND2_X1 sboxTI_f3_U2 ( .A1(sboxTI_g1Reg[1]), .A2(sboxTI_f3_n1), .ZN(
        sboxTI_f3_n3) );
  XOR2_X1 sboxTI_f3_U1 ( .A(sboxTI_g1Reg[0]), .B(sboxTI_g2Reg[0]), .Z(
        sboxTI_f3_n1) );
  XNOR2_X1 sboxTI_g1_U26 ( .A(md1Reg[0]), .B(sboxTI_g1Out[2]), .ZN(
        sboxTI_g1Out[3]) );
  XOR2_X1 sboxTI_g1_U25 ( .A(sboxTI_g1_n22), .B(sboxTI_g1_n21), .Z(
        sboxTI_g1Out[0]) );
  NAND2_X1 sboxTI_g1_U24 ( .A1(sboxTI_g1_n20), .A2(sboxTI_g1_n19), .ZN(
        sboxTI_g1_n21) );
  OR2_X1 sboxTI_g1_U23 ( .A1(md1Reg[2]), .A2(md1Reg[1]), .ZN(sboxTI_g1_n19) );
  NAND2_X1 sboxTI_g1_U22 ( .A1(sboxTI_g1_n18), .A2(sboxTI_g1_n17), .ZN(
        sboxTI_g1_n20) );
  NAND2_X1 sboxTI_g1_U21 ( .A1(md1Reg[2]), .A2(md1Reg[1]), .ZN(sboxTI_g1_n17)
         );
  XNOR2_X1 sboxTI_g1_U20 ( .A(md1Reg[3]), .B(md2Reg[3]), .ZN(sboxTI_g1_n18) );
  XNOR2_X1 sboxTI_g1_U19 ( .A(sboxTI_g1_n16), .B(sboxTI_g1_n15), .ZN(
        sboxTI_g1_n22) );
  NAND2_X1 sboxTI_g1_U18 ( .A1(sboxTI_g1_n14), .A2(md1Reg[3]), .ZN(
        sboxTI_g1_n15) );
  XOR2_X1 sboxTI_g1_U17 ( .A(md2Reg[1]), .B(md2Reg[2]), .Z(sboxTI_g1_n14) );
  XOR2_X1 sboxTI_g1_U16 ( .A(md1Reg[0]), .B(sboxTI_g1_n13), .Z(sboxTI_g1_n16)
         );
  XOR2_X1 sboxTI_g1_U15 ( .A(sboxTI_g1_n12), .B(sboxTI_g1_n11), .Z(
        sboxTI_g1_n13) );
  NAND2_X1 sboxTI_g1_U14 ( .A1(md2Reg[1]), .A2(md1Reg[2]), .ZN(sboxTI_g1_n11)
         );
  NAND2_X1 sboxTI_g1_U13 ( .A1(md2Reg[2]), .A2(md1Reg[1]), .ZN(sboxTI_g1_n12)
         );
  XNOR2_X1 sboxTI_g1_U12 ( .A(sboxTI_g1_n10), .B(sboxTI_g1_n9), .ZN(
        sboxTI_g1Out[1]) );
  XNOR2_X1 sboxTI_g1_U11 ( .A(sboxTI_g1_n8), .B(sboxTI_g1_n7), .ZN(
        sboxTI_g1_n9) );
  XOR2_X1 sboxTI_g1_U10 ( .A(sboxTI_g1_n6), .B(sboxTI_g1_n5), .Z(sboxTI_g1_n7)
         );
  NAND2_X1 sboxTI_g1_U9 ( .A1(md1Reg[0]), .A2(sboxTI_g1_n4), .ZN(sboxTI_g1_n5)
         );
  XNOR2_X1 sboxTI_g1_U8 ( .A(sboxTI_g1_n3), .B(md2Reg[2]), .ZN(sboxTI_g1_n4)
         );
  XOR2_X1 sboxTI_g1_U7 ( .A(md2Reg[1]), .B(sboxTI_g1Out[2]), .Z(sboxTI_g1_n3)
         );
  NAND2_X1 sboxTI_g1_U6 ( .A1(md1Reg[2]), .A2(md2Reg[0]), .ZN(sboxTI_g1_n6) );
  NAND2_X1 sboxTI_g1_U5 ( .A1(sboxTI_g1_n2), .A2(md1Reg[1]), .ZN(sboxTI_g1_n8)
         );
  XNOR2_X1 sboxTI_g1_U4 ( .A(md1Reg[2]), .B(md2Reg[0]), .ZN(sboxTI_g1_n2) );
  XNOR2_X1 sboxTI_g1_U3 ( .A(md2Reg[3]), .B(sboxTI_g1_n1), .ZN(sboxTI_g1_n10)
         );
  NAND2_X1 sboxTI_g1_U2 ( .A1(md2Reg[1]), .A2(md2Reg[2]), .ZN(sboxTI_g1_n1) );
  XNOR2_X1 sboxTI_g1_U1 ( .A(md1Reg[2]), .B(md1Reg[1]), .ZN(sboxTI_g1Out[2])
         );
  XOR2_X1 sboxTI_g2_U27 ( .A(md2Reg[0]), .B(sboxTI_g2Out[2]), .Z(
        sboxTI_g2Out[3]) );
  XNOR2_X1 sboxTI_g2_U26 ( .A(sboxTI_g2_n23), .B(sboxTI_g2_n22), .ZN(
        sboxTI_g2Out[0]) );
  MUX2_X1 sboxTI_g2_U25 ( .A(sboxTI_g2_n21), .B(sboxTI_g2_n20), .S(md2Reg[1]), 
        .Z(sboxTI_g2_n22) );
  XNOR2_X1 sboxTI_g2_U24 ( .A(sboxTI_g2_n19), .B(sboxTI_g2_n18), .ZN(
        sboxTI_g2_n20) );
  NOR2_X1 sboxTI_g2_U23 ( .A1(sboxIn1[2]), .A2(md2Reg[3]), .ZN(sboxTI_g2_n18)
         );
  NAND2_X1 sboxTI_g2_U22 ( .A1(sboxIn1[2]), .A2(md2Reg[3]), .ZN(sboxTI_g2_n21)
         );
  XNOR2_X1 sboxTI_g2_U21 ( .A(md2Reg[0]), .B(sboxTI_g2_n17), .ZN(sboxTI_g2_n23) );
  MUX2_X1 sboxTI_g2_U20 ( .A(sboxTI_g2_n16), .B(sboxTI_g2_n15), .S(
        sboxTI_g2_n14), .Z(sboxTI_g2_n17) );
  MUX2_X1 sboxTI_g2_U19 ( .A(sboxTI_g2_n13), .B(sboxTI_g2_n12), .S(md2Reg[2]), 
        .Z(sboxTI_g2_n14) );
  NOR2_X1 sboxTI_g2_U18 ( .A1(sboxTI_g2_n11), .A2(sboxTI_g2_n10), .ZN(
        sboxTI_g2_n12) );
  NAND2_X1 sboxTI_g2_U17 ( .A1(sboxIn1[1]), .A2(md2Reg[3]), .ZN(sboxTI_g2_n13)
         );
  NAND2_X1 sboxTI_g2_U16 ( .A1(sboxTI_g2_n15), .A2(sboxTI_g2_n9), .ZN(
        sboxTI_g2_n16) );
  NAND2_X1 sboxTI_g2_U15 ( .A1(sboxTI_g2_n11), .A2(sboxTI_g2_n10), .ZN(
        sboxTI_g2_n9) );
  INV_X1 sboxTI_g2_U14 ( .A(sboxIn1[3]), .ZN(sboxTI_g2_n10) );
  NOR2_X1 sboxTI_g2_U13 ( .A1(md2Reg[3]), .A2(sboxIn1[1]), .ZN(sboxTI_g2_n11)
         );
  NAND2_X1 sboxTI_g2_U12 ( .A1(md2Reg[1]), .A2(sboxIn1[3]), .ZN(sboxTI_g2_n15)
         );
  XNOR2_X1 sboxTI_g2_U11 ( .A(sboxTI_g2_n8), .B(sboxTI_g2_n7), .ZN(
        sboxTI_g2Out[1]) );
  NAND2_X1 sboxTI_g2_U10 ( .A1(md2Reg[0]), .A2(sboxTI_g2_n6), .ZN(sboxTI_g2_n7) );
  XOR2_X1 sboxTI_g2_U9 ( .A(sboxIn1[1]), .B(sboxIn1[2]), .Z(sboxTI_g2_n6) );
  XNOR2_X1 sboxTI_g2_U8 ( .A(sboxTI_g2_n5), .B(sboxTI_g2_n4), .ZN(sboxTI_g2_n8) );
  XNOR2_X1 sboxTI_g2_U7 ( .A(sboxTI_g2_n3), .B(sboxTI_g2_n2), .ZN(sboxTI_g2_n4) );
  NAND2_X1 sboxTI_g2_U6 ( .A1(sboxTI_g2_n1), .A2(sboxTI_g2Out[2]), .ZN(
        sboxTI_g2_n2) );
  XOR2_X1 sboxTI_g2_U5 ( .A(md2Reg[0]), .B(sboxIn1[0]), .Z(sboxTI_g2_n1) );
  XOR2_X1 sboxTI_g2_U4 ( .A(sboxIn1[3]), .B(sboxTI_g2_C), .Z(sboxTI_g2_n3) );
  NAND2_X1 sboxTI_g2_U3 ( .A1(md2Reg[1]), .A2(sboxTI_g2_n19), .ZN(sboxTI_g2_n5) );
  XNOR2_X1 sboxTI_g2_U2 ( .A(md2Reg[1]), .B(sboxTI_g2_n19), .ZN(
        sboxTI_g2Out[2]) );
  INV_X1 sboxTI_g2_U1 ( .A(md2Reg[2]), .ZN(sboxTI_g2_n19) );
  AND2_X1 sboxTI_g2_CtermInst_U1 ( .A1(sboxIn1[1]), .A2(sboxIn1[2]), .ZN(
        sboxTI_g2_C) );
  XOR2_X1 sboxTI_g3_U26 ( .A(sboxIn1[0]), .B(sboxTI_g3Out[2]), .Z(
        sboxTI_g3Out[3]) );
  XNOR2_X1 sboxTI_g3_U25 ( .A(sboxTI_g3_n41), .B(sboxTI_g3_n40), .ZN(
        sboxTI_g3Out[0]) );
  XNOR2_X1 sboxTI_g3_U24 ( .A(sboxTI_g3_n39), .B(sboxTI_g3_n38), .ZN(
        sboxTI_g3_n40) );
  NAND2_X1 sboxTI_g3_U23 ( .A1(sboxTI_g3_n37), .A2(sboxIn1[3]), .ZN(
        sboxTI_g3_n38) );
  NOR2_X1 sboxTI_g3_U22 ( .A1(sboxTI_g3_n36), .A2(sboxTI_g3_n35), .ZN(
        sboxTI_g3_n39) );
  NOR2_X1 sboxTI_g3_U21 ( .A1(sboxIn1[1]), .A2(sboxTI_g3_n34), .ZN(
        sboxTI_g3_n35) );
  AND2_X1 sboxTI_g3_U20 ( .A1(sboxIn1[2]), .A2(md1Reg[3]), .ZN(sboxTI_g3_n34)
         );
  NOR2_X1 sboxTI_g3_U19 ( .A1(sboxIn1[2]), .A2(md1Reg[3]), .ZN(sboxTI_g3_n36)
         );
  XNOR2_X1 sboxTI_g3_U18 ( .A(sboxIn1[0]), .B(sboxTI_g3_n33), .ZN(
        sboxTI_g3_n41) );
  XOR2_X1 sboxTI_g3_U17 ( .A(sboxTI_g3_n32), .B(sboxTI_g3_n31), .Z(
        sboxTI_g3_n33) );
  NAND2_X1 sboxTI_g3_U16 ( .A1(md1Reg[2]), .A2(sboxIn1[1]), .ZN(sboxTI_g3_n31)
         );
  NAND2_X1 sboxTI_g3_U15 ( .A1(md1Reg[1]), .A2(sboxIn1[2]), .ZN(sboxTI_g3_n32)
         );
  XNOR2_X1 sboxTI_g3_U14 ( .A(sboxTI_g3_n30), .B(sboxTI_g3_n29), .ZN(
        sboxTI_g3Out[1]) );
  XNOR2_X1 sboxTI_g3_U13 ( .A(sboxTI_g3_n28), .B(sboxTI_g3_n27), .ZN(
        sboxTI_g3_n29) );
  XOR2_X1 sboxTI_g3_U12 ( .A(sboxTI_g3_n26), .B(sboxTI_g3_n25), .Z(
        sboxTI_g3_n27) );
  NAND2_X1 sboxTI_g3_U11 ( .A1(sboxTI_g3_n37), .A2(sboxIn1[0]), .ZN(
        sboxTI_g3_n25) );
  XNOR2_X1 sboxTI_g3_U10 ( .A(sboxTI_g3_n24), .B(sboxTI_g3_n23), .ZN(
        sboxTI_g3_n37) );
  XOR2_X1 sboxTI_g3_U9 ( .A(sboxIn1[2]), .B(md1Reg[2]), .Z(sboxTI_g3_n23) );
  XNOR2_X1 sboxTI_g3_U8 ( .A(md1Reg[1]), .B(sboxIn1[1]), .ZN(sboxTI_g3_n24) );
  NAND2_X1 sboxTI_g3_U7 ( .A1(md1Reg[1]), .A2(md1Reg[2]), .ZN(sboxTI_g3_n26)
         );
  NOR2_X1 sboxTI_g3_U6 ( .A1(md1Reg[0]), .A2(sboxTI_g3_n22), .ZN(sboxTI_g3_n28) );
  XNOR2_X1 sboxTI_g3_U5 ( .A(sboxTI_g3_n21), .B(sboxTI_g3_n20), .ZN(
        sboxTI_g3_n30) );
  NAND2_X1 sboxTI_g3_U4 ( .A1(md1Reg[0]), .A2(sboxIn1[2]), .ZN(sboxTI_g3_n20)
         );
  XOR2_X1 sboxTI_g3_U3 ( .A(md1Reg[3]), .B(sboxTI_g3_C), .Z(sboxTI_g3_n21) );
  XNOR2_X1 sboxTI_g3_U2 ( .A(sboxTI_g3_n22), .B(sboxIn1[2]), .ZN(
        sboxTI_g3Out[2]) );
  INV_X1 sboxTI_g3_U1 ( .A(sboxIn1[1]), .ZN(sboxTI_g3_n22) );
  AND2_X1 sboxTI_g3_CtermInst_U1 ( .A1(sboxIn1[1]), .A2(sboxIn1[2]), .ZN(
        sboxTI_g3_C) );
  MUX2_X1 sboxTI_y3_U5 ( .A(sboxTI_g3Reg[3]), .B(sboxTI_g3Out[3]), .S(
        enSboxReg), .Z(sboxTI_y3_n13) );
  MUX2_X1 sboxTI_y3_U4 ( .A(sboxTI_g3Reg[1]), .B(sboxTI_g3Out[1]), .S(
        enSboxReg), .Z(sboxTI_y3_n11) );
  MUX2_X1 sboxTI_y3_U3 ( .A(sboxTI_g3Reg[2]), .B(sboxTI_g3Out[2]), .S(
        enSboxReg), .Z(sboxTI_y3_n12) );
  MUX2_X1 sboxTI_y3_U2 ( .A(sboxTI_g3Reg[0]), .B(sboxTI_g3Out[0]), .S(
        enSboxReg), .Z(sboxTI_y3_n10) );
  DFF_X1 sboxTI_y3_s_current_state_reg_0_ ( .D(sboxTI_y3_n10), .CK(clk), .Q(
        sboxTI_g3Reg[0]) , .QN() ); 
  DFF_X1 sboxTI_y3_s_current_state_reg_1_ ( .D(sboxTI_y3_n11), .CK(clk), .Q(
        sboxTI_g3Reg[1]) , .QN() ); 
  DFF_X1 sboxTI_y3_s_current_state_reg_2_ ( .D(sboxTI_y3_n12), .CK(clk), .Q(
        sboxTI_g3Reg[2]) , .QN() ); 
  DFF_X1 sboxTI_y3_s_current_state_reg_3_ ( .D(sboxTI_y3_n13), .CK(clk), .Q(
        sboxTI_g3Reg[3]) , .QN() ); 
  MUX2_X1 sboxTI_y2_U5 ( .A(sboxTI_g2Reg[3]), .B(sboxTI_g2Out[3]), .S(
        enSboxReg), .Z(sboxTI_y2_n14) );
  MUX2_X1 sboxTI_y2_U4 ( .A(sboxTI_g2Reg[2]), .B(sboxTI_g2Out[2]), .S(
        enSboxReg), .Z(sboxTI_y2_n15) );
  MUX2_X1 sboxTI_y2_U3 ( .A(sboxTI_g2Reg[1]), .B(sboxTI_g2Out[1]), .S(
        enSboxReg), .Z(sboxTI_y2_n16) );
  MUX2_X1 sboxTI_y2_U2 ( .A(sboxTI_g2Reg[0]), .B(sboxTI_g2Out[0]), .S(
        enSboxReg), .Z(sboxTI_y2_n17) );
  DFF_X1 sboxTI_y2_s_current_state_reg_0_ ( .D(sboxTI_y2_n17), .CK(clk), .Q(
        sboxTI_g2Reg[0]) , .QN() ); 
  DFF_X1 sboxTI_y2_s_current_state_reg_1_ ( .D(sboxTI_y2_n16), .CK(clk), .Q(
        sboxTI_g2Reg[1]) , .QN() ); 
  DFF_X1 sboxTI_y2_s_current_state_reg_2_ ( .D(sboxTI_y2_n15), .CK(clk), .Q(
        sboxTI_g2Reg[2]) , .QN() ); 
  DFF_X1 sboxTI_y2_s_current_state_reg_3_ ( .D(sboxTI_y2_n14), .CK(clk), .Q(
        sboxTI_g2Reg[3]) , .QN() ); 
  MUX2_X1 sboxTI_y1_U5 ( .A(sboxTI_g1Reg[3]), .B(sboxTI_g1Out[3]), .S(
        enSboxReg), .Z(sboxTI_y1_n14) );
  MUX2_X1 sboxTI_y1_U4 ( .A(sboxTI_g1Reg[2]), .B(sboxTI_g1Out[2]), .S(
        enSboxReg), .Z(sboxTI_y1_n15) );
  MUX2_X1 sboxTI_y1_U3 ( .A(sboxTI_g1Reg[1]), .B(sboxTI_g1Out[1]), .S(
        enSboxReg), .Z(sboxTI_y1_n16) );
  MUX2_X1 sboxTI_y1_U2 ( .A(sboxTI_g1Reg[0]), .B(sboxTI_g1Out[0]), .S(
        enSboxReg), .Z(sboxTI_y1_n17) );
  DFF_X1 sboxTI_y1_s_current_state_reg_0_ ( .D(sboxTI_y1_n17), .CK(clk), .Q(
        sboxTI_g1Reg[0]) , .QN() ); 
  DFF_X1 sboxTI_y1_s_current_state_reg_1_ ( .D(sboxTI_y1_n16), .CK(clk), .Q(
        sboxTI_g1Reg[1]) , .QN() ); 
  DFF_X1 sboxTI_y1_s_current_state_reg_2_ ( .D(sboxTI_y1_n15), .CK(clk), .Q(
        sboxTI_g1Reg[2]) , .QN() ); 
  DFF_X1 sboxTI_y1_s_current_state_reg_3_ ( .D(sboxTI_y1_n14), .CK(clk), .Q(
        sboxTI_g1Reg[3]) , .QN() ); 
DFF_X1 DoneReg_s_current_state_reg ( .D(final), .CK(clk), .Q(done) , .QN() );
  MUX2_X1 DataOutReg1_gff_U68 ( .A(data_out1[63]), .B(data_out1[59]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n193) );
  MUX2_X1 DataOutReg1_gff_U67 ( .A(data_out1[62]), .B(data_out1[58]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n192) );
  MUX2_X1 DataOutReg1_gff_U66 ( .A(data_out1[61]), .B(data_out1[57]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n191) );
  MUX2_X1 DataOutReg1_gff_U65 ( .A(data_out1[60]), .B(data_out1[56]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n190) );
  MUX2_X1 DataOutReg1_gff_U64 ( .A(data_out1[59]), .B(data_out1[55]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n189) );
  MUX2_X1 DataOutReg1_gff_U63 ( .A(data_out1[58]), .B(data_out1[54]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n188) );
  MUX2_X1 DataOutReg1_gff_U62 ( .A(data_out1[57]), .B(data_out1[53]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n187) );
  MUX2_X1 DataOutReg1_gff_U61 ( .A(data_out1[56]), .B(data_out1[52]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n186) );
  MUX2_X1 DataOutReg1_gff_U60 ( .A(data_out1[55]), .B(data_out1[51]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n185) );
  MUX2_X1 DataOutReg1_gff_U59 ( .A(data_out1[54]), .B(data_out1[50]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n184) );
  MUX2_X1 DataOutReg1_gff_U58 ( .A(data_out1[53]), .B(data_out1[49]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n183) );
  MUX2_X1 DataOutReg1_gff_U57 ( .A(data_out1[52]), .B(data_out1[48]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n182) );
  MUX2_X1 DataOutReg1_gff_U56 ( .A(data_out1[51]), .B(data_out1[47]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n181) );
  MUX2_X1 DataOutReg1_gff_U55 ( .A(data_out1[50]), .B(data_out1[46]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n180) );
  MUX2_X1 DataOutReg1_gff_U54 ( .A(data_out1[49]), .B(data_out1[45]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n179) );
  MUX2_X1 DataOutReg1_gff_U53 ( .A(data_out1[48]), .B(data_out1[44]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n178) );
  MUX2_X1 DataOutReg1_gff_U52 ( .A(data_out1[47]), .B(data_out1[43]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n177) );
  MUX2_X1 DataOutReg1_gff_U51 ( .A(data_out1[46]), .B(data_out1[42]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n176) );
  MUX2_X1 DataOutReg1_gff_U50 ( .A(data_out1[45]), .B(data_out1[41]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n175) );
  MUX2_X1 DataOutReg1_gff_U49 ( .A(data_out1[44]), .B(data_out1[40]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n174) );
  MUX2_X1 DataOutReg1_gff_U48 ( .A(data_out1[43]), .B(data_out1[39]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n173) );
  MUX2_X1 DataOutReg1_gff_U47 ( .A(data_out1[42]), .B(data_out1[38]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n172) );
  MUX2_X1 DataOutReg1_gff_U46 ( .A(data_out1[41]), .B(data_out1[37]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n171) );
  MUX2_X1 DataOutReg1_gff_U45 ( .A(data_out1[40]), .B(data_out1[36]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n170) );
  MUX2_X1 DataOutReg1_gff_U44 ( .A(data_out1[39]), .B(data_out1[35]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n169) );
  MUX2_X1 DataOutReg1_gff_U43 ( .A(data_out1[38]), .B(data_out1[34]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n168) );
  MUX2_X1 DataOutReg1_gff_U42 ( .A(data_out1[37]), .B(data_out1[33]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n167) );
  MUX2_X1 DataOutReg1_gff_U41 ( .A(data_out1[36]), .B(data_out1[32]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n166) );
  MUX2_X1 DataOutReg1_gff_U40 ( .A(data_out1[35]), .B(data_out1[31]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n165) );
  MUX2_X1 DataOutReg1_gff_U39 ( .A(data_out1[34]), .B(data_out1[30]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n164) );
  MUX2_X1 DataOutReg1_gff_U38 ( .A(data_out1[33]), .B(data_out1[29]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n163) );
  MUX2_X1 DataOutReg1_gff_U37 ( .A(data_out1[32]), .B(data_out1[28]), .S(
        intDone), .Z(DataOutReg1_gff_n162) );
  MUX2_X1 DataOutReg1_gff_U36 ( .A(data_out1[31]), .B(data_out1[27]), .S(
        intDone), .Z(DataOutReg1_gff_n161) );
  MUX2_X1 DataOutReg1_gff_U35 ( .A(data_out1[30]), .B(data_out1[26]), .S(
        intDone), .Z(DataOutReg1_gff_n160) );
  MUX2_X1 DataOutReg1_gff_U34 ( .A(data_out1[29]), .B(data_out1[25]), .S(
        intDone), .Z(DataOutReg1_gff_n159) );
  MUX2_X1 DataOutReg1_gff_U33 ( .A(data_out1[28]), .B(data_out1[24]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n158) );
  MUX2_X1 DataOutReg1_gff_U32 ( .A(data_out1[27]), .B(data_out1[23]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n157) );
  MUX2_X1 DataOutReg1_gff_U31 ( .A(data_out1[26]), .B(data_out1[22]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n156) );
  MUX2_X1 DataOutReg1_gff_U30 ( .A(data_out1[25]), .B(data_out1[21]), .S(
        intDone), .Z(DataOutReg1_gff_n155) );
  MUX2_X1 DataOutReg1_gff_U29 ( .A(data_out1[24]), .B(data_out1[20]), .S(
        intDone), .Z(DataOutReg1_gff_n154) );
  MUX2_X1 DataOutReg1_gff_U28 ( .A(data_out1[23]), .B(data_out1[19]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n153) );
  MUX2_X1 DataOutReg1_gff_U27 ( .A(data_out1[22]), .B(data_out1[18]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n152) );
  MUX2_X1 DataOutReg1_gff_U26 ( .A(data_out1[21]), .B(data_out1[17]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n151) );
  MUX2_X1 DataOutReg1_gff_U25 ( .A(data_out1[20]), .B(data_out1[16]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n150) );
  MUX2_X1 DataOutReg1_gff_U24 ( .A(data_out1[19]), .B(data_out1[15]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n149) );
  MUX2_X1 DataOutReg1_gff_U23 ( .A(data_out1[18]), .B(data_out1[14]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n148) );
  MUX2_X1 DataOutReg1_gff_U22 ( .A(data_out1[17]), .B(data_out1[13]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n147) );
  MUX2_X1 DataOutReg1_gff_U21 ( .A(data_out1[16]), .B(data_out1[12]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n146) );
  MUX2_X1 DataOutReg1_gff_U20 ( .A(data_out1[15]), .B(data_out1[11]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n145) );
  MUX2_X1 DataOutReg1_gff_U19 ( .A(data_out1[14]), .B(data_out1[10]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n144) );
  MUX2_X1 DataOutReg1_gff_U18 ( .A(data_out1[13]), .B(data_out1[9]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n143) );
  MUX2_X1 DataOutReg1_gff_U17 ( .A(data_out1[12]), .B(data_out1[8]), .S(
        DataOutReg1_gff_n200), .Z(DataOutReg1_gff_n142) );
  MUX2_X1 DataOutReg1_gff_U16 ( .A(data_out1[11]), .B(data_out1[7]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n141) );
  MUX2_X1 DataOutReg1_gff_U15 ( .A(data_out1[10]), .B(data_out1[6]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n140) );
  MUX2_X1 DataOutReg1_gff_U14 ( .A(data_out1[9]), .B(data_out1[5]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n139) );
  MUX2_X1 DataOutReg1_gff_U13 ( .A(data_out1[8]), .B(data_out1[4]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n138) );
  MUX2_X1 DataOutReg1_gff_U12 ( .A(data_out1[7]), .B(data_out1[3]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n137) );
  MUX2_X1 DataOutReg1_gff_U11 ( .A(data_out1[6]), .B(data_out1[2]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n136) );
  MUX2_X1 DataOutReg1_gff_U10 ( .A(data_out1[5]), .B(data_out1[1]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n135) );
  MUX2_X1 DataOutReg1_gff_U9 ( .A(data_out1[4]), .B(data_out1[0]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n134) );
  MUX2_X1 DataOutReg1_gff_U8 ( .A(data_out1[0]), .B(sboxIn1[0]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n130) );
  MUX2_X1 DataOutReg1_gff_U7 ( .A(data_out1[3]), .B(sboxIn1[3]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n133) );
  MUX2_X1 DataOutReg1_gff_U6 ( .A(data_out1[2]), .B(sboxIn1[2]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n132) );
  MUX2_X1 DataOutReg1_gff_U5 ( .A(data_out1[1]), .B(sboxIn1[1]), .S(
        DataOutReg1_gff_n199), .Z(DataOutReg1_gff_n131) );
  INV_X2 DataOutReg1_gff_U4 ( .A(DataOutReg1_gff_n198), .ZN(
        DataOutReg1_gff_n199) );
  INV_X1 DataOutReg1_gff_U3 ( .A(DataOutReg1_gff_n198), .ZN(
        DataOutReg1_gff_n200) );
  INV_X1 DataOutReg1_gff_U2 ( .A(intDone), .ZN(DataOutReg1_gff_n198) );
  DFF_X1 DataOutReg1_gff_s_current_state_reg_0_ ( .D(DataOutReg1_gff_n130), 
        .CK(clk), .Q(data_out1[0]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_1_ ( .D(DataOutReg1_gff_n131), 
        .CK(clk), .Q(data_out1[1]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_2_ ( .D(DataOutReg1_gff_n132), 
        .CK(clk), .Q(data_out1[2]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_3_ ( .D(DataOutReg1_gff_n133), 
        .CK(clk), .Q(data_out1[3]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_4_ ( .D(DataOutReg1_gff_n134), 
        .CK(clk), .Q(data_out1[4]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_5_ ( .D(DataOutReg1_gff_n135), 
        .CK(clk), .Q(data_out1[5]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_6_ ( .D(DataOutReg1_gff_n136), 
        .CK(clk), .Q(data_out1[6]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_7_ ( .D(DataOutReg1_gff_n137), 
        .CK(clk), .Q(data_out1[7]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_8_ ( .D(DataOutReg1_gff_n138), 
        .CK(clk), .Q(data_out1[8]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_9_ ( .D(DataOutReg1_gff_n139), 
        .CK(clk), .Q(data_out1[9]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_10_ ( .D(DataOutReg1_gff_n140), 
        .CK(clk), .Q(data_out1[10]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_11_ ( .D(DataOutReg1_gff_n141), 
        .CK(clk), .Q(data_out1[11]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_12_ ( .D(DataOutReg1_gff_n142), 
        .CK(clk), .Q(data_out1[12]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_13_ ( .D(DataOutReg1_gff_n143), 
        .CK(clk), .Q(data_out1[13]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_14_ ( .D(DataOutReg1_gff_n144), 
        .CK(clk), .Q(data_out1[14]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_15_ ( .D(DataOutReg1_gff_n145), 
        .CK(clk), .Q(data_out1[15]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_16_ ( .D(DataOutReg1_gff_n146), 
        .CK(clk), .Q(data_out1[16]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_17_ ( .D(DataOutReg1_gff_n147), 
        .CK(clk), .Q(data_out1[17]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_18_ ( .D(DataOutReg1_gff_n148), 
        .CK(clk), .Q(data_out1[18]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_19_ ( .D(DataOutReg1_gff_n149), 
        .CK(clk), .Q(data_out1[19]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_20_ ( .D(DataOutReg1_gff_n150), 
        .CK(clk), .Q(data_out1[20]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_21_ ( .D(DataOutReg1_gff_n151), 
        .CK(clk), .Q(data_out1[21]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_22_ ( .D(DataOutReg1_gff_n152), 
        .CK(clk), .Q(data_out1[22]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_23_ ( .D(DataOutReg1_gff_n153), 
        .CK(clk), .Q(data_out1[23]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_24_ ( .D(DataOutReg1_gff_n154), 
        .CK(clk), .Q(data_out1[24]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_25_ ( .D(DataOutReg1_gff_n155), 
        .CK(clk), .Q(data_out1[25]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_26_ ( .D(DataOutReg1_gff_n156), 
        .CK(clk), .Q(data_out1[26]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_27_ ( .D(DataOutReg1_gff_n157), 
        .CK(clk), .Q(data_out1[27]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_28_ ( .D(DataOutReg1_gff_n158), 
        .CK(clk), .Q(data_out1[28]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_29_ ( .D(DataOutReg1_gff_n159), 
        .CK(clk), .Q(data_out1[29]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_30_ ( .D(DataOutReg1_gff_n160), 
        .CK(clk), .Q(data_out1[30]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_31_ ( .D(DataOutReg1_gff_n161), 
        .CK(clk), .Q(data_out1[31]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_32_ ( .D(DataOutReg1_gff_n162), 
        .CK(clk), .Q(data_out1[32]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_33_ ( .D(DataOutReg1_gff_n163), 
        .CK(clk), .Q(data_out1[33]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_34_ ( .D(DataOutReg1_gff_n164), 
        .CK(clk), .Q(data_out1[34]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_35_ ( .D(DataOutReg1_gff_n165), 
        .CK(clk), .Q(data_out1[35]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_36_ ( .D(DataOutReg1_gff_n166), 
        .CK(clk), .Q(data_out1[36]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_37_ ( .D(DataOutReg1_gff_n167), 
        .CK(clk), .Q(data_out1[37]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_38_ ( .D(DataOutReg1_gff_n168), 
        .CK(clk), .Q(data_out1[38]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_39_ ( .D(DataOutReg1_gff_n169), 
        .CK(clk), .Q(data_out1[39]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_40_ ( .D(DataOutReg1_gff_n170), 
        .CK(clk), .Q(data_out1[40]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_41_ ( .D(DataOutReg1_gff_n171), 
        .CK(clk), .Q(data_out1[41]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_42_ ( .D(DataOutReg1_gff_n172), 
        .CK(clk), .Q(data_out1[42]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_43_ ( .D(DataOutReg1_gff_n173), 
        .CK(clk), .Q(data_out1[43]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_44_ ( .D(DataOutReg1_gff_n174), 
        .CK(clk), .Q(data_out1[44]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_45_ ( .D(DataOutReg1_gff_n175), 
        .CK(clk), .Q(data_out1[45]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_46_ ( .D(DataOutReg1_gff_n176), 
        .CK(clk), .Q(data_out1[46]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_47_ ( .D(DataOutReg1_gff_n177), 
        .CK(clk), .Q(data_out1[47]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_48_ ( .D(DataOutReg1_gff_n178), 
        .CK(clk), .Q(data_out1[48]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_49_ ( .D(DataOutReg1_gff_n179), 
        .CK(clk), .Q(data_out1[49]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_50_ ( .D(DataOutReg1_gff_n180), 
        .CK(clk), .Q(data_out1[50]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_51_ ( .D(DataOutReg1_gff_n181), 
        .CK(clk), .Q(data_out1[51]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_52_ ( .D(DataOutReg1_gff_n182), 
        .CK(clk), .Q(data_out1[52]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_53_ ( .D(DataOutReg1_gff_n183), 
        .CK(clk), .Q(data_out1[53]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_54_ ( .D(DataOutReg1_gff_n184), 
        .CK(clk), .Q(data_out1[54]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_55_ ( .D(DataOutReg1_gff_n185), 
        .CK(clk), .Q(data_out1[55]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_56_ ( .D(DataOutReg1_gff_n186), 
        .CK(clk), .Q(data_out1[56]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_57_ ( .D(DataOutReg1_gff_n187), 
        .CK(clk), .Q(data_out1[57]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_58_ ( .D(DataOutReg1_gff_n188), 
        .CK(clk), .Q(data_out1[58]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_59_ ( .D(DataOutReg1_gff_n189), 
        .CK(clk), .Q(data_out1[59]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_60_ ( .D(DataOutReg1_gff_n190), 
        .CK(clk), .Q(data_out1[60]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_61_ ( .D(DataOutReg1_gff_n191), 
        .CK(clk), .Q(data_out1[61]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_62_ ( .D(DataOutReg1_gff_n192), 
        .CK(clk), .Q(data_out1[62]) , .QN() ); 
  DFF_X1 DataOutReg1_gff_s_current_state_reg_63_ ( .D(DataOutReg1_gff_n193), 
        .CK(clk), .Q(data_out1[63]) , .QN() ); 
  MUX2_X1 DataOutReg2_gff_U67 ( .A(data_out2[63]), .B(data_out2[59]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n199) );
  MUX2_X1 DataOutReg2_gff_U66 ( .A(data_out2[62]), .B(data_out2[58]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n200) );
  MUX2_X1 DataOutReg2_gff_U65 ( .A(data_out2[61]), .B(data_out2[57]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n201) );
  MUX2_X1 DataOutReg2_gff_U64 ( .A(data_out2[60]), .B(data_out2[56]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n202) );
  MUX2_X1 DataOutReg2_gff_U63 ( .A(data_out2[59]), .B(data_out2[55]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n203) );
  MUX2_X1 DataOutReg2_gff_U62 ( .A(data_out2[58]), .B(data_out2[54]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n204) );
  MUX2_X1 DataOutReg2_gff_U61 ( .A(data_out2[57]), .B(data_out2[53]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n205) );
  MUX2_X1 DataOutReg2_gff_U60 ( .A(data_out2[56]), .B(data_out2[52]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n206) );
  MUX2_X1 DataOutReg2_gff_U59 ( .A(data_out2[55]), .B(data_out2[51]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n207) );
  MUX2_X1 DataOutReg2_gff_U58 ( .A(data_out2[54]), .B(data_out2[50]), .S(
        intDone), .Z(DataOutReg2_gff_n208) );
  MUX2_X1 DataOutReg2_gff_U57 ( .A(data_out2[53]), .B(data_out2[49]), .S(
        intDone), .Z(DataOutReg2_gff_n209) );
  MUX2_X1 DataOutReg2_gff_U56 ( .A(data_out2[52]), .B(data_out2[48]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n210) );
  MUX2_X1 DataOutReg2_gff_U55 ( .A(data_out2[51]), .B(data_out2[47]), .S(
        intDone), .Z(DataOutReg2_gff_n211) );
  MUX2_X1 DataOutReg2_gff_U54 ( .A(data_out2[50]), .B(data_out2[46]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n212) );
  MUX2_X1 DataOutReg2_gff_U53 ( .A(data_out2[49]), .B(data_out2[45]), .S(
        intDone), .Z(DataOutReg2_gff_n213) );
  MUX2_X1 DataOutReg2_gff_U52 ( .A(data_out2[48]), .B(data_out2[44]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n214) );
  MUX2_X1 DataOutReg2_gff_U51 ( .A(data_out2[47]), .B(data_out2[43]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n215) );
  MUX2_X1 DataOutReg2_gff_U50 ( .A(data_out2[46]), .B(data_out2[42]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n216) );
  MUX2_X1 DataOutReg2_gff_U49 ( .A(data_out2[45]), .B(data_out2[41]), .S(
        intDone), .Z(DataOutReg2_gff_n217) );
  MUX2_X1 DataOutReg2_gff_U48 ( .A(data_out2[44]), .B(data_out2[40]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n218) );
  MUX2_X1 DataOutReg2_gff_U47 ( .A(data_out2[43]), .B(data_out2[39]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n219) );
  MUX2_X1 DataOutReg2_gff_U46 ( .A(data_out2[42]), .B(data_out2[38]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n220) );
  MUX2_X1 DataOutReg2_gff_U45 ( .A(data_out2[41]), .B(data_out2[37]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n221) );
  MUX2_X1 DataOutReg2_gff_U44 ( .A(data_out2[40]), .B(data_out2[36]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n222) );
  MUX2_X1 DataOutReg2_gff_U43 ( .A(data_out2[39]), .B(data_out2[35]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n223) );
  MUX2_X1 DataOutReg2_gff_U42 ( .A(data_out2[38]), .B(data_out2[34]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n224) );
  MUX2_X1 DataOutReg2_gff_U41 ( .A(data_out2[37]), .B(data_out2[33]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n225) );
  MUX2_X1 DataOutReg2_gff_U40 ( .A(data_out2[36]), .B(data_out2[32]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n226) );
  MUX2_X1 DataOutReg2_gff_U39 ( .A(data_out2[35]), .B(data_out2[31]), .S(
        intDone), .Z(DataOutReg2_gff_n227) );
  MUX2_X1 DataOutReg2_gff_U38 ( .A(data_out2[34]), .B(data_out2[30]), .S(
        intDone), .Z(DataOutReg2_gff_n228) );
  MUX2_X1 DataOutReg2_gff_U37 ( .A(data_out2[33]), .B(data_out2[29]), .S(
        intDone), .Z(DataOutReg2_gff_n229) );
  MUX2_X1 DataOutReg2_gff_U36 ( .A(data_out2[32]), .B(data_out2[28]), .S(
        intDone), .Z(DataOutReg2_gff_n230) );
  MUX2_X1 DataOutReg2_gff_U35 ( .A(data_out2[31]), .B(data_out2[27]), .S(
        intDone), .Z(DataOutReg2_gff_n231) );
  MUX2_X1 DataOutReg2_gff_U34 ( .A(data_out2[30]), .B(data_out2[26]), .S(
        intDone), .Z(DataOutReg2_gff_n232) );
  MUX2_X1 DataOutReg2_gff_U33 ( .A(data_out2[29]), .B(data_out2[25]), .S(
        intDone), .Z(DataOutReg2_gff_n233) );
  MUX2_X1 DataOutReg2_gff_U32 ( .A(data_out2[28]), .B(data_out2[24]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n234) );
  MUX2_X1 DataOutReg2_gff_U31 ( .A(data_out2[27]), .B(data_out2[23]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n235) );
  MUX2_X1 DataOutReg2_gff_U30 ( .A(data_out2[26]), .B(data_out2[22]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n236) );
  MUX2_X1 DataOutReg2_gff_U29 ( .A(data_out2[25]), .B(data_out2[21]), .S(
        intDone), .Z(DataOutReg2_gff_n237) );
  MUX2_X1 DataOutReg2_gff_U28 ( .A(data_out2[24]), .B(data_out2[20]), .S(
        intDone), .Z(DataOutReg2_gff_n238) );
  MUX2_X1 DataOutReg2_gff_U27 ( .A(data_out2[23]), .B(data_out2[19]), .S(
        intDone), .Z(DataOutReg2_gff_n239) );
  MUX2_X1 DataOutReg2_gff_U26 ( .A(data_out2[22]), .B(data_out2[18]), .S(
        intDone), .Z(DataOutReg2_gff_n240) );
  MUX2_X1 DataOutReg2_gff_U25 ( .A(data_out2[21]), .B(data_out2[17]), .S(
        intDone), .Z(DataOutReg2_gff_n241) );
  MUX2_X1 DataOutReg2_gff_U24 ( .A(data_out2[20]), .B(data_out2[16]), .S(
        intDone), .Z(DataOutReg2_gff_n242) );
  MUX2_X1 DataOutReg2_gff_U23 ( .A(data_out2[19]), .B(data_out2[15]), .S(
        intDone), .Z(DataOutReg2_gff_n243) );
  MUX2_X1 DataOutReg2_gff_U22 ( .A(data_out2[18]), .B(data_out2[14]), .S(
        intDone), .Z(DataOutReg2_gff_n244) );
  MUX2_X1 DataOutReg2_gff_U21 ( .A(data_out2[17]), .B(data_out2[13]), .S(
        intDone), .Z(DataOutReg2_gff_n245) );
  MUX2_X1 DataOutReg2_gff_U20 ( .A(data_out2[16]), .B(data_out2[12]), .S(
        intDone), .Z(DataOutReg2_gff_n246) );
  MUX2_X1 DataOutReg2_gff_U19 ( .A(data_out2[15]), .B(data_out2[11]), .S(
        intDone), .Z(DataOutReg2_gff_n247) );
  MUX2_X1 DataOutReg2_gff_U18 ( .A(data_out2[14]), .B(data_out2[10]), .S(
        intDone), .Z(DataOutReg2_gff_n248) );
  MUX2_X1 DataOutReg2_gff_U17 ( .A(data_out2[13]), .B(data_out2[9]), .S(
        intDone), .Z(DataOutReg2_gff_n249) );
  MUX2_X1 DataOutReg2_gff_U16 ( .A(data_out2[12]), .B(data_out2[8]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n250) );
  MUX2_X1 DataOutReg2_gff_U15 ( .A(data_out2[11]), .B(data_out2[7]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n251) );
  MUX2_X1 DataOutReg2_gff_U14 ( .A(data_out2[10]), .B(data_out2[6]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n252) );
  MUX2_X1 DataOutReg2_gff_U13 ( .A(data_out2[9]), .B(data_out2[5]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n253) );
  MUX2_X1 DataOutReg2_gff_U12 ( .A(data_out2[8]), .B(data_out2[4]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n254) );
  MUX2_X1 DataOutReg2_gff_U11 ( .A(data_out2[7]), .B(data_out2[3]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n255) );
  MUX2_X1 DataOutReg2_gff_U10 ( .A(data_out2[6]), .B(data_out2[2]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n256) );
  MUX2_X1 DataOutReg2_gff_U9 ( .A(data_out2[5]), .B(data_out2[1]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n257) );
  MUX2_X1 DataOutReg2_gff_U8 ( .A(data_out2[4]), .B(data_out2[0]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n258) );
  MUX2_X1 DataOutReg2_gff_U7 ( .A(data_out2[0]), .B(md1Reg[0]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n262) );
  MUX2_X1 DataOutReg2_gff_U6 ( .A(data_out2[3]), .B(md1Reg[3]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n259) );
  MUX2_X1 DataOutReg2_gff_U5 ( .A(data_out2[2]), .B(md1Reg[2]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n260) );
  MUX2_X1 DataOutReg2_gff_U4 ( .A(data_out2[1]), .B(md1Reg[1]), .S(
        DataOutReg2_gff_n392), .Z(DataOutReg2_gff_n261) );
  INV_X2 DataOutReg2_gff_U3 ( .A(DataOutReg2_gff_n391), .ZN(
        DataOutReg2_gff_n392) );
  INV_X1 DataOutReg2_gff_U2 ( .A(intDone), .ZN(DataOutReg2_gff_n391) );
  DFF_X1 DataOutReg2_gff_s_current_state_reg_0_ ( .D(DataOutReg2_gff_n262), 
        .CK(clk), .Q(data_out2[0]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_1_ ( .D(DataOutReg2_gff_n261), 
        .CK(clk), .Q(data_out2[1]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_2_ ( .D(DataOutReg2_gff_n260), 
        .CK(clk), .Q(data_out2[2]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_3_ ( .D(DataOutReg2_gff_n259), 
        .CK(clk), .Q(data_out2[3]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_4_ ( .D(DataOutReg2_gff_n258), 
        .CK(clk), .Q(data_out2[4]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_5_ ( .D(DataOutReg2_gff_n257), 
        .CK(clk), .Q(data_out2[5]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_6_ ( .D(DataOutReg2_gff_n256), 
        .CK(clk), .Q(data_out2[6]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_7_ ( .D(DataOutReg2_gff_n255), 
        .CK(clk), .Q(data_out2[7]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_8_ ( .D(DataOutReg2_gff_n254), 
        .CK(clk), .Q(data_out2[8]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_9_ ( .D(DataOutReg2_gff_n253), 
        .CK(clk), .Q(data_out2[9]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_10_ ( .D(DataOutReg2_gff_n252), 
        .CK(clk), .Q(data_out2[10]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_11_ ( .D(DataOutReg2_gff_n251), 
        .CK(clk), .Q(data_out2[11]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_12_ ( .D(DataOutReg2_gff_n250), 
        .CK(clk), .Q(data_out2[12]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_13_ ( .D(DataOutReg2_gff_n249), 
        .CK(clk), .Q(data_out2[13]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_14_ ( .D(DataOutReg2_gff_n248), 
        .CK(clk), .Q(data_out2[14]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_15_ ( .D(DataOutReg2_gff_n247), 
        .CK(clk), .Q(data_out2[15]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_16_ ( .D(DataOutReg2_gff_n246), 
        .CK(clk), .Q(data_out2[16]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_17_ ( .D(DataOutReg2_gff_n245), 
        .CK(clk), .Q(data_out2[17]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_18_ ( .D(DataOutReg2_gff_n244), 
        .CK(clk), .Q(data_out2[18]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_19_ ( .D(DataOutReg2_gff_n243), 
        .CK(clk), .Q(data_out2[19]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_20_ ( .D(DataOutReg2_gff_n242), 
        .CK(clk), .Q(data_out2[20]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_21_ ( .D(DataOutReg2_gff_n241), 
        .CK(clk), .Q(data_out2[21]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_22_ ( .D(DataOutReg2_gff_n240), 
        .CK(clk), .Q(data_out2[22]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_23_ ( .D(DataOutReg2_gff_n239), 
        .CK(clk), .Q(data_out2[23]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_24_ ( .D(DataOutReg2_gff_n238), 
        .CK(clk), .Q(data_out2[24]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_25_ ( .D(DataOutReg2_gff_n237), 
        .CK(clk), .Q(data_out2[25]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_26_ ( .D(DataOutReg2_gff_n236), 
        .CK(clk), .Q(data_out2[26]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_27_ ( .D(DataOutReg2_gff_n235), 
        .CK(clk), .Q(data_out2[27]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_28_ ( .D(DataOutReg2_gff_n234), 
        .CK(clk), .Q(data_out2[28]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_29_ ( .D(DataOutReg2_gff_n233), 
        .CK(clk), .Q(data_out2[29]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_30_ ( .D(DataOutReg2_gff_n232), 
        .CK(clk), .Q(data_out2[30]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_31_ ( .D(DataOutReg2_gff_n231), 
        .CK(clk), .Q(data_out2[31]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_32_ ( .D(DataOutReg2_gff_n230), 
        .CK(clk), .Q(data_out2[32]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_33_ ( .D(DataOutReg2_gff_n229), 
        .CK(clk), .Q(data_out2[33]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_34_ ( .D(DataOutReg2_gff_n228), 
        .CK(clk), .Q(data_out2[34]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_35_ ( .D(DataOutReg2_gff_n227), 
        .CK(clk), .Q(data_out2[35]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_36_ ( .D(DataOutReg2_gff_n226), 
        .CK(clk), .Q(data_out2[36]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_37_ ( .D(DataOutReg2_gff_n225), 
        .CK(clk), .Q(data_out2[37]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_38_ ( .D(DataOutReg2_gff_n224), 
        .CK(clk), .Q(data_out2[38]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_39_ ( .D(DataOutReg2_gff_n223), 
        .CK(clk), .Q(data_out2[39]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_40_ ( .D(DataOutReg2_gff_n222), 
        .CK(clk), .Q(data_out2[40]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_41_ ( .D(DataOutReg2_gff_n221), 
        .CK(clk), .Q(data_out2[41]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_42_ ( .D(DataOutReg2_gff_n220), 
        .CK(clk), .Q(data_out2[42]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_43_ ( .D(DataOutReg2_gff_n219), 
        .CK(clk), .Q(data_out2[43]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_44_ ( .D(DataOutReg2_gff_n218), 
        .CK(clk), .Q(data_out2[44]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_45_ ( .D(DataOutReg2_gff_n217), 
        .CK(clk), .Q(data_out2[45]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_46_ ( .D(DataOutReg2_gff_n216), 
        .CK(clk), .Q(data_out2[46]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_47_ ( .D(DataOutReg2_gff_n215), 
        .CK(clk), .Q(data_out2[47]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_48_ ( .D(DataOutReg2_gff_n214), 
        .CK(clk), .Q(data_out2[48]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_49_ ( .D(DataOutReg2_gff_n213), 
        .CK(clk), .Q(data_out2[49]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_50_ ( .D(DataOutReg2_gff_n212), 
        .CK(clk), .Q(data_out2[50]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_51_ ( .D(DataOutReg2_gff_n211), 
        .CK(clk), .Q(data_out2[51]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_52_ ( .D(DataOutReg2_gff_n210), 
        .CK(clk), .Q(data_out2[52]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_53_ ( .D(DataOutReg2_gff_n209), 
        .CK(clk), .Q(data_out2[53]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_54_ ( .D(DataOutReg2_gff_n208), 
        .CK(clk), .Q(data_out2[54]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_55_ ( .D(DataOutReg2_gff_n207), 
        .CK(clk), .Q(data_out2[55]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_56_ ( .D(DataOutReg2_gff_n206), 
        .CK(clk), .Q(data_out2[56]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_57_ ( .D(DataOutReg2_gff_n205), 
        .CK(clk), .Q(data_out2[57]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_58_ ( .D(DataOutReg2_gff_n204), 
        .CK(clk), .Q(data_out2[58]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_59_ ( .D(DataOutReg2_gff_n203), 
        .CK(clk), .Q(data_out2[59]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_60_ ( .D(DataOutReg2_gff_n202), 
        .CK(clk), .Q(data_out2[60]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_61_ ( .D(DataOutReg2_gff_n201), 
        .CK(clk), .Q(data_out2[61]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_62_ ( .D(DataOutReg2_gff_n200), 
        .CK(clk), .Q(data_out2[62]) , .QN() ); 
  DFF_X1 DataOutReg2_gff_s_current_state_reg_63_ ( .D(DataOutReg2_gff_n199), 
        .CK(clk), .Q(data_out2[63]) , .QN() ); 
  MUX2_X1 DataOutReg3_gff_U68 ( .A(data_out3[63]), .B(data_out3[59]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n199) );
  MUX2_X1 DataOutReg3_gff_U67 ( .A(data_out3[62]), .B(data_out3[58]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n200) );
  MUX2_X1 DataOutReg3_gff_U66 ( .A(data_out3[61]), .B(data_out3[57]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n201) );
  MUX2_X1 DataOutReg3_gff_U65 ( .A(data_out3[60]), .B(data_out3[56]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n202) );
  MUX2_X1 DataOutReg3_gff_U64 ( .A(data_out3[59]), .B(data_out3[55]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n203) );
  MUX2_X1 DataOutReg3_gff_U63 ( .A(data_out3[58]), .B(data_out3[54]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n204) );
  MUX2_X1 DataOutReg3_gff_U62 ( .A(data_out3[57]), .B(data_out3[53]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n205) );
  MUX2_X1 DataOutReg3_gff_U61 ( .A(data_out3[56]), .B(data_out3[52]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n206) );
  MUX2_X1 DataOutReg3_gff_U60 ( .A(data_out3[55]), .B(data_out3[51]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n207) );
  MUX2_X1 DataOutReg3_gff_U59 ( .A(data_out3[54]), .B(data_out3[50]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n208) );
  MUX2_X1 DataOutReg3_gff_U58 ( .A(data_out3[53]), .B(data_out3[49]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n209) );
  MUX2_X1 DataOutReg3_gff_U57 ( .A(data_out3[52]), .B(data_out3[48]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n210) );
  MUX2_X1 DataOutReg3_gff_U56 ( .A(data_out3[51]), .B(data_out3[47]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n211) );
  MUX2_X1 DataOutReg3_gff_U55 ( .A(data_out3[50]), .B(data_out3[46]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n212) );
  MUX2_X1 DataOutReg3_gff_U54 ( .A(data_out3[49]), .B(data_out3[45]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n213) );
  MUX2_X1 DataOutReg3_gff_U53 ( .A(data_out3[48]), .B(data_out3[44]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n214) );
  MUX2_X1 DataOutReg3_gff_U52 ( .A(data_out3[47]), .B(data_out3[43]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n215) );
  MUX2_X1 DataOutReg3_gff_U51 ( .A(data_out3[46]), .B(data_out3[42]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n216) );
  MUX2_X1 DataOutReg3_gff_U50 ( .A(data_out3[45]), .B(data_out3[41]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n217) );
  MUX2_X1 DataOutReg3_gff_U49 ( .A(data_out3[44]), .B(data_out3[40]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n218) );
  MUX2_X1 DataOutReg3_gff_U48 ( .A(data_out3[43]), .B(data_out3[39]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n219) );
  MUX2_X1 DataOutReg3_gff_U47 ( .A(data_out3[42]), .B(data_out3[38]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n220) );
  MUX2_X1 DataOutReg3_gff_U46 ( .A(data_out3[41]), .B(data_out3[37]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n221) );
  MUX2_X1 DataOutReg3_gff_U45 ( .A(data_out3[40]), .B(data_out3[36]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n222) );
  MUX2_X1 DataOutReg3_gff_U44 ( .A(data_out3[39]), .B(data_out3[35]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n223) );
  MUX2_X1 DataOutReg3_gff_U43 ( .A(data_out3[38]), .B(data_out3[34]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n224) );
  MUX2_X1 DataOutReg3_gff_U42 ( .A(data_out3[37]), .B(data_out3[33]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n225) );
  MUX2_X1 DataOutReg3_gff_U41 ( .A(data_out3[36]), .B(data_out3[32]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n226) );
  MUX2_X1 DataOutReg3_gff_U40 ( .A(data_out3[35]), .B(data_out3[31]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n227) );
  MUX2_X1 DataOutReg3_gff_U39 ( .A(data_out3[34]), .B(data_out3[30]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n228) );
  MUX2_X1 DataOutReg3_gff_U38 ( .A(data_out3[33]), .B(data_out3[29]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n229) );
  MUX2_X1 DataOutReg3_gff_U37 ( .A(data_out3[32]), .B(data_out3[28]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n230) );
  MUX2_X1 DataOutReg3_gff_U36 ( .A(data_out3[31]), .B(data_out3[27]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n231) );
  MUX2_X1 DataOutReg3_gff_U35 ( .A(data_out3[30]), .B(data_out3[26]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n232) );
  MUX2_X1 DataOutReg3_gff_U34 ( .A(data_out3[29]), .B(data_out3[25]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n233) );
  MUX2_X1 DataOutReg3_gff_U33 ( .A(data_out3[28]), .B(data_out3[24]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n234) );
  MUX2_X1 DataOutReg3_gff_U32 ( .A(data_out3[27]), .B(data_out3[23]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n235) );
  MUX2_X1 DataOutReg3_gff_U31 ( .A(data_out3[26]), .B(data_out3[22]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n236) );
  MUX2_X1 DataOutReg3_gff_U30 ( .A(data_out3[25]), .B(data_out3[21]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n237) );
  MUX2_X1 DataOutReg3_gff_U29 ( .A(data_out3[24]), .B(data_out3[20]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n238) );
  MUX2_X1 DataOutReg3_gff_U28 ( .A(data_out3[23]), .B(data_out3[19]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n239) );
  MUX2_X1 DataOutReg3_gff_U27 ( .A(data_out3[22]), .B(data_out3[18]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n240) );
  MUX2_X1 DataOutReg3_gff_U26 ( .A(data_out3[21]), .B(data_out3[17]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n241) );
  MUX2_X1 DataOutReg3_gff_U25 ( .A(data_out3[20]), .B(data_out3[16]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n242) );
  MUX2_X1 DataOutReg3_gff_U24 ( .A(data_out3[19]), .B(data_out3[15]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n243) );
  MUX2_X1 DataOutReg3_gff_U23 ( .A(data_out3[18]), .B(data_out3[14]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n244) );
  MUX2_X1 DataOutReg3_gff_U22 ( .A(data_out3[17]), .B(data_out3[13]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n245) );
  MUX2_X1 DataOutReg3_gff_U21 ( .A(data_out3[16]), .B(data_out3[12]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n246) );
  MUX2_X1 DataOutReg3_gff_U20 ( .A(data_out3[15]), .B(data_out3[11]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n247) );
  MUX2_X1 DataOutReg3_gff_U19 ( .A(data_out3[14]), .B(data_out3[10]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n248) );
  MUX2_X1 DataOutReg3_gff_U18 ( .A(data_out3[13]), .B(data_out3[9]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n249) );
  MUX2_X1 DataOutReg3_gff_U17 ( .A(data_out3[12]), .B(data_out3[8]), .S(
        DataOutReg3_gff_n392), .Z(DataOutReg3_gff_n250) );
  MUX2_X1 DataOutReg3_gff_U16 ( .A(data_out3[11]), .B(data_out3[7]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n251) );
  MUX2_X1 DataOutReg3_gff_U15 ( .A(data_out3[10]), .B(data_out3[6]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n252) );
  MUX2_X1 DataOutReg3_gff_U14 ( .A(data_out3[9]), .B(data_out3[5]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n253) );
  MUX2_X1 DataOutReg3_gff_U13 ( .A(data_out3[8]), .B(data_out3[4]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n254) );
  MUX2_X1 DataOutReg3_gff_U12 ( .A(data_out3[7]), .B(data_out3[3]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n255) );
  MUX2_X1 DataOutReg3_gff_U11 ( .A(data_out3[6]), .B(data_out3[2]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n256) );
  MUX2_X1 DataOutReg3_gff_U10 ( .A(data_out3[5]), .B(data_out3[1]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n257) );
  MUX2_X1 DataOutReg3_gff_U9 ( .A(data_out3[4]), .B(data_out3[0]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n258) );
  MUX2_X1 DataOutReg3_gff_U8 ( .A(data_out3[0]), .B(md2Reg[0]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n262) );
  MUX2_X1 DataOutReg3_gff_U7 ( .A(data_out3[3]), .B(md2Reg[3]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n259) );
  MUX2_X1 DataOutReg3_gff_U6 ( .A(data_out3[2]), .B(md2Reg[2]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n260) );
  MUX2_X1 DataOutReg3_gff_U5 ( .A(data_out3[1]), .B(md2Reg[1]), .S(
        DataOutReg3_gff_n393), .Z(DataOutReg3_gff_n261) );
  INV_X2 DataOutReg3_gff_U4 ( .A(DataOutReg3_gff_n391), .ZN(
        DataOutReg3_gff_n392) );
  INV_X1 DataOutReg3_gff_U3 ( .A(intDone), .ZN(DataOutReg3_gff_n391) );
  INV_X2 DataOutReg3_gff_U2 ( .A(DataOutReg3_gff_n391), .ZN(
        DataOutReg3_gff_n393) );
  DFF_X1 DataOutReg3_gff_s_current_state_reg_0_ ( .D(DataOutReg3_gff_n262), 
        .CK(clk), .Q(data_out3[0]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_1_ ( .D(DataOutReg3_gff_n261), 
        .CK(clk), .Q(data_out3[1]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_2_ ( .D(DataOutReg3_gff_n260), 
        .CK(clk), .Q(data_out3[2]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_3_ ( .D(DataOutReg3_gff_n259), 
        .CK(clk), .Q(data_out3[3]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_4_ ( .D(DataOutReg3_gff_n258), 
        .CK(clk), .Q(data_out3[4]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_5_ ( .D(DataOutReg3_gff_n257), 
        .CK(clk), .Q(data_out3[5]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_6_ ( .D(DataOutReg3_gff_n256), 
        .CK(clk), .Q(data_out3[6]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_7_ ( .D(DataOutReg3_gff_n255), 
        .CK(clk), .Q(data_out3[7]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_8_ ( .D(DataOutReg3_gff_n254), 
        .CK(clk), .Q(data_out3[8]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_9_ ( .D(DataOutReg3_gff_n253), 
        .CK(clk), .Q(data_out3[9]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_10_ ( .D(DataOutReg3_gff_n252), 
        .CK(clk), .Q(data_out3[10]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_11_ ( .D(DataOutReg3_gff_n251), 
        .CK(clk), .Q(data_out3[11]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_12_ ( .D(DataOutReg3_gff_n250), 
        .CK(clk), .Q(data_out3[12]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_13_ ( .D(DataOutReg3_gff_n249), 
        .CK(clk), .Q(data_out3[13]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_14_ ( .D(DataOutReg3_gff_n248), 
        .CK(clk), .Q(data_out3[14]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_15_ ( .D(DataOutReg3_gff_n247), 
        .CK(clk), .Q(data_out3[15]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_16_ ( .D(DataOutReg3_gff_n246), 
        .CK(clk), .Q(data_out3[16]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_17_ ( .D(DataOutReg3_gff_n245), 
        .CK(clk), .Q(data_out3[17]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_18_ ( .D(DataOutReg3_gff_n244), 
        .CK(clk), .Q(data_out3[18]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_19_ ( .D(DataOutReg3_gff_n243), 
        .CK(clk), .Q(data_out3[19]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_20_ ( .D(DataOutReg3_gff_n242), 
        .CK(clk), .Q(data_out3[20]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_21_ ( .D(DataOutReg3_gff_n241), 
        .CK(clk), .Q(data_out3[21]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_22_ ( .D(DataOutReg3_gff_n240), 
        .CK(clk), .Q(data_out3[22]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_23_ ( .D(DataOutReg3_gff_n239), 
        .CK(clk), .Q(data_out3[23]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_24_ ( .D(DataOutReg3_gff_n238), 
        .CK(clk), .Q(data_out3[24]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_25_ ( .D(DataOutReg3_gff_n237), 
        .CK(clk), .Q(data_out3[25]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_26_ ( .D(DataOutReg3_gff_n236), 
        .CK(clk), .Q(data_out3[26]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_27_ ( .D(DataOutReg3_gff_n235), 
        .CK(clk), .Q(data_out3[27]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_28_ ( .D(DataOutReg3_gff_n234), 
        .CK(clk), .Q(data_out3[28]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_29_ ( .D(DataOutReg3_gff_n233), 
        .CK(clk), .Q(data_out3[29]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_30_ ( .D(DataOutReg3_gff_n232), 
        .CK(clk), .Q(data_out3[30]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_31_ ( .D(DataOutReg3_gff_n231), 
        .CK(clk), .Q(data_out3[31]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_32_ ( .D(DataOutReg3_gff_n230), 
        .CK(clk), .Q(data_out3[32]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_33_ ( .D(DataOutReg3_gff_n229), 
        .CK(clk), .Q(data_out3[33]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_34_ ( .D(DataOutReg3_gff_n228), 
        .CK(clk), .Q(data_out3[34]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_35_ ( .D(DataOutReg3_gff_n227), 
        .CK(clk), .Q(data_out3[35]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_36_ ( .D(DataOutReg3_gff_n226), 
        .CK(clk), .Q(data_out3[36]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_37_ ( .D(DataOutReg3_gff_n225), 
        .CK(clk), .Q(data_out3[37]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_38_ ( .D(DataOutReg3_gff_n224), 
        .CK(clk), .Q(data_out3[38]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_39_ ( .D(DataOutReg3_gff_n223), 
        .CK(clk), .Q(data_out3[39]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_40_ ( .D(DataOutReg3_gff_n222), 
        .CK(clk), .Q(data_out3[40]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_41_ ( .D(DataOutReg3_gff_n221), 
        .CK(clk), .Q(data_out3[41]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_42_ ( .D(DataOutReg3_gff_n220), 
        .CK(clk), .Q(data_out3[42]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_43_ ( .D(DataOutReg3_gff_n219), 
        .CK(clk), .Q(data_out3[43]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_44_ ( .D(DataOutReg3_gff_n218), 
        .CK(clk), .Q(data_out3[44]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_45_ ( .D(DataOutReg3_gff_n217), 
        .CK(clk), .Q(data_out3[45]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_46_ ( .D(DataOutReg3_gff_n216), 
        .CK(clk), .Q(data_out3[46]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_47_ ( .D(DataOutReg3_gff_n215), 
        .CK(clk), .Q(data_out3[47]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_48_ ( .D(DataOutReg3_gff_n214), 
        .CK(clk), .Q(data_out3[48]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_49_ ( .D(DataOutReg3_gff_n213), 
        .CK(clk), .Q(data_out3[49]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_50_ ( .D(DataOutReg3_gff_n212), 
        .CK(clk), .Q(data_out3[50]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_51_ ( .D(DataOutReg3_gff_n211), 
        .CK(clk), .Q(data_out3[51]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_52_ ( .D(DataOutReg3_gff_n210), 
        .CK(clk), .Q(data_out3[52]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_53_ ( .D(DataOutReg3_gff_n209), 
        .CK(clk), .Q(data_out3[53]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_54_ ( .D(DataOutReg3_gff_n208), 
        .CK(clk), .Q(data_out3[54]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_55_ ( .D(DataOutReg3_gff_n207), 
        .CK(clk), .Q(data_out3[55]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_56_ ( .D(DataOutReg3_gff_n206), 
        .CK(clk), .Q(data_out3[56]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_57_ ( .D(DataOutReg3_gff_n205), 
        .CK(clk), .Q(data_out3[57]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_58_ ( .D(DataOutReg3_gff_n204), 
        .CK(clk), .Q(data_out3[58]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_59_ ( .D(DataOutReg3_gff_n203), 
        .CK(clk), .Q(data_out3[59]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_60_ ( .D(DataOutReg3_gff_n202), 
        .CK(clk), .Q(data_out3[60]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_61_ ( .D(DataOutReg3_gff_n201), 
        .CK(clk), .Q(data_out3[61]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_62_ ( .D(DataOutReg3_gff_n200), 
        .CK(clk), .Q(data_out3[62]) , .QN() ); 
  DFF_X1 DataOutReg3_gff_s_current_state_reg_63_ ( .D(DataOutReg3_gff_n199), 
        .CK(clk), .Q(data_out3[63]) , .QN() ); 
endmodule