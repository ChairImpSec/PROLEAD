module circuit ( clk, nReset, r, dataIn1, dataIn2, dataIn3, key1, key2, key3, 
        dataOut1, dataOut2, dataOut3, done );
  input [7:0] r;
  input [3:0] dataIn1;
  input [3:0] dataIn2;
  input [3:0] dataIn3;
  input [3:0] key1;
  input [3:0] key2;
  input [3:0] key3;
  output [3:0] dataOut1;
  output [3:0] dataOut2;
  output [3:0] dataOut3;
  input clk, nReset;
  output done;
  wire   selInit, selP, selSbox, enKey, enData, n4, fsm_n31, fsm_n30, fsm_n29,
         fsm_n28, fsm_n27, fsm_n26, fsm_n25, fsm_n24, fsm_n20, fsm_n19,
         fsm_n18, fsm_n17, fsm_n16, fsm_n15, fsm_n14, fsm_n13, fsm_n12,
         fsm_n11, fsm_n10, fsm_n9, fsm_n23, fsm_n22, fsm_n21, fsm_ps_state_0_,
         fsm_ps_state_1_, fsm_ps_state_2_, fsm_countSerial_0_,
         fsm_countSerial_1_, fsm_countSerial_2_, fsm_countSerial_3_,
         fsm_countSerial_4_, fsm_en_countSerial, fsm_rst_countSerial,
         fsm_en_countRound, fsm_cnt_rnd_n38, fsm_cnt_rnd_n37, fsm_cnt_rnd_n36,
         fsm_cnt_rnd_n35, fsm_cnt_rnd_n34, fsm_cnt_rnd_n33, fsm_cnt_rnd_n32,
         fsm_cnt_rnd_n31, fsm_cnt_rnd_n30, fsm_cnt_rnd_n29, fsm_cnt_rnd_n28,
         fsm_cnt_rnd_n27, fsm_cnt_rnd_n26, fsm_cnt_rnd_n25, fsm_cnt_rnd_n24,
         fsm_cnt_rnd_n23, fsm_cnt_rnd_n20, fsm_cnt_rnd_n22, fsm_cnt_rnd_n21,
         fsm_cnt_rnd_n19, fsm_cnt_rnd_n2, fsm_cnt_ser_n43, fsm_cnt_ser_n42,
         fsm_cnt_ser_n41, fsm_cnt_ser_n40, fsm_cnt_ser_n39, fsm_cnt_ser_n38,
         fsm_cnt_ser_n37, fsm_cnt_ser_n36, fsm_cnt_ser_n35, fsm_cnt_ser_n34,
         fsm_cnt_ser_n33, fsm_cnt_ser_n32, fsm_cnt_ser_n31, fsm_cnt_ser_n30,
         fsm_cnt_ser_n29, fsm_cnt_ser_n28, fsm_cnt_ser_n26, fsm_cnt_ser_n25,
         fsm_cnt_ser_n23, fsm_cnt_ser_n22, fsm_cnt_ser_n20, fsm_cnt_ser_n5,
         state1FF_n4, state1FF_n3, state1FF_n2, state1FF_n1,
         state1FF_state_n13, state1FF_state_n12, state1FF_state_n11,
         state1FF_state_n10, state1FF_state_n9, state1FF_state_n8,
         state1FF_state_n7, state1FF_state_n6, state1FF_state_gff_1_SFF_0_n10,
         state1FF_state_gff_1_SFF_0_n9, state1FF_state_gff_1_SFF_0_n7,
         state1FF_state_gff_1_SFF_0_n6, state1FF_state_gff_1_SFF_1_n11,
         state1FF_state_gff_1_SFF_1_n10, state1FF_state_gff_1_SFF_1_n8,
         state1FF_state_gff_1_SFF_1_n7, state1FF_state_gff_1_SFF_2_n12,
         state1FF_state_gff_1_SFF_2_n11, state1FF_state_gff_1_SFF_2_n10,
         state1FF_state_gff_1_SFF_2_n8, state1FF_state_gff_1_SFF_2_n7,
         state1FF_state_gff_1_SFF_3_n12, state1FF_state_gff_1_SFF_3_n11,
         state1FF_state_gff_1_SFF_3_n10, state1FF_state_gff_1_SFF_3_n8,
         state1FF_state_gff_1_SFF_3_n7, state1FF_state_gff_2_SFF_0_n12,
         state1FF_state_gff_2_SFF_0_n11, state1FF_state_gff_2_SFF_0_n10,
         state1FF_state_gff_2_SFF_0_n8, state1FF_state_gff_2_SFF_0_n7,
         state1FF_state_gff_2_SFF_1_n12, state1FF_state_gff_2_SFF_1_n11,
         state1FF_state_gff_2_SFF_1_n10, state1FF_state_gff_2_SFF_1_n8,
         state1FF_state_gff_2_SFF_1_n7, state1FF_state_gff_2_SFF_2_n11,
         state1FF_state_gff_2_SFF_2_n10, state1FF_state_gff_2_SFF_2_n8,
         state1FF_state_gff_2_SFF_2_n7, state1FF_state_gff_2_SFF_3_n11,
         state1FF_state_gff_2_SFF_3_n10, state1FF_state_gff_2_SFF_3_n8,
         state1FF_state_gff_2_SFF_3_n7, state1FF_state_gff_3_SFF_0_n12,
         state1FF_state_gff_3_SFF_0_n11, state1FF_state_gff_3_SFF_0_n10,
         state1FF_state_gff_3_SFF_0_n8, state1FF_state_gff_3_SFF_0_n7,
         state1FF_state_gff_3_SFF_1_n12, state1FF_state_gff_3_SFF_1_n11,
         state1FF_state_gff_3_SFF_1_n10, state1FF_state_gff_3_SFF_1_n8,
         state1FF_state_gff_3_SFF_1_n7, state1FF_state_gff_3_SFF_2_n12,
         state1FF_state_gff_3_SFF_2_n11, state1FF_state_gff_3_SFF_2_n10,
         state1FF_state_gff_3_SFF_2_n8, state1FF_state_gff_3_SFF_2_n7,
         state1FF_state_gff_3_SFF_3_n12, state1FF_state_gff_3_SFF_3_n11,
         state1FF_state_gff_3_SFF_3_n10, state1FF_state_gff_3_SFF_3_n8,
         state1FF_state_gff_3_SFF_3_n7, state1FF_state_gff_4_SFF_0_n11,
         state1FF_state_gff_4_SFF_0_n10, state1FF_state_gff_4_SFF_0_n8,
         state1FF_state_gff_4_SFF_0_n7, state1FF_state_gff_4_SFF_1_n11,
         state1FF_state_gff_4_SFF_1_n10, state1FF_state_gff_4_SFF_1_n8,
         state1FF_state_gff_4_SFF_1_n7, state1FF_state_gff_4_SFF_2_n11,
         state1FF_state_gff_4_SFF_2_n10, state1FF_state_gff_4_SFF_2_n9,
         state1FF_state_gff_4_SFF_2_n7, state1FF_state_gff_4_SFF_2_n6,
         state1FF_state_gff_4_SFF_3_n11, state1FF_state_gff_4_SFF_3_n10,
         state1FF_state_gff_4_SFF_3_n9, state1FF_state_gff_4_SFF_3_n7,
         state1FF_state_gff_4_SFF_3_n6, state1FF_state_gff_5_SFF_0_n11,
         state1FF_state_gff_5_SFF_0_n10, state1FF_state_gff_5_SFF_0_n9,
         state1FF_state_gff_5_SFF_0_n7, state1FF_state_gff_5_SFF_0_n6,
         state1FF_state_gff_5_SFF_1_n11, state1FF_state_gff_5_SFF_1_n10,
         state1FF_state_gff_5_SFF_1_n9, state1FF_state_gff_5_SFF_1_n7,
         state1FF_state_gff_5_SFF_1_n6, state1FF_state_gff_5_SFF_2_n11,
         state1FF_state_gff_5_SFF_2_n10, state1FF_state_gff_5_SFF_2_n9,
         state1FF_state_gff_5_SFF_2_n7, state1FF_state_gff_5_SFF_2_n6,
         state1FF_state_gff_5_SFF_3_n11, state1FF_state_gff_5_SFF_3_n10,
         state1FF_state_gff_5_SFF_3_n9, state1FF_state_gff_5_SFF_3_n7,
         state1FF_state_gff_5_SFF_3_n6, state1FF_state_gff_6_SFF_0_n12,
         state1FF_state_gff_6_SFF_0_n11, state1FF_state_gff_6_SFF_0_n10,
         state1FF_state_gff_6_SFF_0_n8, state1FF_state_gff_6_SFF_0_n7,
         state1FF_state_gff_6_SFF_1_n12, state1FF_state_gff_6_SFF_1_n11,
         state1FF_state_gff_6_SFF_1_n10, state1FF_state_gff_6_SFF_1_n8,
         state1FF_state_gff_6_SFF_1_n7, state1FF_state_gff_6_SFF_2_n12,
         state1FF_state_gff_6_SFF_2_n11, state1FF_state_gff_6_SFF_2_n10,
         state1FF_state_gff_6_SFF_2_n8, state1FF_state_gff_6_SFF_2_n7,
         state1FF_state_gff_6_SFF_3_n12, state1FF_state_gff_6_SFF_3_n11,
         state1FF_state_gff_6_SFF_3_n10, state1FF_state_gff_6_SFF_3_n8,
         state1FF_state_gff_6_SFF_3_n7, state1FF_state_gff_7_SFF_0_n12,
         state1FF_state_gff_7_SFF_0_n11, state1FF_state_gff_7_SFF_0_n10,
         state1FF_state_gff_7_SFF_0_n8, state1FF_state_gff_7_SFF_0_n7,
         state1FF_state_gff_7_SFF_1_n12, state1FF_state_gff_7_SFF_1_n11,
         state1FF_state_gff_7_SFF_1_n10, state1FF_state_gff_7_SFF_1_n8,
         state1FF_state_gff_7_SFF_1_n7, state1FF_state_gff_7_SFF_2_n11,
         state1FF_state_gff_7_SFF_2_n10, state1FF_state_gff_7_SFF_2_n8,
         state1FF_state_gff_7_SFF_2_n7, state1FF_state_gff_7_SFF_3_n11,
         state1FF_state_gff_7_SFF_3_n10, state1FF_state_gff_7_SFF_3_n8,
         state1FF_state_gff_7_SFF_3_n7, state1FF_state_gff_8_SFF_0_n12,
         state1FF_state_gff_8_SFF_0_n11, state1FF_state_gff_8_SFF_0_n10,
         state1FF_state_gff_8_SFF_0_n8, state1FF_state_gff_8_SFF_0_n7,
         state1FF_state_gff_8_SFF_1_n12, state1FF_state_gff_8_SFF_1_n11,
         state1FF_state_gff_8_SFF_1_n10, state1FF_state_gff_8_SFF_1_n8,
         state1FF_state_gff_8_SFF_1_n7, state1FF_state_gff_8_SFF_2_n11,
         state1FF_state_gff_8_SFF_2_n10, state1FF_state_gff_8_SFF_2_n9,
         state1FF_state_gff_8_SFF_2_n7, state1FF_state_gff_8_SFF_2_n6,
         state1FF_state_gff_8_SFF_3_n11, state1FF_state_gff_8_SFF_3_n10,
         state1FF_state_gff_8_SFF_3_n9, state1FF_state_gff_8_SFF_3_n7,
         state1FF_state_gff_8_SFF_3_n6, state1FF_state_gff_9_SFF_0_n11,
         state1FF_state_gff_9_SFF_0_n10, state1FF_state_gff_9_SFF_0_n9,
         state1FF_state_gff_9_SFF_0_n7, state1FF_state_gff_9_SFF_0_n6,
         state1FF_state_gff_9_SFF_1_n11, state1FF_state_gff_9_SFF_1_n10,
         state1FF_state_gff_9_SFF_1_n9, state1FF_state_gff_9_SFF_1_n7,
         state1FF_state_gff_9_SFF_1_n6, state1FF_state_gff_9_SFF_2_n11,
         state1FF_state_gff_9_SFF_2_n10, state1FF_state_gff_9_SFF_2_n9,
         state1FF_state_gff_9_SFF_2_n7, state1FF_state_gff_9_SFF_2_n6,
         state1FF_state_gff_9_SFF_3_n11, state1FF_state_gff_9_SFF_3_n10,
         state1FF_state_gff_9_SFF_3_n9, state1FF_state_gff_9_SFF_3_n7,
         state1FF_state_gff_9_SFF_3_n6, state1FF_state_gff_10_SFF_0_n11,
         state1FF_state_gff_10_SFF_0_n10, state1FF_state_gff_10_SFF_0_n8,
         state1FF_state_gff_10_SFF_0_n7, state1FF_state_gff_10_SFF_1_n11,
         state1FF_state_gff_10_SFF_1_n10, state1FF_state_gff_10_SFF_1_n8,
         state1FF_state_gff_10_SFF_1_n7, state1FF_state_gff_10_SFF_2_n11,
         state1FF_state_gff_10_SFF_2_n10, state1FF_state_gff_10_SFF_2_n8,
         state1FF_state_gff_10_SFF_2_n7, state1FF_state_gff_10_SFF_3_n11,
         state1FF_state_gff_10_SFF_3_n10, state1FF_state_gff_10_SFF_3_n8,
         state1FF_state_gff_10_SFF_3_n7, state1FF_state_gff_11_SFF_0_n12,
         state1FF_state_gff_11_SFF_0_n11, state1FF_state_gff_11_SFF_0_n10,
         state1FF_state_gff_11_SFF_0_n8, state1FF_state_gff_11_SFF_0_n7,
         state1FF_state_gff_11_SFF_1_n12, state1FF_state_gff_11_SFF_1_n11,
         state1FF_state_gff_11_SFF_1_n10, state1FF_state_gff_11_SFF_1_n8,
         state1FF_state_gff_11_SFF_1_n7, state1FF_state_gff_11_SFF_2_n12,
         state1FF_state_gff_11_SFF_2_n11, state1FF_state_gff_11_SFF_2_n10,
         state1FF_state_gff_11_SFF_2_n8, state1FF_state_gff_11_SFF_2_n7,
         state1FF_state_gff_11_SFF_3_n12, state1FF_state_gff_11_SFF_3_n11,
         state1FF_state_gff_11_SFF_3_n10, state1FF_state_gff_11_SFF_3_n8,
         state1FF_state_gff_11_SFF_3_n7, state1FF_state_gff_12_SFF_0_n11,
         state1FF_state_gff_12_SFF_0_n10, state1FF_state_gff_12_SFF_0_n8,
         state1FF_state_gff_12_SFF_0_n7, state1FF_state_gff_12_SFF_1_n11,
         state1FF_state_gff_12_SFF_1_n10, state1FF_state_gff_12_SFF_1_n8,
         state1FF_state_gff_12_SFF_1_n7, state1FF_state_gff_12_SFF_2_n11,
         state1FF_state_gff_12_SFF_2_n10, state1FF_state_gff_12_SFF_2_n9,
         state1FF_state_gff_12_SFF_2_n7, state1FF_state_gff_12_SFF_2_n6,
         state1FF_state_gff_12_SFF_3_n11, state1FF_state_gff_12_SFF_3_n10,
         state1FF_state_gff_12_SFF_3_n9, state1FF_state_gff_12_SFF_3_n7,
         state1FF_state_gff_12_SFF_3_n6, state1FF_state_gff_13_SFF_0_n11,
         state1FF_state_gff_13_SFF_0_n10, state1FF_state_gff_13_SFF_0_n9,
         state1FF_state_gff_13_SFF_0_n7, state1FF_state_gff_13_SFF_0_n6,
         state1FF_state_gff_13_SFF_1_n11, state1FF_state_gff_13_SFF_1_n10,
         state1FF_state_gff_13_SFF_1_n9, state1FF_state_gff_13_SFF_1_n7,
         state1FF_state_gff_13_SFF_1_n6, state1FF_state_gff_13_SFF_2_n11,
         state1FF_state_gff_13_SFF_2_n10, state1FF_state_gff_13_SFF_2_n9,
         state1FF_state_gff_13_SFF_2_n7, state1FF_state_gff_13_SFF_2_n6,
         state1FF_state_gff_13_SFF_3_n11, state1FF_state_gff_13_SFF_3_n10,
         state1FF_state_gff_13_SFF_3_n9, state1FF_state_gff_13_SFF_3_n7,
         state1FF_state_gff_13_SFF_3_n6, state1FF_state_gff_14_SFF_0_n11,
         state1FF_state_gff_14_SFF_0_n10, state1FF_state_gff_14_SFF_0_n8,
         state1FF_state_gff_14_SFF_0_n7, state1FF_state_gff_14_SFF_1_n11,
         state1FF_state_gff_14_SFF_1_n10, state1FF_state_gff_14_SFF_1_n8,
         state1FF_state_gff_14_SFF_1_n7, state1FF_state_gff_14_SFF_2_n11,
         state1FF_state_gff_14_SFF_2_n10, state1FF_state_gff_14_SFF_2_n8,
         state1FF_state_gff_14_SFF_2_n7, state1FF_state_gff_14_SFF_3_n11,
         state1FF_state_gff_14_SFF_3_n10, state1FF_state_gff_14_SFF_3_n8,
         state1FF_state_gff_14_SFF_3_n7, state1FF_state_gff_15_SFF_0_n11,
         state1FF_state_gff_15_SFF_0_n10, state1FF_state_gff_15_SFF_0_n8,
         state1FF_state_gff_15_SFF_0_n7, state1FF_state_gff_15_SFF_1_n11,
         state1FF_state_gff_15_SFF_1_n10, state1FF_state_gff_15_SFF_1_n8,
         state1FF_state_gff_15_SFF_1_n7, state1FF_state_gff_15_SFF_2_n11,
         state1FF_state_gff_15_SFF_2_n10, state1FF_state_gff_15_SFF_2_n8,
         state1FF_state_gff_15_SFF_2_n7, state1FF_state_gff_15_SFF_3_n11,
         state1FF_state_gff_15_SFF_3_n10, state1FF_state_gff_15_SFF_3_n9,
         state1FF_state_gff_15_SFF_3_n7, state1FF_state_gff_15_SFF_3_n6,
         state1FF_state_gff_16_SFF_0_n11, state1FF_state_gff_16_SFF_0_n10,
         state1FF_state_gff_16_SFF_0_n9, state1FF_state_gff_16_SFF_0_n7,
         state1FF_state_gff_16_SFF_0_n6, state1FF_state_gff_16_SFF_1_n10,
         state1FF_state_gff_16_SFF_1_n9, state1FF_state_gff_16_SFF_1_n7,
         state1FF_state_gff_16_SFF_1_n6, state1FF_state_gff_16_SFF_2_n10,
         state1FF_state_gff_16_SFF_2_n9, state1FF_state_gff_16_SFF_2_n7,
         state1FF_state_gff_16_SFF_2_n6, state1FF_state_gff_16_SFF_3_n10,
         state1FF_state_gff_16_SFF_3_n9, state1FF_state_gff_16_SFF_3_n7,
         state1FF_state_gff_16_SFF_3_n6, state2FF_n4, state2FF_n3, state2FF_n2,
         state2FF_n1, state2FF_state_n13, state2FF_state_n12,
         state2FF_state_n11, state2FF_state_n10, state2FF_state_n9,
         state2FF_state_n8, state2FF_state_n7, state2FF_state_n6,
         state2FF_state_gff_1_SFF_0_n12, state2FF_state_gff_1_SFF_0_n11,
         state2FF_state_gff_1_SFF_0_n10, state2FF_state_gff_1_SFF_0_n8,
         state2FF_state_gff_1_SFF_0_n7, state2FF_state_gff_1_SFF_1_n12,
         state2FF_state_gff_1_SFF_1_n11, state2FF_state_gff_1_SFF_1_n10,
         state2FF_state_gff_1_SFF_1_n8, state2FF_state_gff_1_SFF_1_n7,
         state2FF_state_gff_1_SFF_2_n12, state2FF_state_gff_1_SFF_2_n11,
         state2FF_state_gff_1_SFF_2_n10, state2FF_state_gff_1_SFF_2_n8,
         state2FF_state_gff_1_SFF_2_n7, state2FF_state_gff_1_SFF_3_n12,
         state2FF_state_gff_1_SFF_3_n11, state2FF_state_gff_1_SFF_3_n10,
         state2FF_state_gff_1_SFF_3_n8, state2FF_state_gff_1_SFF_3_n7,
         state2FF_state_gff_2_SFF_0_n12, state2FF_state_gff_2_SFF_0_n11,
         state2FF_state_gff_2_SFF_0_n10, state2FF_state_gff_2_SFF_0_n8,
         state2FF_state_gff_2_SFF_0_n7, state2FF_state_gff_2_SFF_1_n12,
         state2FF_state_gff_2_SFF_1_n11, state2FF_state_gff_2_SFF_1_n10,
         state2FF_state_gff_2_SFF_1_n8, state2FF_state_gff_2_SFF_1_n7,
         state2FF_state_gff_2_SFF_2_n12, state2FF_state_gff_2_SFF_2_n11,
         state2FF_state_gff_2_SFF_2_n10, state2FF_state_gff_2_SFF_2_n8,
         state2FF_state_gff_2_SFF_2_n7, state2FF_state_gff_2_SFF_3_n12,
         state2FF_state_gff_2_SFF_3_n11, state2FF_state_gff_2_SFF_3_n10,
         state2FF_state_gff_2_SFF_3_n8, state2FF_state_gff_2_SFF_3_n7,
         state2FF_state_gff_3_SFF_0_n12, state2FF_state_gff_3_SFF_0_n11,
         state2FF_state_gff_3_SFF_0_n10, state2FF_state_gff_3_SFF_0_n8,
         state2FF_state_gff_3_SFF_0_n7, state2FF_state_gff_3_SFF_1_n12,
         state2FF_state_gff_3_SFF_1_n11, state2FF_state_gff_3_SFF_1_n10,
         state2FF_state_gff_3_SFF_1_n8, state2FF_state_gff_3_SFF_1_n7,
         state2FF_state_gff_3_SFF_2_n11, state2FF_state_gff_3_SFF_2_n10,
         state2FF_state_gff_3_SFF_2_n9, state2FF_state_gff_3_SFF_2_n7,
         state2FF_state_gff_3_SFF_2_n6, state2FF_state_gff_3_SFF_3_n11,
         state2FF_state_gff_3_SFF_3_n10, state2FF_state_gff_3_SFF_3_n9,
         state2FF_state_gff_3_SFF_3_n7, state2FF_state_gff_3_SFF_3_n6,
         state2FF_state_gff_4_SFF_0_n11, state2FF_state_gff_4_SFF_0_n10,
         state2FF_state_gff_4_SFF_0_n9, state2FF_state_gff_4_SFF_0_n7,
         state2FF_state_gff_4_SFF_0_n6, state2FF_state_gff_4_SFF_1_n11,
         state2FF_state_gff_4_SFF_1_n10, state2FF_state_gff_4_SFF_1_n9,
         state2FF_state_gff_4_SFF_1_n7, state2FF_state_gff_4_SFF_1_n6,
         state2FF_state_gff_4_SFF_2_n11, state2FF_state_gff_4_SFF_2_n10,
         state2FF_state_gff_4_SFF_2_n9, state2FF_state_gff_4_SFF_2_n7,
         state2FF_state_gff_4_SFF_2_n6, state2FF_state_gff_4_SFF_3_n11,
         state2FF_state_gff_4_SFF_3_n10, state2FF_state_gff_4_SFF_3_n9,
         state2FF_state_gff_4_SFF_3_n7, state2FF_state_gff_4_SFF_3_n6,
         state2FF_state_gff_5_SFF_0_n12, state2FF_state_gff_5_SFF_0_n11,
         state2FF_state_gff_5_SFF_0_n10, state2FF_state_gff_5_SFF_0_n8,
         state2FF_state_gff_5_SFF_0_n7, state2FF_state_gff_5_SFF_1_n12,
         state2FF_state_gff_5_SFF_1_n11, state2FF_state_gff_5_SFF_1_n10,
         state2FF_state_gff_5_SFF_1_n8, state2FF_state_gff_5_SFF_1_n7,
         state2FF_state_gff_5_SFF_2_n11, state2FF_state_gff_5_SFF_2_n10,
         state2FF_state_gff_5_SFF_2_n8, state2FF_state_gff_5_SFF_2_n7,
         state2FF_state_gff_5_SFF_3_n11, state2FF_state_gff_5_SFF_3_n10,
         state2FF_state_gff_5_SFF_3_n8, state2FF_state_gff_5_SFF_3_n7,
         state2FF_state_gff_6_SFF_0_n11, state2FF_state_gff_6_SFF_0_n10,
         state2FF_state_gff_6_SFF_0_n8, state2FF_state_gff_6_SFF_0_n7,
         state2FF_state_gff_6_SFF_1_n11, state2FF_state_gff_6_SFF_1_n10,
         state2FF_state_gff_6_SFF_1_n8, state2FF_state_gff_6_SFF_1_n7,
         state2FF_state_gff_6_SFF_2_n11, state2FF_state_gff_6_SFF_2_n10,
         state2FF_state_gff_6_SFF_2_n8, state2FF_state_gff_6_SFF_2_n7,
         state2FF_state_gff_6_SFF_3_n11, state2FF_state_gff_6_SFF_3_n10,
         state2FF_state_gff_6_SFF_3_n8, state2FF_state_gff_6_SFF_3_n7,
         state2FF_state_gff_7_SFF_0_n11, state2FF_state_gff_7_SFF_0_n10,
         state2FF_state_gff_7_SFF_0_n8, state2FF_state_gff_7_SFF_0_n7,
         state2FF_state_gff_7_SFF_1_n11, state2FF_state_gff_7_SFF_1_n10,
         state2FF_state_gff_7_SFF_1_n8, state2FF_state_gff_7_SFF_1_n7,
         state2FF_state_gff_7_SFF_2_n11, state2FF_state_gff_7_SFF_2_n10,
         state2FF_state_gff_7_SFF_2_n9, state2FF_state_gff_7_SFF_2_n7,
         state2FF_state_gff_7_SFF_2_n6, state2FF_state_gff_7_SFF_3_n11,
         state2FF_state_gff_7_SFF_3_n10, state2FF_state_gff_7_SFF_3_n9,
         state2FF_state_gff_7_SFF_3_n7, state2FF_state_gff_7_SFF_3_n6,
         state2FF_state_gff_8_SFF_0_n11, state2FF_state_gff_8_SFF_0_n10,
         state2FF_state_gff_8_SFF_0_n9, state2FF_state_gff_8_SFF_0_n7,
         state2FF_state_gff_8_SFF_0_n6, state2FF_state_gff_8_SFF_1_n11,
         state2FF_state_gff_8_SFF_1_n10, state2FF_state_gff_8_SFF_1_n9,
         state2FF_state_gff_8_SFF_1_n7, state2FF_state_gff_8_SFF_1_n6,
         state2FF_state_gff_8_SFF_2_n11, state2FF_state_gff_8_SFF_2_n10,
         state2FF_state_gff_8_SFF_2_n9, state2FF_state_gff_8_SFF_2_n7,
         state2FF_state_gff_8_SFF_2_n6, state2FF_state_gff_8_SFF_3_n11,
         state2FF_state_gff_8_SFF_3_n10, state2FF_state_gff_8_SFF_3_n9,
         state2FF_state_gff_8_SFF_3_n7, state2FF_state_gff_8_SFF_3_n6,
         state2FF_state_gff_9_SFF_0_n12, state2FF_state_gff_9_SFF_0_n11,
         state2FF_state_gff_9_SFF_0_n10, state2FF_state_gff_9_SFF_0_n8,
         state2FF_state_gff_9_SFF_0_n7, state2FF_state_gff_9_SFF_1_n12,
         state2FF_state_gff_9_SFF_1_n11, state2FF_state_gff_9_SFF_1_n10,
         state2FF_state_gff_9_SFF_1_n8, state2FF_state_gff_9_SFF_1_n7,
         state2FF_state_gff_9_SFF_2_n12, state2FF_state_gff_9_SFF_2_n11,
         state2FF_state_gff_9_SFF_2_n10, state2FF_state_gff_9_SFF_2_n8,
         state2FF_state_gff_9_SFF_2_n7, state2FF_state_gff_9_SFF_3_n12,
         state2FF_state_gff_9_SFF_3_n11, state2FF_state_gff_9_SFF_3_n10,
         state2FF_state_gff_9_SFF_3_n8, state2FF_state_gff_9_SFF_3_n7,
         state2FF_state_gff_10_SFF_0_n12, state2FF_state_gff_10_SFF_0_n11,
         state2FF_state_gff_10_SFF_0_n10, state2FF_state_gff_10_SFF_0_n8,
         state2FF_state_gff_10_SFF_0_n7, state2FF_state_gff_10_SFF_1_n12,
         state2FF_state_gff_10_SFF_1_n11, state2FF_state_gff_10_SFF_1_n10,
         state2FF_state_gff_10_SFF_1_n8, state2FF_state_gff_10_SFF_1_n7,
         state2FF_state_gff_10_SFF_2_n12, state2FF_state_gff_10_SFF_2_n11,
         state2FF_state_gff_10_SFF_2_n10, state2FF_state_gff_10_SFF_2_n8,
         state2FF_state_gff_10_SFF_2_n7, state2FF_state_gff_10_SFF_3_n12,
         state2FF_state_gff_10_SFF_3_n11, state2FF_state_gff_10_SFF_3_n10,
         state2FF_state_gff_10_SFF_3_n8, state2FF_state_gff_10_SFF_3_n7,
         state2FF_state_gff_11_SFF_0_n11, state2FF_state_gff_11_SFF_0_n10,
         state2FF_state_gff_11_SFF_0_n8, state2FF_state_gff_11_SFF_0_n7,
         state2FF_state_gff_11_SFF_1_n11, state2FF_state_gff_11_SFF_1_n10,
         state2FF_state_gff_11_SFF_1_n8, state2FF_state_gff_11_SFF_1_n7,
         state2FF_state_gff_11_SFF_2_n11, state2FF_state_gff_11_SFF_2_n10,
         state2FF_state_gff_11_SFF_2_n9, state2FF_state_gff_11_SFF_2_n7,
         state2FF_state_gff_11_SFF_2_n6, state2FF_state_gff_11_SFF_3_n11,
         state2FF_state_gff_11_SFF_3_n10, state2FF_state_gff_11_SFF_3_n9,
         state2FF_state_gff_11_SFF_3_n7, state2FF_state_gff_11_SFF_3_n6,
         state2FF_state_gff_12_SFF_0_n11, state2FF_state_gff_12_SFF_0_n10,
         state2FF_state_gff_12_SFF_0_n9, state2FF_state_gff_12_SFF_0_n7,
         state2FF_state_gff_12_SFF_0_n6, state2FF_state_gff_12_SFF_1_n11,
         state2FF_state_gff_12_SFF_1_n10, state2FF_state_gff_12_SFF_1_n9,
         state2FF_state_gff_12_SFF_1_n7, state2FF_state_gff_12_SFF_1_n6,
         state2FF_state_gff_12_SFF_2_n10, state2FF_state_gff_12_SFF_2_n9,
         state2FF_state_gff_12_SFF_2_n7, state2FF_state_gff_12_SFF_2_n6,
         state2FF_state_gff_12_SFF_3_n10, state2FF_state_gff_12_SFF_3_n9,
         state2FF_state_gff_12_SFF_3_n7, state2FF_state_gff_12_SFF_3_n6,
         state2FF_state_gff_13_SFF_0_n12, state2FF_state_gff_13_SFF_0_n11,
         state2FF_state_gff_13_SFF_0_n10, state2FF_state_gff_13_SFF_0_n8,
         state2FF_state_gff_13_SFF_0_n7, state2FF_state_gff_13_SFF_1_n12,
         state2FF_state_gff_13_SFF_1_n11, state2FF_state_gff_13_SFF_1_n10,
         state2FF_state_gff_13_SFF_1_n8, state2FF_state_gff_13_SFF_1_n7,
         state2FF_state_gff_13_SFF_2_n11, state2FF_state_gff_13_SFF_2_n10,
         state2FF_state_gff_13_SFF_2_n8, state2FF_state_gff_13_SFF_2_n7,
         state2FF_state_gff_13_SFF_3_n11, state2FF_state_gff_13_SFF_3_n10,
         state2FF_state_gff_13_SFF_3_n8, state2FF_state_gff_13_SFF_3_n7,
         state2FF_state_gff_14_SFF_0_n11, state2FF_state_gff_14_SFF_0_n10,
         state2FF_state_gff_14_SFF_0_n8, state2FF_state_gff_14_SFF_0_n7,
         state2FF_state_gff_14_SFF_1_n11, state2FF_state_gff_14_SFF_1_n10,
         state2FF_state_gff_14_SFF_1_n8, state2FF_state_gff_14_SFF_1_n7,
         state2FF_state_gff_14_SFF_2_n11, state2FF_state_gff_14_SFF_2_n10,
         state2FF_state_gff_14_SFF_2_n8, state2FF_state_gff_14_SFF_2_n7,
         state2FF_state_gff_14_SFF_3_n11, state2FF_state_gff_14_SFF_3_n10,
         state2FF_state_gff_14_SFF_3_n8, state2FF_state_gff_14_SFF_3_n7,
         state2FF_state_gff_15_SFF_0_n11, state2FF_state_gff_15_SFF_0_n10,
         state2FF_state_gff_15_SFF_0_n8, state2FF_state_gff_15_SFF_0_n7,
         state2FF_state_gff_15_SFF_1_n11, state2FF_state_gff_15_SFF_1_n10,
         state2FF_state_gff_15_SFF_1_n8, state2FF_state_gff_15_SFF_1_n7,
         state2FF_state_gff_15_SFF_2_n11, state2FF_state_gff_15_SFF_2_n10,
         state2FF_state_gff_15_SFF_2_n9, state2FF_state_gff_15_SFF_2_n7,
         state2FF_state_gff_15_SFF_2_n6, state2FF_state_gff_15_SFF_3_n11,
         state2FF_state_gff_15_SFF_3_n10, state2FF_state_gff_15_SFF_3_n9,
         state2FF_state_gff_15_SFF_3_n7, state2FF_state_gff_15_SFF_3_n6,
         state2FF_state_gff_16_SFF_0_n10, state2FF_state_gff_16_SFF_0_n9,
         state2FF_state_gff_16_SFF_0_n7, state2FF_state_gff_16_SFF_0_n6,
         state2FF_state_gff_16_SFF_1_n10, state2FF_state_gff_16_SFF_1_n9,
         state2FF_state_gff_16_SFF_1_n7, state2FF_state_gff_16_SFF_1_n6,
         state2FF_state_gff_16_SFF_2_n10, state2FF_state_gff_16_SFF_2_n9,
         state2FF_state_gff_16_SFF_2_n7, state2FF_state_gff_16_SFF_2_n6,
         state2FF_state_gff_16_SFF_3_n10, state2FF_state_gff_16_SFF_3_n9,
         state2FF_state_gff_16_SFF_3_n7, state2FF_state_gff_16_SFF_3_n6,
         state3FF_n4, state3FF_n3, state3FF_n2, state3FF_n1,
         state3FF_state_n12, state3FF_state_n11, state3FF_state_n10,
         state3FF_state_n9, state3FF_state_n8, state3FF_state_n7,
         state3FF_state_n6, state3FF_state_gff_1_SFF_0_n12,
         state3FF_state_gff_1_SFF_0_n11, state3FF_state_gff_1_SFF_0_n10,
         state3FF_state_gff_1_SFF_0_n8, state3FF_state_gff_1_SFF_0_n7,
         state3FF_state_gff_1_SFF_1_n12, state3FF_state_gff_1_SFF_1_n11,
         state3FF_state_gff_1_SFF_1_n10, state3FF_state_gff_1_SFF_1_n8,
         state3FF_state_gff_1_SFF_1_n7, state3FF_state_gff_1_SFF_2_n12,
         state3FF_state_gff_1_SFF_2_n11, state3FF_state_gff_1_SFF_2_n10,
         state3FF_state_gff_1_SFF_2_n8, state3FF_state_gff_1_SFF_2_n7,
         state3FF_state_gff_1_SFF_3_n12, state3FF_state_gff_1_SFF_3_n11,
         state3FF_state_gff_1_SFF_3_n10, state3FF_state_gff_1_SFF_3_n8,
         state3FF_state_gff_1_SFF_3_n7, state3FF_state_gff_2_SFF_0_n12,
         state3FF_state_gff_2_SFF_0_n11, state3FF_state_gff_2_SFF_0_n10,
         state3FF_state_gff_2_SFF_0_n8, state3FF_state_gff_2_SFF_0_n7,
         state3FF_state_gff_2_SFF_1_n12, state3FF_state_gff_2_SFF_1_n11,
         state3FF_state_gff_2_SFF_1_n10, state3FF_state_gff_2_SFF_1_n8,
         state3FF_state_gff_2_SFF_1_n7, state3FF_state_gff_2_SFF_2_n12,
         state3FF_state_gff_2_SFF_2_n11, state3FF_state_gff_2_SFF_2_n10,
         state3FF_state_gff_2_SFF_2_n8, state3FF_state_gff_2_SFF_2_n7,
         state3FF_state_gff_2_SFF_3_n12, state3FF_state_gff_2_SFF_3_n11,
         state3FF_state_gff_2_SFF_3_n10, state3FF_state_gff_2_SFF_3_n8,
         state3FF_state_gff_2_SFF_3_n7, state3FF_state_gff_3_SFF_0_n12,
         state3FF_state_gff_3_SFF_0_n11, state3FF_state_gff_3_SFF_0_n10,
         state3FF_state_gff_3_SFF_0_n8, state3FF_state_gff_3_SFF_0_n7,
         state3FF_state_gff_3_SFF_1_n12, state3FF_state_gff_3_SFF_1_n11,
         state3FF_state_gff_3_SFF_1_n10, state3FF_state_gff_3_SFF_1_n8,
         state3FF_state_gff_3_SFF_1_n7, state3FF_state_gff_3_SFF_2_n11,
         state3FF_state_gff_3_SFF_2_n10, state3FF_state_gff_3_SFF_2_n9,
         state3FF_state_gff_3_SFF_2_n7, state3FF_state_gff_3_SFF_2_n6,
         state3FF_state_gff_3_SFF_3_n11, state3FF_state_gff_3_SFF_3_n10,
         state3FF_state_gff_3_SFF_3_n9, state3FF_state_gff_3_SFF_3_n7,
         state3FF_state_gff_3_SFF_3_n6, state3FF_state_gff_4_SFF_0_n11,
         state3FF_state_gff_4_SFF_0_n10, state3FF_state_gff_4_SFF_0_n9,
         state3FF_state_gff_4_SFF_0_n7, state3FF_state_gff_4_SFF_0_n6,
         state3FF_state_gff_4_SFF_1_n11, state3FF_state_gff_4_SFF_1_n10,
         state3FF_state_gff_4_SFF_1_n9, state3FF_state_gff_4_SFF_1_n7,
         state3FF_state_gff_4_SFF_1_n6, state3FF_state_gff_4_SFF_2_n11,
         state3FF_state_gff_4_SFF_2_n10, state3FF_state_gff_4_SFF_2_n9,
         state3FF_state_gff_4_SFF_2_n7, state3FF_state_gff_4_SFF_2_n6,
         state3FF_state_gff_4_SFF_3_n11, state3FF_state_gff_4_SFF_3_n10,
         state3FF_state_gff_4_SFF_3_n9, state3FF_state_gff_4_SFF_3_n7,
         state3FF_state_gff_4_SFF_3_n6, state3FF_state_gff_5_SFF_0_n12,
         state3FF_state_gff_5_SFF_0_n11, state3FF_state_gff_5_SFF_0_n10,
         state3FF_state_gff_5_SFF_0_n8, state3FF_state_gff_5_SFF_0_n7,
         state3FF_state_gff_5_SFF_1_n12, state3FF_state_gff_5_SFF_1_n11,
         state3FF_state_gff_5_SFF_1_n10, state3FF_state_gff_5_SFF_1_n8,
         state3FF_state_gff_5_SFF_1_n7, state3FF_state_gff_5_SFF_2_n11,
         state3FF_state_gff_5_SFF_2_n10, state3FF_state_gff_5_SFF_2_n8,
         state3FF_state_gff_5_SFF_2_n7, state3FF_state_gff_5_SFF_3_n11,
         state3FF_state_gff_5_SFF_3_n10, state3FF_state_gff_5_SFF_3_n8,
         state3FF_state_gff_5_SFF_3_n7, state3FF_state_gff_6_SFF_0_n11,
         state3FF_state_gff_6_SFF_0_n10, state3FF_state_gff_6_SFF_0_n8,
         state3FF_state_gff_6_SFF_0_n7, state3FF_state_gff_6_SFF_1_n11,
         state3FF_state_gff_6_SFF_1_n10, state3FF_state_gff_6_SFF_1_n8,
         state3FF_state_gff_6_SFF_1_n7, state3FF_state_gff_6_SFF_2_n11,
         state3FF_state_gff_6_SFF_2_n10, state3FF_state_gff_6_SFF_2_n8,
         state3FF_state_gff_6_SFF_2_n7, state3FF_state_gff_6_SFF_3_n11,
         state3FF_state_gff_6_SFF_3_n10, state3FF_state_gff_6_SFF_3_n8,
         state3FF_state_gff_6_SFF_3_n7, state3FF_state_gff_7_SFF_0_n11,
         state3FF_state_gff_7_SFF_0_n10, state3FF_state_gff_7_SFF_0_n8,
         state3FF_state_gff_7_SFF_0_n7, state3FF_state_gff_7_SFF_1_n11,
         state3FF_state_gff_7_SFF_1_n10, state3FF_state_gff_7_SFF_1_n8,
         state3FF_state_gff_7_SFF_1_n7, state3FF_state_gff_7_SFF_2_n11,
         state3FF_state_gff_7_SFF_2_n10, state3FF_state_gff_7_SFF_2_n9,
         state3FF_state_gff_7_SFF_2_n7, state3FF_state_gff_7_SFF_2_n6,
         state3FF_state_gff_7_SFF_3_n11, state3FF_state_gff_7_SFF_3_n10,
         state3FF_state_gff_7_SFF_3_n9, state3FF_state_gff_7_SFF_3_n7,
         state3FF_state_gff_7_SFF_3_n6, state3FF_state_gff_8_SFF_0_n11,
         state3FF_state_gff_8_SFF_0_n10, state3FF_state_gff_8_SFF_0_n9,
         state3FF_state_gff_8_SFF_0_n7, state3FF_state_gff_8_SFF_0_n6,
         state3FF_state_gff_8_SFF_1_n11, state3FF_state_gff_8_SFF_1_n10,
         state3FF_state_gff_8_SFF_1_n9, state3FF_state_gff_8_SFF_1_n7,
         state3FF_state_gff_8_SFF_1_n6, state3FF_state_gff_8_SFF_2_n11,
         state3FF_state_gff_8_SFF_2_n10, state3FF_state_gff_8_SFF_2_n9,
         state3FF_state_gff_8_SFF_2_n7, state3FF_state_gff_8_SFF_2_n6,
         state3FF_state_gff_8_SFF_3_n11, state3FF_state_gff_8_SFF_3_n10,
         state3FF_state_gff_8_SFF_3_n9, state3FF_state_gff_8_SFF_3_n7,
         state3FF_state_gff_8_SFF_3_n6, state3FF_state_gff_9_SFF_0_n12,
         state3FF_state_gff_9_SFF_0_n11, state3FF_state_gff_9_SFF_0_n10,
         state3FF_state_gff_9_SFF_0_n8, state3FF_state_gff_9_SFF_0_n7,
         state3FF_state_gff_9_SFF_1_n12, state3FF_state_gff_9_SFF_1_n11,
         state3FF_state_gff_9_SFF_1_n10, state3FF_state_gff_9_SFF_1_n8,
         state3FF_state_gff_9_SFF_1_n7, state3FF_state_gff_9_SFF_2_n12,
         state3FF_state_gff_9_SFF_2_n11, state3FF_state_gff_9_SFF_2_n10,
         state3FF_state_gff_9_SFF_2_n8, state3FF_state_gff_9_SFF_2_n7,
         state3FF_state_gff_9_SFF_3_n12, state3FF_state_gff_9_SFF_3_n11,
         state3FF_state_gff_9_SFF_3_n10, state3FF_state_gff_9_SFF_3_n8,
         state3FF_state_gff_9_SFF_3_n7, state3FF_state_gff_10_SFF_0_n12,
         state3FF_state_gff_10_SFF_0_n11, state3FF_state_gff_10_SFF_0_n10,
         state3FF_state_gff_10_SFF_0_n8, state3FF_state_gff_10_SFF_0_n7,
         state3FF_state_gff_10_SFF_1_n12, state3FF_state_gff_10_SFF_1_n11,
         state3FF_state_gff_10_SFF_1_n10, state3FF_state_gff_10_SFF_1_n8,
         state3FF_state_gff_10_SFF_1_n7, state3FF_state_gff_10_SFF_2_n12,
         state3FF_state_gff_10_SFF_2_n11, state3FF_state_gff_10_SFF_2_n10,
         state3FF_state_gff_10_SFF_2_n8, state3FF_state_gff_10_SFF_2_n7,
         state3FF_state_gff_10_SFF_3_n12, state3FF_state_gff_10_SFF_3_n11,
         state3FF_state_gff_10_SFF_3_n10, state3FF_state_gff_10_SFF_3_n8,
         state3FF_state_gff_10_SFF_3_n7, state3FF_state_gff_11_SFF_0_n11,
         state3FF_state_gff_11_SFF_0_n10, state3FF_state_gff_11_SFF_0_n8,
         state3FF_state_gff_11_SFF_0_n7, state3FF_state_gff_11_SFF_1_n11,
         state3FF_state_gff_11_SFF_1_n10, state3FF_state_gff_11_SFF_1_n8,
         state3FF_state_gff_11_SFF_1_n7, state3FF_state_gff_11_SFF_2_n11,
         state3FF_state_gff_11_SFF_2_n10, state3FF_state_gff_11_SFF_2_n9,
         state3FF_state_gff_11_SFF_2_n7, state3FF_state_gff_11_SFF_2_n6,
         state3FF_state_gff_11_SFF_3_n11, state3FF_state_gff_11_SFF_3_n10,
         state3FF_state_gff_11_SFF_3_n9, state3FF_state_gff_11_SFF_3_n7,
         state3FF_state_gff_11_SFF_3_n6, state3FF_state_gff_12_SFF_0_n11,
         state3FF_state_gff_12_SFF_0_n10, state3FF_state_gff_12_SFF_0_n9,
         state3FF_state_gff_12_SFF_0_n7, state3FF_state_gff_12_SFF_0_n6,
         state3FF_state_gff_12_SFF_1_n11, state3FF_state_gff_12_SFF_1_n10,
         state3FF_state_gff_12_SFF_1_n9, state3FF_state_gff_12_SFF_1_n7,
         state3FF_state_gff_12_SFF_1_n6, state3FF_state_gff_12_SFF_2_n10,
         state3FF_state_gff_12_SFF_2_n9, state3FF_state_gff_12_SFF_2_n7,
         state3FF_state_gff_12_SFF_2_n6, state3FF_state_gff_12_SFF_3_n10,
         state3FF_state_gff_12_SFF_3_n9, state3FF_state_gff_12_SFF_3_n7,
         state3FF_state_gff_12_SFF_3_n6, state3FF_state_gff_13_SFF_0_n12,
         state3FF_state_gff_13_SFF_0_n11, state3FF_state_gff_13_SFF_0_n10,
         state3FF_state_gff_13_SFF_0_n8, state3FF_state_gff_13_SFF_0_n7,
         state3FF_state_gff_13_SFF_1_n12, state3FF_state_gff_13_SFF_1_n11,
         state3FF_state_gff_13_SFF_1_n10, state3FF_state_gff_13_SFF_1_n8,
         state3FF_state_gff_13_SFF_1_n7, state3FF_state_gff_13_SFF_2_n11,
         state3FF_state_gff_13_SFF_2_n10, state3FF_state_gff_13_SFF_2_n8,
         state3FF_state_gff_13_SFF_2_n7, state3FF_state_gff_13_SFF_3_n11,
         state3FF_state_gff_13_SFF_3_n10, state3FF_state_gff_13_SFF_3_n8,
         state3FF_state_gff_13_SFF_3_n7, state3FF_state_gff_14_SFF_0_n11,
         state3FF_state_gff_14_SFF_0_n10, state3FF_state_gff_14_SFF_0_n8,
         state3FF_state_gff_14_SFF_0_n7, state3FF_state_gff_14_SFF_1_n11,
         state3FF_state_gff_14_SFF_1_n10, state3FF_state_gff_14_SFF_1_n8,
         state3FF_state_gff_14_SFF_1_n7, state3FF_state_gff_14_SFF_2_n11,
         state3FF_state_gff_14_SFF_2_n10, state3FF_state_gff_14_SFF_2_n8,
         state3FF_state_gff_14_SFF_2_n7, state3FF_state_gff_14_SFF_3_n11,
         state3FF_state_gff_14_SFF_3_n10, state3FF_state_gff_14_SFF_3_n8,
         state3FF_state_gff_14_SFF_3_n7, state3FF_state_gff_15_SFF_0_n11,
         state3FF_state_gff_15_SFF_0_n10, state3FF_state_gff_15_SFF_0_n8,
         state3FF_state_gff_15_SFF_0_n7, state3FF_state_gff_15_SFF_1_n11,
         state3FF_state_gff_15_SFF_1_n10, state3FF_state_gff_15_SFF_1_n8,
         state3FF_state_gff_15_SFF_1_n7, state3FF_state_gff_15_SFF_2_n11,
         state3FF_state_gff_15_SFF_2_n10, state3FF_state_gff_15_SFF_2_n9,
         state3FF_state_gff_15_SFF_2_n7, state3FF_state_gff_15_SFF_2_n6,
         state3FF_state_gff_15_SFF_3_n11, state3FF_state_gff_15_SFF_3_n10,
         state3FF_state_gff_15_SFF_3_n9, state3FF_state_gff_15_SFF_3_n7,
         state3FF_state_gff_15_SFF_3_n6, state3FF_state_gff_16_SFF_0_n10,
         state3FF_state_gff_16_SFF_0_n9, state3FF_state_gff_16_SFF_0_n7,
         state3FF_state_gff_16_SFF_0_n6, state3FF_state_gff_16_SFF_1_n10,
         state3FF_state_gff_16_SFF_1_n9, state3FF_state_gff_16_SFF_1_n7,
         state3FF_state_gff_16_SFF_1_n6, state3FF_state_gff_16_SFF_2_n10,
         state3FF_state_gff_16_SFF_2_n9, state3FF_state_gff_16_SFF_2_n7,
         state3FF_state_gff_16_SFF_2_n6, state3FF_state_gff_16_SFF_3_n10,
         state3FF_state_gff_16_SFF_3_n9, state3FF_state_gff_16_SFF_3_n7,
         state3FF_state_gff_16_SFF_3_n6, key1FF_n4, key1FF_n3, key1FF_n2,
         key1FF_n1, key1FF_keystate_n18, key1FF_keystate_n17,
         key1FF_keystate_n16, key1FF_keystate_n15, key1FF_keystate_n14,
         key1FF_keystate_n13, key1FF_keystate_n12, key1FF_keystate_n11,
         key1FF_keystate_n10, key1FF_keystate_gff_1_SFF_0_n12,
         key1FF_keystate_gff_1_SFF_0_n11, key1FF_keystate_gff_1_SFF_0_n10,
         key1FF_keystate_gff_1_SFF_0_n8, key1FF_keystate_gff_1_SFF_0_n7,
         key1FF_keystate_gff_1_SFF_1_n12, key1FF_keystate_gff_1_SFF_1_n11,
         key1FF_keystate_gff_1_SFF_1_n10, key1FF_keystate_gff_1_SFF_1_n8,
         key1FF_keystate_gff_1_SFF_1_n7, key1FF_keystate_gff_1_SFF_2_n12,
         key1FF_keystate_gff_1_SFF_2_n11, key1FF_keystate_gff_1_SFF_2_n10,
         key1FF_keystate_gff_1_SFF_2_n8, key1FF_keystate_gff_1_SFF_2_n7,
         key1FF_keystate_gff_1_SFF_3_n12, key1FF_keystate_gff_1_SFF_3_n11,
         key1FF_keystate_gff_1_SFF_3_n10, key1FF_keystate_gff_1_SFF_3_n8,
         key1FF_keystate_gff_1_SFF_3_n7, key1FF_keystate_gff_2_SFF_0_n12,
         key1FF_keystate_gff_2_SFF_0_n11, key1FF_keystate_gff_2_SFF_0_n10,
         key1FF_keystate_gff_2_SFF_0_n8, key1FF_keystate_gff_2_SFF_0_n7,
         key1FF_keystate_gff_2_SFF_1_n12, key1FF_keystate_gff_2_SFF_1_n11,
         key1FF_keystate_gff_2_SFF_1_n10, key1FF_keystate_gff_2_SFF_1_n8,
         key1FF_keystate_gff_2_SFF_1_n7, key1FF_keystate_gff_2_SFF_2_n12,
         key1FF_keystate_gff_2_SFF_2_n11, key1FF_keystate_gff_2_SFF_2_n10,
         key1FF_keystate_gff_2_SFF_2_n8, key1FF_keystate_gff_2_SFF_2_n7,
         key1FF_keystate_gff_2_SFF_3_n12, key1FF_keystate_gff_2_SFF_3_n11,
         key1FF_keystate_gff_2_SFF_3_n10, key1FF_keystate_gff_2_SFF_3_n8,
         key1FF_keystate_gff_2_SFF_3_n7, key1FF_keystate_gff_3_SFF_0_n12,
         key1FF_keystate_gff_3_SFF_0_n11, key1FF_keystate_gff_3_SFF_0_n10,
         key1FF_keystate_gff_3_SFF_0_n8, key1FF_keystate_gff_3_SFF_0_n7,
         key1FF_keystate_gff_3_SFF_1_n12, key1FF_keystate_gff_3_SFF_1_n11,
         key1FF_keystate_gff_3_SFF_1_n10, key1FF_keystate_gff_3_SFF_1_n8,
         key1FF_keystate_gff_3_SFF_1_n7, key1FF_keystate_gff_3_SFF_2_n11,
         key1FF_keystate_gff_3_SFF_2_n10, key1FF_keystate_gff_3_SFF_2_n9,
         key1FF_keystate_gff_3_SFF_2_n7, key1FF_keystate_gff_3_SFF_2_n6,
         key1FF_keystate_gff_3_SFF_3_n11, key1FF_keystate_gff_3_SFF_3_n10,
         key1FF_keystate_gff_3_SFF_3_n9, key1FF_keystate_gff_3_SFF_3_n7,
         key1FF_keystate_gff_3_SFF_3_n6, key1FF_keystate_gff_4_SFF_0_n11,
         key1FF_keystate_gff_4_SFF_0_n10, key1FF_keystate_gff_4_SFF_0_n9,
         key1FF_keystate_gff_4_SFF_0_n7, key1FF_keystate_gff_4_SFF_0_n6,
         key1FF_keystate_gff_4_SFF_1_n11, key1FF_keystate_gff_4_SFF_1_n10,
         key1FF_keystate_gff_4_SFF_1_n9, key1FF_keystate_gff_4_SFF_1_n7,
         key1FF_keystate_gff_4_SFF_1_n6, key1FF_keystate_gff_4_SFF_2_n11,
         key1FF_keystate_gff_4_SFF_2_n10, key1FF_keystate_gff_4_SFF_2_n9,
         key1FF_keystate_gff_4_SFF_2_n7, key1FF_keystate_gff_4_SFF_2_n6,
         key1FF_keystate_gff_4_SFF_3_n11, key1FF_keystate_gff_4_SFF_3_n10,
         key1FF_keystate_gff_4_SFF_3_n9, key1FF_keystate_gff_4_SFF_3_n7,
         key1FF_keystate_gff_4_SFF_3_n6, key1FF_keystate_gff_5_SFF_0_n12,
         key1FF_keystate_gff_5_SFF_0_n11, key1FF_keystate_gff_5_SFF_0_n10,
         key1FF_keystate_gff_5_SFF_0_n8, key1FF_keystate_gff_5_SFF_0_n7,
         key1FF_keystate_gff_5_SFF_1_n12, key1FF_keystate_gff_5_SFF_1_n11,
         key1FF_keystate_gff_5_SFF_1_n10, key1FF_keystate_gff_5_SFF_1_n8,
         key1FF_keystate_gff_5_SFF_1_n7, key1FF_keystate_gff_5_SFF_2_n11,
         key1FF_keystate_gff_5_SFF_2_n10, key1FF_keystate_gff_5_SFF_2_n8,
         key1FF_keystate_gff_5_SFF_2_n7, key1FF_keystate_gff_5_SFF_3_n11,
         key1FF_keystate_gff_5_SFF_3_n10, key1FF_keystate_gff_5_SFF_3_n8,
         key1FF_keystate_gff_5_SFF_3_n7, key1FF_keystate_gff_6_SFF_0_n11,
         key1FF_keystate_gff_6_SFF_0_n10, key1FF_keystate_gff_6_SFF_0_n8,
         key1FF_keystate_gff_6_SFF_0_n7, key1FF_keystate_gff_6_SFF_1_n11,
         key1FF_keystate_gff_6_SFF_1_n10, key1FF_keystate_gff_6_SFF_1_n8,
         key1FF_keystate_gff_6_SFF_1_n7, key1FF_keystate_gff_6_SFF_2_n11,
         key1FF_keystate_gff_6_SFF_2_n10, key1FF_keystate_gff_6_SFF_2_n8,
         key1FF_keystate_gff_6_SFF_2_n7, key1FF_keystate_gff_6_SFF_3_n11,
         key1FF_keystate_gff_6_SFF_3_n10, key1FF_keystate_gff_6_SFF_3_n8,
         key1FF_keystate_gff_6_SFF_3_n7, key1FF_keystate_gff_7_SFF_0_n12,
         key1FF_keystate_gff_7_SFF_0_n11, key1FF_keystate_gff_7_SFF_0_n10,
         key1FF_keystate_gff_7_SFF_0_n8, key1FF_keystate_gff_7_SFF_0_n7,
         key1FF_keystate_gff_7_SFF_1_n12, key1FF_keystate_gff_7_SFF_1_n11,
         key1FF_keystate_gff_7_SFF_1_n10, key1FF_keystate_gff_7_SFF_1_n8,
         key1FF_keystate_gff_7_SFF_1_n7, key1FF_keystate_gff_7_SFF_2_n11,
         key1FF_keystate_gff_7_SFF_2_n10, key1FF_keystate_gff_7_SFF_2_n9,
         key1FF_keystate_gff_7_SFF_2_n7, key1FF_keystate_gff_7_SFF_2_n6,
         key1FF_keystate_gff_7_SFF_3_n11, key1FF_keystate_gff_7_SFF_3_n10,
         key1FF_keystate_gff_7_SFF_3_n9, key1FF_keystate_gff_7_SFF_3_n7,
         key1FF_keystate_gff_7_SFF_3_n6, key1FF_keystate_gff_8_SFF_0_n11,
         key1FF_keystate_gff_8_SFF_0_n10, key1FF_keystate_gff_8_SFF_0_n9,
         key1FF_keystate_gff_8_SFF_0_n7, key1FF_keystate_gff_8_SFF_0_n6,
         key1FF_keystate_gff_8_SFF_1_n11, key1FF_keystate_gff_8_SFF_1_n10,
         key1FF_keystate_gff_8_SFF_1_n9, key1FF_keystate_gff_8_SFF_1_n7,
         key1FF_keystate_gff_8_SFF_1_n6, key1FF_keystate_gff_8_SFF_2_n11,
         key1FF_keystate_gff_8_SFF_2_n10, key1FF_keystate_gff_8_SFF_2_n9,
         key1FF_keystate_gff_8_SFF_2_n7, key1FF_keystate_gff_8_SFF_2_n6,
         key1FF_keystate_gff_8_SFF_3_n11, key1FF_keystate_gff_8_SFF_3_n10,
         key1FF_keystate_gff_8_SFF_3_n9, key1FF_keystate_gff_8_SFF_3_n7,
         key1FF_keystate_gff_8_SFF_3_n6, key1FF_keystate_gff_9_SFF_0_n12,
         key1FF_keystate_gff_9_SFF_0_n11, key1FF_keystate_gff_9_SFF_0_n10,
         key1FF_keystate_gff_9_SFF_0_n8, key1FF_keystate_gff_9_SFF_0_n7,
         key1FF_keystate_gff_9_SFF_1_n12, key1FF_keystate_gff_9_SFF_1_n11,
         key1FF_keystate_gff_9_SFF_1_n10, key1FF_keystate_gff_9_SFF_1_n8,
         key1FF_keystate_gff_9_SFF_1_n7, key1FF_keystate_gff_9_SFF_2_n12,
         key1FF_keystate_gff_9_SFF_2_n11, key1FF_keystate_gff_9_SFF_2_n10,
         key1FF_keystate_gff_9_SFF_2_n8, key1FF_keystate_gff_9_SFF_2_n7,
         key1FF_keystate_gff_9_SFF_3_n12, key1FF_keystate_gff_9_SFF_3_n11,
         key1FF_keystate_gff_9_SFF_3_n10, key1FF_keystate_gff_9_SFF_3_n8,
         key1FF_keystate_gff_9_SFF_3_n7, key1FF_keystate_gff_10_SFF_0_n12,
         key1FF_keystate_gff_10_SFF_0_n11, key1FF_keystate_gff_10_SFF_0_n10,
         key1FF_keystate_gff_10_SFF_0_n8, key1FF_keystate_gff_10_SFF_0_n7,
         key1FF_keystate_gff_10_SFF_1_n12, key1FF_keystate_gff_10_SFF_1_n11,
         key1FF_keystate_gff_10_SFF_1_n10, key1FF_keystate_gff_10_SFF_1_n8,
         key1FF_keystate_gff_10_SFF_1_n7, key1FF_keystate_gff_10_SFF_2_n12,
         key1FF_keystate_gff_10_SFF_2_n11, key1FF_keystate_gff_10_SFF_2_n10,
         key1FF_keystate_gff_10_SFF_2_n8, key1FF_keystate_gff_10_SFF_2_n7,
         key1FF_keystate_gff_10_SFF_3_n12, key1FF_keystate_gff_10_SFF_3_n11,
         key1FF_keystate_gff_10_SFF_3_n10, key1FF_keystate_gff_10_SFF_3_n8,
         key1FF_keystate_gff_10_SFF_3_n7, key1FF_keystate_gff_11_SFF_0_n11,
         key1FF_keystate_gff_11_SFF_0_n10, key1FF_keystate_gff_11_SFF_0_n8,
         key1FF_keystate_gff_11_SFF_0_n7, key1FF_keystate_gff_11_SFF_1_n11,
         key1FF_keystate_gff_11_SFF_1_n10, key1FF_keystate_gff_11_SFF_1_n8,
         key1FF_keystate_gff_11_SFF_1_n7, key1FF_keystate_gff_11_SFF_2_n11,
         key1FF_keystate_gff_11_SFF_2_n10, key1FF_keystate_gff_11_SFF_2_n9,
         key1FF_keystate_gff_11_SFF_2_n7, key1FF_keystate_gff_11_SFF_2_n6,
         key1FF_keystate_gff_11_SFF_3_n11, key1FF_keystate_gff_11_SFF_3_n10,
         key1FF_keystate_gff_11_SFF_3_n9, key1FF_keystate_gff_11_SFF_3_n7,
         key1FF_keystate_gff_11_SFF_3_n6, key1FF_keystate_gff_12_SFF_0_n11,
         key1FF_keystate_gff_12_SFF_0_n10, key1FF_keystate_gff_12_SFF_0_n9,
         key1FF_keystate_gff_12_SFF_0_n7, key1FF_keystate_gff_12_SFF_0_n6,
         key1FF_keystate_gff_12_SFF_1_n11, key1FF_keystate_gff_12_SFF_1_n10,
         key1FF_keystate_gff_12_SFF_1_n9, key1FF_keystate_gff_12_SFF_1_n7,
         key1FF_keystate_gff_12_SFF_1_n6, key1FF_keystate_gff_12_SFF_2_n11,
         key1FF_keystate_gff_12_SFF_2_n10, key1FF_keystate_gff_12_SFF_2_n9,
         key1FF_keystate_gff_12_SFF_2_n7, key1FF_keystate_gff_12_SFF_2_n6,
         key1FF_keystate_gff_12_SFF_3_n11, key1FF_keystate_gff_12_SFF_3_n10,
         key1FF_keystate_gff_12_SFF_3_n9, key1FF_keystate_gff_12_SFF_3_n7,
         key1FF_keystate_gff_12_SFF_3_n6, key1FF_keystate_gff_13_SFF_0_n12,
         key1FF_keystate_gff_13_SFF_0_n11, key1FF_keystate_gff_13_SFF_0_n10,
         key1FF_keystate_gff_13_SFF_0_n8, key1FF_keystate_gff_13_SFF_0_n7,
         key1FF_keystate_gff_13_SFF_1_n12, key1FF_keystate_gff_13_SFF_1_n11,
         key1FF_keystate_gff_13_SFF_1_n10, key1FF_keystate_gff_13_SFF_1_n8,
         key1FF_keystate_gff_13_SFF_1_n7, key1FF_keystate_gff_13_SFF_2_n11,
         key1FF_keystate_gff_13_SFF_2_n10, key1FF_keystate_gff_13_SFF_2_n8,
         key1FF_keystate_gff_13_SFF_2_n7, key1FF_keystate_gff_13_SFF_3_n11,
         key1FF_keystate_gff_13_SFF_3_n10, key1FF_keystate_gff_13_SFF_3_n8,
         key1FF_keystate_gff_13_SFF_3_n7, key1FF_keystate_gff_14_SFF_0_n11,
         key1FF_keystate_gff_14_SFF_0_n10, key1FF_keystate_gff_14_SFF_0_n8,
         key1FF_keystate_gff_14_SFF_0_n7, key1FF_keystate_gff_14_SFF_1_n11,
         key1FF_keystate_gff_14_SFF_1_n10, key1FF_keystate_gff_14_SFF_1_n8,
         key1FF_keystate_gff_14_SFF_1_n7, key1FF_keystate_gff_14_SFF_2_n11,
         key1FF_keystate_gff_14_SFF_2_n10, key1FF_keystate_gff_14_SFF_2_n8,
         key1FF_keystate_gff_14_SFF_2_n7, key1FF_keystate_gff_14_SFF_3_n11,
         key1FF_keystate_gff_14_SFF_3_n10, key1FF_keystate_gff_14_SFF_3_n8,
         key1FF_keystate_gff_14_SFF_3_n7, key1FF_keystate_gff_15_SFF_0_n11,
         key1FF_keystate_gff_15_SFF_0_n10, key1FF_keystate_gff_15_SFF_0_n8,
         key1FF_keystate_gff_15_SFF_0_n7, key1FF_keystate_gff_15_SFF_1_n11,
         key1FF_keystate_gff_15_SFF_1_n10, key1FF_keystate_gff_15_SFF_1_n8,
         key1FF_keystate_gff_15_SFF_1_n7, key1FF_keystate_gff_15_SFF_2_n11,
         key1FF_keystate_gff_15_SFF_2_n10, key1FF_keystate_gff_15_SFF_2_n9,
         key1FF_keystate_gff_15_SFF_2_n7, key1FF_keystate_gff_15_SFF_2_n6,
         key1FF_keystate_gff_15_SFF_3_n11, key1FF_keystate_gff_15_SFF_3_n10,
         key1FF_keystate_gff_15_SFF_3_n9, key1FF_keystate_gff_15_SFF_3_n7,
         key1FF_keystate_gff_15_SFF_3_n6, key1FF_keystate_gff_16_SFF_0_n11,
         key1FF_keystate_gff_16_SFF_0_n10, key1FF_keystate_gff_16_SFF_0_n9,
         key1FF_keystate_gff_16_SFF_0_n7, key1FF_keystate_gff_16_SFF_0_n6,
         key1FF_keystate_gff_16_SFF_1_n11, key1FF_keystate_gff_16_SFF_1_n10,
         key1FF_keystate_gff_16_SFF_1_n9, key1FF_keystate_gff_16_SFF_1_n7,
         key1FF_keystate_gff_16_SFF_1_n6, key1FF_keystate_gff_16_SFF_2_n10,
         key1FF_keystate_gff_16_SFF_2_n9, key1FF_keystate_gff_16_SFF_2_n7,
         key1FF_keystate_gff_16_SFF_2_n6, key1FF_keystate_gff_16_SFF_3_n10,
         key1FF_keystate_gff_16_SFF_3_n9, key1FF_keystate_gff_16_SFF_3_n7,
         key1FF_keystate_gff_16_SFF_3_n6, key1FF_keystate_gff_17_SFF_0_n12,
         key1FF_keystate_gff_17_SFF_0_n11, key1FF_keystate_gff_17_SFF_0_n10,
         key1FF_keystate_gff_17_SFF_0_n8, key1FF_keystate_gff_17_SFF_0_n7,
         key1FF_keystate_gff_17_SFF_1_n12, key1FF_keystate_gff_17_SFF_1_n11,
         key1FF_keystate_gff_17_SFF_1_n10, key1FF_keystate_gff_17_SFF_1_n8,
         key1FF_keystate_gff_17_SFF_1_n7, key1FF_keystate_gff_17_SFF_2_n11,
         key1FF_keystate_gff_17_SFF_2_n10, key1FF_keystate_gff_17_SFF_2_n8,
         key1FF_keystate_gff_17_SFF_2_n7, key1FF_keystate_gff_17_SFF_3_n11,
         key1FF_keystate_gff_17_SFF_3_n10, key1FF_keystate_gff_17_SFF_3_n8,
         key1FF_keystate_gff_17_SFF_3_n7, key1FF_keystate_gff_18_SFF_0_n11,
         key1FF_keystate_gff_18_SFF_0_n10, key1FF_keystate_gff_18_SFF_0_n8,
         key1FF_keystate_gff_18_SFF_0_n7, key1FF_keystate_gff_18_SFF_1_n11,
         key1FF_keystate_gff_18_SFF_1_n10, key1FF_keystate_gff_18_SFF_1_n8,
         key1FF_keystate_gff_18_SFF_1_n7, key1FF_keystate_gff_18_SFF_2_n11,
         key1FF_keystate_gff_18_SFF_2_n10, key1FF_keystate_gff_18_SFF_2_n8,
         key1FF_keystate_gff_18_SFF_2_n7, key1FF_keystate_gff_18_SFF_3_n11,
         key1FF_keystate_gff_18_SFF_3_n10, key1FF_keystate_gff_18_SFF_3_n8,
         key1FF_keystate_gff_18_SFF_3_n7, key1FF_keystate_gff_19_SFF_0_n11,
         key1FF_keystate_gff_19_SFF_0_n10, key1FF_keystate_gff_19_SFF_0_n8,
         key1FF_keystate_gff_19_SFF_0_n7, key1FF_keystate_gff_19_SFF_1_n11,
         key1FF_keystate_gff_19_SFF_1_n10, key1FF_keystate_gff_19_SFF_1_n8,
         key1FF_keystate_gff_19_SFF_1_n7, key1FF_keystate_gff_19_SFF_2_n11,
         key1FF_keystate_gff_19_SFF_2_n10, key1FF_keystate_gff_19_SFF_2_n9,
         key1FF_keystate_gff_19_SFF_2_n7, key1FF_keystate_gff_19_SFF_2_n6,
         key1FF_keystate_gff_19_SFF_3_n11, key1FF_keystate_gff_19_SFF_3_n10,
         key1FF_keystate_gff_19_SFF_3_n9, key1FF_keystate_gff_19_SFF_3_n7,
         key1FF_keystate_gff_19_SFF_3_n6, key1FF_keystate_gff_20_SFF_0_n10,
         key1FF_keystate_gff_20_SFF_0_n9, key1FF_keystate_gff_20_SFF_0_n7,
         key1FF_keystate_gff_20_SFF_0_n6, key1FF_keystate_gff_20_SFF_1_n10,
         key1FF_keystate_gff_20_SFF_1_n9, key1FF_keystate_gff_20_SFF_1_n7,
         key1FF_keystate_gff_20_SFF_1_n6, key1FF_keystate_gff_20_SFF_2_n10,
         key1FF_keystate_gff_20_SFF_2_n9, key1FF_keystate_gff_20_SFF_2_n7,
         key1FF_keystate_gff_20_SFF_2_n6, key1FF_keystate_gff_20_SFF_3_n10,
         key1FF_keystate_gff_20_SFF_3_n9, key1FF_keystate_gff_20_SFF_3_n7,
         key1FF_keystate_gff_20_SFF_3_n6, key2FF_n4, key2FF_n3, key2FF_n2,
         key2FF_n1, key2FF_keystate_n18, key2FF_keystate_n17,
         key2FF_keystate_n16, key2FF_keystate_n15, key2FF_keystate_n14,
         key2FF_keystate_n13, key2FF_keystate_n12, key2FF_keystate_n11,
         key2FF_keystate_n10, key2FF_keystate_gff_1_SFF_0_n12,
         key2FF_keystate_gff_1_SFF_0_n11, key2FF_keystate_gff_1_SFF_0_n10,
         key2FF_keystate_gff_1_SFF_0_n8, key2FF_keystate_gff_1_SFF_0_n7,
         key2FF_keystate_gff_1_SFF_1_n12, key2FF_keystate_gff_1_SFF_1_n11,
         key2FF_keystate_gff_1_SFF_1_n10, key2FF_keystate_gff_1_SFF_1_n8,
         key2FF_keystate_gff_1_SFF_1_n7, key2FF_keystate_gff_1_SFF_2_n12,
         key2FF_keystate_gff_1_SFF_2_n11, key2FF_keystate_gff_1_SFF_2_n10,
         key2FF_keystate_gff_1_SFF_2_n8, key2FF_keystate_gff_1_SFF_2_n7,
         key2FF_keystate_gff_1_SFF_3_n12, key2FF_keystate_gff_1_SFF_3_n11,
         key2FF_keystate_gff_1_SFF_3_n10, key2FF_keystate_gff_1_SFF_3_n8,
         key2FF_keystate_gff_1_SFF_3_n7, key2FF_keystate_gff_2_SFF_0_n12,
         key2FF_keystate_gff_2_SFF_0_n11, key2FF_keystate_gff_2_SFF_0_n10,
         key2FF_keystate_gff_2_SFF_0_n8, key2FF_keystate_gff_2_SFF_0_n7,
         key2FF_keystate_gff_2_SFF_1_n12, key2FF_keystate_gff_2_SFF_1_n11,
         key2FF_keystate_gff_2_SFF_1_n10, key2FF_keystate_gff_2_SFF_1_n8,
         key2FF_keystate_gff_2_SFF_1_n7, key2FF_keystate_gff_2_SFF_2_n12,
         key2FF_keystate_gff_2_SFF_2_n11, key2FF_keystate_gff_2_SFF_2_n10,
         key2FF_keystate_gff_2_SFF_2_n8, key2FF_keystate_gff_2_SFF_2_n7,
         key2FF_keystate_gff_2_SFF_3_n12, key2FF_keystate_gff_2_SFF_3_n11,
         key2FF_keystate_gff_2_SFF_3_n10, key2FF_keystate_gff_2_SFF_3_n8,
         key2FF_keystate_gff_2_SFF_3_n7, key2FF_keystate_gff_3_SFF_0_n12,
         key2FF_keystate_gff_3_SFF_0_n11, key2FF_keystate_gff_3_SFF_0_n10,
         key2FF_keystate_gff_3_SFF_0_n8, key2FF_keystate_gff_3_SFF_0_n7,
         key2FF_keystate_gff_3_SFF_1_n12, key2FF_keystate_gff_3_SFF_1_n11,
         key2FF_keystate_gff_3_SFF_1_n10, key2FF_keystate_gff_3_SFF_1_n8,
         key2FF_keystate_gff_3_SFF_1_n7, key2FF_keystate_gff_3_SFF_2_n11,
         key2FF_keystate_gff_3_SFF_2_n10, key2FF_keystate_gff_3_SFF_2_n9,
         key2FF_keystate_gff_3_SFF_2_n7, key2FF_keystate_gff_3_SFF_2_n6,
         key2FF_keystate_gff_3_SFF_3_n11, key2FF_keystate_gff_3_SFF_3_n10,
         key2FF_keystate_gff_3_SFF_3_n9, key2FF_keystate_gff_3_SFF_3_n7,
         key2FF_keystate_gff_3_SFF_3_n6, key2FF_keystate_gff_4_SFF_0_n11,
         key2FF_keystate_gff_4_SFF_0_n10, key2FF_keystate_gff_4_SFF_0_n9,
         key2FF_keystate_gff_4_SFF_0_n7, key2FF_keystate_gff_4_SFF_0_n6,
         key2FF_keystate_gff_4_SFF_1_n11, key2FF_keystate_gff_4_SFF_1_n10,
         key2FF_keystate_gff_4_SFF_1_n9, key2FF_keystate_gff_4_SFF_1_n7,
         key2FF_keystate_gff_4_SFF_1_n6, key2FF_keystate_gff_4_SFF_2_n11,
         key2FF_keystate_gff_4_SFF_2_n10, key2FF_keystate_gff_4_SFF_2_n9,
         key2FF_keystate_gff_4_SFF_2_n7, key2FF_keystate_gff_4_SFF_2_n6,
         key2FF_keystate_gff_4_SFF_3_n11, key2FF_keystate_gff_4_SFF_3_n10,
         key2FF_keystate_gff_4_SFF_3_n9, key2FF_keystate_gff_4_SFF_3_n7,
         key2FF_keystate_gff_4_SFF_3_n6, key2FF_keystate_gff_5_SFF_0_n12,
         key2FF_keystate_gff_5_SFF_0_n11, key2FF_keystate_gff_5_SFF_0_n10,
         key2FF_keystate_gff_5_SFF_0_n8, key2FF_keystate_gff_5_SFF_0_n7,
         key2FF_keystate_gff_5_SFF_1_n12, key2FF_keystate_gff_5_SFF_1_n11,
         key2FF_keystate_gff_5_SFF_1_n10, key2FF_keystate_gff_5_SFF_1_n8,
         key2FF_keystate_gff_5_SFF_1_n7, key2FF_keystate_gff_5_SFF_2_n11,
         key2FF_keystate_gff_5_SFF_2_n10, key2FF_keystate_gff_5_SFF_2_n8,
         key2FF_keystate_gff_5_SFF_2_n7, key2FF_keystate_gff_5_SFF_3_n11,
         key2FF_keystate_gff_5_SFF_3_n10, key2FF_keystate_gff_5_SFF_3_n8,
         key2FF_keystate_gff_5_SFF_3_n7, key2FF_keystate_gff_6_SFF_0_n11,
         key2FF_keystate_gff_6_SFF_0_n10, key2FF_keystate_gff_6_SFF_0_n8,
         key2FF_keystate_gff_6_SFF_0_n7, key2FF_keystate_gff_6_SFF_1_n11,
         key2FF_keystate_gff_6_SFF_1_n10, key2FF_keystate_gff_6_SFF_1_n8,
         key2FF_keystate_gff_6_SFF_1_n7, key2FF_keystate_gff_6_SFF_2_n11,
         key2FF_keystate_gff_6_SFF_2_n10, key2FF_keystate_gff_6_SFF_2_n8,
         key2FF_keystate_gff_6_SFF_2_n7, key2FF_keystate_gff_6_SFF_3_n11,
         key2FF_keystate_gff_6_SFF_3_n10, key2FF_keystate_gff_6_SFF_3_n8,
         key2FF_keystate_gff_6_SFF_3_n7, key2FF_keystate_gff_7_SFF_0_n12,
         key2FF_keystate_gff_7_SFF_0_n11, key2FF_keystate_gff_7_SFF_0_n10,
         key2FF_keystate_gff_7_SFF_0_n8, key2FF_keystate_gff_7_SFF_0_n7,
         key2FF_keystate_gff_7_SFF_1_n12, key2FF_keystate_gff_7_SFF_1_n11,
         key2FF_keystate_gff_7_SFF_1_n10, key2FF_keystate_gff_7_SFF_1_n8,
         key2FF_keystate_gff_7_SFF_1_n7, key2FF_keystate_gff_7_SFF_2_n11,
         key2FF_keystate_gff_7_SFF_2_n10, key2FF_keystate_gff_7_SFF_2_n9,
         key2FF_keystate_gff_7_SFF_2_n7, key2FF_keystate_gff_7_SFF_2_n6,
         key2FF_keystate_gff_7_SFF_3_n11, key2FF_keystate_gff_7_SFF_3_n10,
         key2FF_keystate_gff_7_SFF_3_n9, key2FF_keystate_gff_7_SFF_3_n7,
         key2FF_keystate_gff_7_SFF_3_n6, key2FF_keystate_gff_8_SFF_0_n11,
         key2FF_keystate_gff_8_SFF_0_n10, key2FF_keystate_gff_8_SFF_0_n9,
         key2FF_keystate_gff_8_SFF_0_n7, key2FF_keystate_gff_8_SFF_0_n6,
         key2FF_keystate_gff_8_SFF_1_n11, key2FF_keystate_gff_8_SFF_1_n10,
         key2FF_keystate_gff_8_SFF_1_n9, key2FF_keystate_gff_8_SFF_1_n7,
         key2FF_keystate_gff_8_SFF_1_n6, key2FF_keystate_gff_8_SFF_2_n11,
         key2FF_keystate_gff_8_SFF_2_n10, key2FF_keystate_gff_8_SFF_2_n9,
         key2FF_keystate_gff_8_SFF_2_n7, key2FF_keystate_gff_8_SFF_2_n6,
         key2FF_keystate_gff_8_SFF_3_n11, key2FF_keystate_gff_8_SFF_3_n10,
         key2FF_keystate_gff_8_SFF_3_n9, key2FF_keystate_gff_8_SFF_3_n7,
         key2FF_keystate_gff_8_SFF_3_n6, key2FF_keystate_gff_9_SFF_0_n12,
         key2FF_keystate_gff_9_SFF_0_n11, key2FF_keystate_gff_9_SFF_0_n10,
         key2FF_keystate_gff_9_SFF_0_n8, key2FF_keystate_gff_9_SFF_0_n7,
         key2FF_keystate_gff_9_SFF_1_n12, key2FF_keystate_gff_9_SFF_1_n11,
         key2FF_keystate_gff_9_SFF_1_n10, key2FF_keystate_gff_9_SFF_1_n8,
         key2FF_keystate_gff_9_SFF_1_n7, key2FF_keystate_gff_9_SFF_2_n12,
         key2FF_keystate_gff_9_SFF_2_n11, key2FF_keystate_gff_9_SFF_2_n10,
         key2FF_keystate_gff_9_SFF_2_n8, key2FF_keystate_gff_9_SFF_2_n7,
         key2FF_keystate_gff_9_SFF_3_n12, key2FF_keystate_gff_9_SFF_3_n11,
         key2FF_keystate_gff_9_SFF_3_n10, key2FF_keystate_gff_9_SFF_3_n8,
         key2FF_keystate_gff_9_SFF_3_n7, key2FF_keystate_gff_10_SFF_0_n12,
         key2FF_keystate_gff_10_SFF_0_n11, key2FF_keystate_gff_10_SFF_0_n10,
         key2FF_keystate_gff_10_SFF_0_n8, key2FF_keystate_gff_10_SFF_0_n7,
         key2FF_keystate_gff_10_SFF_1_n12, key2FF_keystate_gff_10_SFF_1_n11,
         key2FF_keystate_gff_10_SFF_1_n10, key2FF_keystate_gff_10_SFF_1_n8,
         key2FF_keystate_gff_10_SFF_1_n7, key2FF_keystate_gff_10_SFF_2_n12,
         key2FF_keystate_gff_10_SFF_2_n11, key2FF_keystate_gff_10_SFF_2_n10,
         key2FF_keystate_gff_10_SFF_2_n8, key2FF_keystate_gff_10_SFF_2_n7,
         key2FF_keystate_gff_10_SFF_3_n12, key2FF_keystate_gff_10_SFF_3_n11,
         key2FF_keystate_gff_10_SFF_3_n10, key2FF_keystate_gff_10_SFF_3_n8,
         key2FF_keystate_gff_10_SFF_3_n7, key2FF_keystate_gff_11_SFF_0_n11,
         key2FF_keystate_gff_11_SFF_0_n10, key2FF_keystate_gff_11_SFF_0_n8,
         key2FF_keystate_gff_11_SFF_0_n7, key2FF_keystate_gff_11_SFF_1_n11,
         key2FF_keystate_gff_11_SFF_1_n10, key2FF_keystate_gff_11_SFF_1_n8,
         key2FF_keystate_gff_11_SFF_1_n7, key2FF_keystate_gff_11_SFF_2_n11,
         key2FF_keystate_gff_11_SFF_2_n10, key2FF_keystate_gff_11_SFF_2_n9,
         key2FF_keystate_gff_11_SFF_2_n7, key2FF_keystate_gff_11_SFF_2_n6,
         key2FF_keystate_gff_11_SFF_3_n11, key2FF_keystate_gff_11_SFF_3_n10,
         key2FF_keystate_gff_11_SFF_3_n9, key2FF_keystate_gff_11_SFF_3_n7,
         key2FF_keystate_gff_11_SFF_3_n6, key2FF_keystate_gff_12_SFF_0_n11,
         key2FF_keystate_gff_12_SFF_0_n10, key2FF_keystate_gff_12_SFF_0_n9,
         key2FF_keystate_gff_12_SFF_0_n7, key2FF_keystate_gff_12_SFF_0_n6,
         key2FF_keystate_gff_12_SFF_1_n11, key2FF_keystate_gff_12_SFF_1_n10,
         key2FF_keystate_gff_12_SFF_1_n9, key2FF_keystate_gff_12_SFF_1_n7,
         key2FF_keystate_gff_12_SFF_1_n6, key2FF_keystate_gff_12_SFF_2_n11,
         key2FF_keystate_gff_12_SFF_2_n10, key2FF_keystate_gff_12_SFF_2_n9,
         key2FF_keystate_gff_12_SFF_2_n7, key2FF_keystate_gff_12_SFF_2_n6,
         key2FF_keystate_gff_12_SFF_3_n11, key2FF_keystate_gff_12_SFF_3_n10,
         key2FF_keystate_gff_12_SFF_3_n9, key2FF_keystate_gff_12_SFF_3_n7,
         key2FF_keystate_gff_12_SFF_3_n6, key2FF_keystate_gff_13_SFF_0_n12,
         key2FF_keystate_gff_13_SFF_0_n11, key2FF_keystate_gff_13_SFF_0_n10,
         key2FF_keystate_gff_13_SFF_0_n8, key2FF_keystate_gff_13_SFF_0_n7,
         key2FF_keystate_gff_13_SFF_1_n12, key2FF_keystate_gff_13_SFF_1_n11,
         key2FF_keystate_gff_13_SFF_1_n10, key2FF_keystate_gff_13_SFF_1_n8,
         key2FF_keystate_gff_13_SFF_1_n7, key2FF_keystate_gff_13_SFF_2_n11,
         key2FF_keystate_gff_13_SFF_2_n10, key2FF_keystate_gff_13_SFF_2_n8,
         key2FF_keystate_gff_13_SFF_2_n7, key2FF_keystate_gff_13_SFF_3_n11,
         key2FF_keystate_gff_13_SFF_3_n10, key2FF_keystate_gff_13_SFF_3_n8,
         key2FF_keystate_gff_13_SFF_3_n7, key2FF_keystate_gff_14_SFF_0_n11,
         key2FF_keystate_gff_14_SFF_0_n10, key2FF_keystate_gff_14_SFF_0_n8,
         key2FF_keystate_gff_14_SFF_0_n7, key2FF_keystate_gff_14_SFF_1_n11,
         key2FF_keystate_gff_14_SFF_1_n10, key2FF_keystate_gff_14_SFF_1_n8,
         key2FF_keystate_gff_14_SFF_1_n7, key2FF_keystate_gff_14_SFF_2_n11,
         key2FF_keystate_gff_14_SFF_2_n10, key2FF_keystate_gff_14_SFF_2_n8,
         key2FF_keystate_gff_14_SFF_2_n7, key2FF_keystate_gff_14_SFF_3_n11,
         key2FF_keystate_gff_14_SFF_3_n10, key2FF_keystate_gff_14_SFF_3_n8,
         key2FF_keystate_gff_14_SFF_3_n7, key2FF_keystate_gff_15_SFF_0_n11,
         key2FF_keystate_gff_15_SFF_0_n10, key2FF_keystate_gff_15_SFF_0_n8,
         key2FF_keystate_gff_15_SFF_0_n7, key2FF_keystate_gff_15_SFF_1_n11,
         key2FF_keystate_gff_15_SFF_1_n10, key2FF_keystate_gff_15_SFF_1_n8,
         key2FF_keystate_gff_15_SFF_1_n7, key2FF_keystate_gff_15_SFF_2_n11,
         key2FF_keystate_gff_15_SFF_2_n10, key2FF_keystate_gff_15_SFF_2_n9,
         key2FF_keystate_gff_15_SFF_2_n7, key2FF_keystate_gff_15_SFF_2_n6,
         key2FF_keystate_gff_15_SFF_3_n11, key2FF_keystate_gff_15_SFF_3_n10,
         key2FF_keystate_gff_15_SFF_3_n9, key2FF_keystate_gff_15_SFF_3_n7,
         key2FF_keystate_gff_15_SFF_3_n6, key2FF_keystate_gff_16_SFF_0_n11,
         key2FF_keystate_gff_16_SFF_0_n10, key2FF_keystate_gff_16_SFF_0_n9,
         key2FF_keystate_gff_16_SFF_0_n7, key2FF_keystate_gff_16_SFF_0_n6,
         key2FF_keystate_gff_16_SFF_1_n11, key2FF_keystate_gff_16_SFF_1_n10,
         key2FF_keystate_gff_16_SFF_1_n9, key2FF_keystate_gff_16_SFF_1_n7,
         key2FF_keystate_gff_16_SFF_1_n6, key2FF_keystate_gff_16_SFF_2_n10,
         key2FF_keystate_gff_16_SFF_2_n9, key2FF_keystate_gff_16_SFF_2_n7,
         key2FF_keystate_gff_16_SFF_2_n6, key2FF_keystate_gff_16_SFF_3_n10,
         key2FF_keystate_gff_16_SFF_3_n9, key2FF_keystate_gff_16_SFF_3_n7,
         key2FF_keystate_gff_16_SFF_3_n6, key2FF_keystate_gff_17_SFF_0_n12,
         key2FF_keystate_gff_17_SFF_0_n11, key2FF_keystate_gff_17_SFF_0_n10,
         key2FF_keystate_gff_17_SFF_0_n8, key2FF_keystate_gff_17_SFF_0_n7,
         key2FF_keystate_gff_17_SFF_1_n12, key2FF_keystate_gff_17_SFF_1_n11,
         key2FF_keystate_gff_17_SFF_1_n10, key2FF_keystate_gff_17_SFF_1_n8,
         key2FF_keystate_gff_17_SFF_1_n7, key2FF_keystate_gff_17_SFF_2_n11,
         key2FF_keystate_gff_17_SFF_2_n10, key2FF_keystate_gff_17_SFF_2_n8,
         key2FF_keystate_gff_17_SFF_2_n7, key2FF_keystate_gff_17_SFF_3_n11,
         key2FF_keystate_gff_17_SFF_3_n10, key2FF_keystate_gff_17_SFF_3_n8,
         key2FF_keystate_gff_17_SFF_3_n7, key2FF_keystate_gff_18_SFF_0_n11,
         key2FF_keystate_gff_18_SFF_0_n10, key2FF_keystate_gff_18_SFF_0_n8,
         key2FF_keystate_gff_18_SFF_0_n7, key2FF_keystate_gff_18_SFF_1_n11,
         key2FF_keystate_gff_18_SFF_1_n10, key2FF_keystate_gff_18_SFF_1_n8,
         key2FF_keystate_gff_18_SFF_1_n7, key2FF_keystate_gff_18_SFF_2_n11,
         key2FF_keystate_gff_18_SFF_2_n10, key2FF_keystate_gff_18_SFF_2_n8,
         key2FF_keystate_gff_18_SFF_2_n7, key2FF_keystate_gff_18_SFF_3_n11,
         key2FF_keystate_gff_18_SFF_3_n10, key2FF_keystate_gff_18_SFF_3_n8,
         key2FF_keystate_gff_18_SFF_3_n7, key2FF_keystate_gff_19_SFF_0_n11,
         key2FF_keystate_gff_19_SFF_0_n10, key2FF_keystate_gff_19_SFF_0_n8,
         key2FF_keystate_gff_19_SFF_0_n7, key2FF_keystate_gff_19_SFF_1_n11,
         key2FF_keystate_gff_19_SFF_1_n10, key2FF_keystate_gff_19_SFF_1_n8,
         key2FF_keystate_gff_19_SFF_1_n7, key2FF_keystate_gff_19_SFF_2_n11,
         key2FF_keystate_gff_19_SFF_2_n10, key2FF_keystate_gff_19_SFF_2_n9,
         key2FF_keystate_gff_19_SFF_2_n7, key2FF_keystate_gff_19_SFF_2_n6,
         key2FF_keystate_gff_19_SFF_3_n11, key2FF_keystate_gff_19_SFF_3_n10,
         key2FF_keystate_gff_19_SFF_3_n9, key2FF_keystate_gff_19_SFF_3_n7,
         key2FF_keystate_gff_19_SFF_3_n6, key2FF_keystate_gff_20_SFF_0_n10,
         key2FF_keystate_gff_20_SFF_0_n9, key2FF_keystate_gff_20_SFF_0_n7,
         key2FF_keystate_gff_20_SFF_0_n6, key2FF_keystate_gff_20_SFF_1_n10,
         key2FF_keystate_gff_20_SFF_1_n9, key2FF_keystate_gff_20_SFF_1_n7,
         key2FF_keystate_gff_20_SFF_1_n6, key2FF_keystate_gff_20_SFF_2_n10,
         key2FF_keystate_gff_20_SFF_2_n9, key2FF_keystate_gff_20_SFF_2_n7,
         key2FF_keystate_gff_20_SFF_2_n6, key2FF_keystate_gff_20_SFF_3_n10,
         key2FF_keystate_gff_20_SFF_3_n9, key2FF_keystate_gff_20_SFF_3_n7,
         key2FF_keystate_gff_20_SFF_3_n6, key3FF_n4, key3FF_n3, key3FF_n2,
         key3FF_n1, key3FF_keystate_n18, key3FF_keystate_n17,
         key3FF_keystate_n16, key3FF_keystate_n15, key3FF_keystate_n14,
         key3FF_keystate_n13, key3FF_keystate_n12, key3FF_keystate_n11,
         key3FF_keystate_n10, key3FF_keystate_gff_1_SFF_0_n12,
         key3FF_keystate_gff_1_SFF_0_n11, key3FF_keystate_gff_1_SFF_0_n10,
         key3FF_keystate_gff_1_SFF_0_n8, key3FF_keystate_gff_1_SFF_0_n7,
         key3FF_keystate_gff_1_SFF_1_n12, key3FF_keystate_gff_1_SFF_1_n11,
         key3FF_keystate_gff_1_SFF_1_n10, key3FF_keystate_gff_1_SFF_1_n8,
         key3FF_keystate_gff_1_SFF_1_n7, key3FF_keystate_gff_1_SFF_2_n12,
         key3FF_keystate_gff_1_SFF_2_n11, key3FF_keystate_gff_1_SFF_2_n10,
         key3FF_keystate_gff_1_SFF_2_n8, key3FF_keystate_gff_1_SFF_2_n7,
         key3FF_keystate_gff_1_SFF_3_n12, key3FF_keystate_gff_1_SFF_3_n11,
         key3FF_keystate_gff_1_SFF_3_n10, key3FF_keystate_gff_1_SFF_3_n8,
         key3FF_keystate_gff_1_SFF_3_n7, key3FF_keystate_gff_2_SFF_0_n12,
         key3FF_keystate_gff_2_SFF_0_n11, key3FF_keystate_gff_2_SFF_0_n10,
         key3FF_keystate_gff_2_SFF_0_n8, key3FF_keystate_gff_2_SFF_0_n7,
         key3FF_keystate_gff_2_SFF_1_n12, key3FF_keystate_gff_2_SFF_1_n11,
         key3FF_keystate_gff_2_SFF_1_n10, key3FF_keystate_gff_2_SFF_1_n8,
         key3FF_keystate_gff_2_SFF_1_n7, key3FF_keystate_gff_2_SFF_2_n12,
         key3FF_keystate_gff_2_SFF_2_n11, key3FF_keystate_gff_2_SFF_2_n10,
         key3FF_keystate_gff_2_SFF_2_n8, key3FF_keystate_gff_2_SFF_2_n7,
         key3FF_keystate_gff_2_SFF_3_n12, key3FF_keystate_gff_2_SFF_3_n11,
         key3FF_keystate_gff_2_SFF_3_n10, key3FF_keystate_gff_2_SFF_3_n8,
         key3FF_keystate_gff_2_SFF_3_n7, key3FF_keystate_gff_3_SFF_0_n12,
         key3FF_keystate_gff_3_SFF_0_n11, key3FF_keystate_gff_3_SFF_0_n10,
         key3FF_keystate_gff_3_SFF_0_n8, key3FF_keystate_gff_3_SFF_0_n7,
         key3FF_keystate_gff_3_SFF_1_n12, key3FF_keystate_gff_3_SFF_1_n11,
         key3FF_keystate_gff_3_SFF_1_n10, key3FF_keystate_gff_3_SFF_1_n8,
         key3FF_keystate_gff_3_SFF_1_n7, key3FF_keystate_gff_3_SFF_2_n11,
         key3FF_keystate_gff_3_SFF_2_n10, key3FF_keystate_gff_3_SFF_2_n9,
         key3FF_keystate_gff_3_SFF_2_n7, key3FF_keystate_gff_3_SFF_2_n6,
         key3FF_keystate_gff_3_SFF_3_n11, key3FF_keystate_gff_3_SFF_3_n10,
         key3FF_keystate_gff_3_SFF_3_n9, key3FF_keystate_gff_3_SFF_3_n7,
         key3FF_keystate_gff_3_SFF_3_n6, key3FF_keystate_gff_4_SFF_0_n11,
         key3FF_keystate_gff_4_SFF_0_n10, key3FF_keystate_gff_4_SFF_0_n9,
         key3FF_keystate_gff_4_SFF_0_n7, key3FF_keystate_gff_4_SFF_0_n6,
         key3FF_keystate_gff_4_SFF_1_n11, key3FF_keystate_gff_4_SFF_1_n10,
         key3FF_keystate_gff_4_SFF_1_n9, key3FF_keystate_gff_4_SFF_1_n7,
         key3FF_keystate_gff_4_SFF_1_n6, key3FF_keystate_gff_4_SFF_2_n11,
         key3FF_keystate_gff_4_SFF_2_n10, key3FF_keystate_gff_4_SFF_2_n9,
         key3FF_keystate_gff_4_SFF_2_n7, key3FF_keystate_gff_4_SFF_2_n6,
         key3FF_keystate_gff_4_SFF_3_n11, key3FF_keystate_gff_4_SFF_3_n10,
         key3FF_keystate_gff_4_SFF_3_n9, key3FF_keystate_gff_4_SFF_3_n7,
         key3FF_keystate_gff_4_SFF_3_n6, key3FF_keystate_gff_5_SFF_0_n12,
         key3FF_keystate_gff_5_SFF_0_n11, key3FF_keystate_gff_5_SFF_0_n10,
         key3FF_keystate_gff_5_SFF_0_n8, key3FF_keystate_gff_5_SFF_0_n7,
         key3FF_keystate_gff_5_SFF_1_n12, key3FF_keystate_gff_5_SFF_1_n11,
         key3FF_keystate_gff_5_SFF_1_n10, key3FF_keystate_gff_5_SFF_1_n8,
         key3FF_keystate_gff_5_SFF_1_n7, key3FF_keystate_gff_5_SFF_2_n11,
         key3FF_keystate_gff_5_SFF_2_n10, key3FF_keystate_gff_5_SFF_2_n8,
         key3FF_keystate_gff_5_SFF_2_n7, key3FF_keystate_gff_5_SFF_3_n11,
         key3FF_keystate_gff_5_SFF_3_n10, key3FF_keystate_gff_5_SFF_3_n8,
         key3FF_keystate_gff_5_SFF_3_n7, key3FF_keystate_gff_6_SFF_0_n11,
         key3FF_keystate_gff_6_SFF_0_n10, key3FF_keystate_gff_6_SFF_0_n8,
         key3FF_keystate_gff_6_SFF_0_n7, key3FF_keystate_gff_6_SFF_1_n11,
         key3FF_keystate_gff_6_SFF_1_n10, key3FF_keystate_gff_6_SFF_1_n8,
         key3FF_keystate_gff_6_SFF_1_n7, key3FF_keystate_gff_6_SFF_2_n11,
         key3FF_keystate_gff_6_SFF_2_n10, key3FF_keystate_gff_6_SFF_2_n8,
         key3FF_keystate_gff_6_SFF_2_n7, key3FF_keystate_gff_6_SFF_3_n11,
         key3FF_keystate_gff_6_SFF_3_n10, key3FF_keystate_gff_6_SFF_3_n8,
         key3FF_keystate_gff_6_SFF_3_n7, key3FF_keystate_gff_7_SFF_0_n12,
         key3FF_keystate_gff_7_SFF_0_n11, key3FF_keystate_gff_7_SFF_0_n10,
         key3FF_keystate_gff_7_SFF_0_n8, key3FF_keystate_gff_7_SFF_0_n7,
         key3FF_keystate_gff_7_SFF_1_n12, key3FF_keystate_gff_7_SFF_1_n11,
         key3FF_keystate_gff_7_SFF_1_n10, key3FF_keystate_gff_7_SFF_1_n8,
         key3FF_keystate_gff_7_SFF_1_n7, key3FF_keystate_gff_7_SFF_2_n11,
         key3FF_keystate_gff_7_SFF_2_n10, key3FF_keystate_gff_7_SFF_2_n9,
         key3FF_keystate_gff_7_SFF_2_n7, key3FF_keystate_gff_7_SFF_2_n6,
         key3FF_keystate_gff_7_SFF_3_n11, key3FF_keystate_gff_7_SFF_3_n10,
         key3FF_keystate_gff_7_SFF_3_n9, key3FF_keystate_gff_7_SFF_3_n7,
         key3FF_keystate_gff_7_SFF_3_n6, key3FF_keystate_gff_8_SFF_0_n11,
         key3FF_keystate_gff_8_SFF_0_n10, key3FF_keystate_gff_8_SFF_0_n9,
         key3FF_keystate_gff_8_SFF_0_n7, key3FF_keystate_gff_8_SFF_0_n6,
         key3FF_keystate_gff_8_SFF_1_n11, key3FF_keystate_gff_8_SFF_1_n10,
         key3FF_keystate_gff_8_SFF_1_n9, key3FF_keystate_gff_8_SFF_1_n7,
         key3FF_keystate_gff_8_SFF_1_n6, key3FF_keystate_gff_8_SFF_2_n11,
         key3FF_keystate_gff_8_SFF_2_n10, key3FF_keystate_gff_8_SFF_2_n9,
         key3FF_keystate_gff_8_SFF_2_n7, key3FF_keystate_gff_8_SFF_2_n6,
         key3FF_keystate_gff_8_SFF_3_n11, key3FF_keystate_gff_8_SFF_3_n10,
         key3FF_keystate_gff_8_SFF_3_n9, key3FF_keystate_gff_8_SFF_3_n7,
         key3FF_keystate_gff_8_SFF_3_n6, key3FF_keystate_gff_9_SFF_0_n12,
         key3FF_keystate_gff_9_SFF_0_n11, key3FF_keystate_gff_9_SFF_0_n10,
         key3FF_keystate_gff_9_SFF_0_n8, key3FF_keystate_gff_9_SFF_0_n7,
         key3FF_keystate_gff_9_SFF_1_n12, key3FF_keystate_gff_9_SFF_1_n11,
         key3FF_keystate_gff_9_SFF_1_n10, key3FF_keystate_gff_9_SFF_1_n8,
         key3FF_keystate_gff_9_SFF_1_n7, key3FF_keystate_gff_9_SFF_2_n12,
         key3FF_keystate_gff_9_SFF_2_n11, key3FF_keystate_gff_9_SFF_2_n10,
         key3FF_keystate_gff_9_SFF_2_n8, key3FF_keystate_gff_9_SFF_2_n7,
         key3FF_keystate_gff_9_SFF_3_n12, key3FF_keystate_gff_9_SFF_3_n11,
         key3FF_keystate_gff_9_SFF_3_n10, key3FF_keystate_gff_9_SFF_3_n8,
         key3FF_keystate_gff_9_SFF_3_n7, key3FF_keystate_gff_10_SFF_0_n12,
         key3FF_keystate_gff_10_SFF_0_n11, key3FF_keystate_gff_10_SFF_0_n10,
         key3FF_keystate_gff_10_SFF_0_n8, key3FF_keystate_gff_10_SFF_0_n7,
         key3FF_keystate_gff_10_SFF_1_n12, key3FF_keystate_gff_10_SFF_1_n11,
         key3FF_keystate_gff_10_SFF_1_n10, key3FF_keystate_gff_10_SFF_1_n8,
         key3FF_keystate_gff_10_SFF_1_n7, key3FF_keystate_gff_10_SFF_2_n12,
         key3FF_keystate_gff_10_SFF_2_n11, key3FF_keystate_gff_10_SFF_2_n10,
         key3FF_keystate_gff_10_SFF_2_n8, key3FF_keystate_gff_10_SFF_2_n7,
         key3FF_keystate_gff_10_SFF_3_n12, key3FF_keystate_gff_10_SFF_3_n11,
         key3FF_keystate_gff_10_SFF_3_n10, key3FF_keystate_gff_10_SFF_3_n8,
         key3FF_keystate_gff_10_SFF_3_n7, key3FF_keystate_gff_11_SFF_0_n11,
         key3FF_keystate_gff_11_SFF_0_n10, key3FF_keystate_gff_11_SFF_0_n8,
         key3FF_keystate_gff_11_SFF_0_n7, key3FF_keystate_gff_11_SFF_1_n11,
         key3FF_keystate_gff_11_SFF_1_n10, key3FF_keystate_gff_11_SFF_1_n8,
         key3FF_keystate_gff_11_SFF_1_n7, key3FF_keystate_gff_11_SFF_2_n11,
         key3FF_keystate_gff_11_SFF_2_n10, key3FF_keystate_gff_11_SFF_2_n9,
         key3FF_keystate_gff_11_SFF_2_n7, key3FF_keystate_gff_11_SFF_2_n6,
         key3FF_keystate_gff_11_SFF_3_n11, key3FF_keystate_gff_11_SFF_3_n10,
         key3FF_keystate_gff_11_SFF_3_n9, key3FF_keystate_gff_11_SFF_3_n7,
         key3FF_keystate_gff_11_SFF_3_n6, key3FF_keystate_gff_12_SFF_0_n11,
         key3FF_keystate_gff_12_SFF_0_n10, key3FF_keystate_gff_12_SFF_0_n9,
         key3FF_keystate_gff_12_SFF_0_n7, key3FF_keystate_gff_12_SFF_0_n6,
         key3FF_keystate_gff_12_SFF_1_n11, key3FF_keystate_gff_12_SFF_1_n10,
         key3FF_keystate_gff_12_SFF_1_n9, key3FF_keystate_gff_12_SFF_1_n7,
         key3FF_keystate_gff_12_SFF_1_n6, key3FF_keystate_gff_12_SFF_2_n11,
         key3FF_keystate_gff_12_SFF_2_n10, key3FF_keystate_gff_12_SFF_2_n9,
         key3FF_keystate_gff_12_SFF_2_n7, key3FF_keystate_gff_12_SFF_2_n6,
         key3FF_keystate_gff_12_SFF_3_n11, key3FF_keystate_gff_12_SFF_3_n10,
         key3FF_keystate_gff_12_SFF_3_n9, key3FF_keystate_gff_12_SFF_3_n7,
         key3FF_keystate_gff_12_SFF_3_n6, key3FF_keystate_gff_13_SFF_0_n12,
         key3FF_keystate_gff_13_SFF_0_n11, key3FF_keystate_gff_13_SFF_0_n10,
         key3FF_keystate_gff_13_SFF_0_n8, key3FF_keystate_gff_13_SFF_0_n7,
         key3FF_keystate_gff_13_SFF_1_n12, key3FF_keystate_gff_13_SFF_1_n11,
         key3FF_keystate_gff_13_SFF_1_n10, key3FF_keystate_gff_13_SFF_1_n8,
         key3FF_keystate_gff_13_SFF_1_n7, key3FF_keystate_gff_13_SFF_2_n11,
         key3FF_keystate_gff_13_SFF_2_n10, key3FF_keystate_gff_13_SFF_2_n8,
         key3FF_keystate_gff_13_SFF_2_n7, key3FF_keystate_gff_13_SFF_3_n11,
         key3FF_keystate_gff_13_SFF_3_n10, key3FF_keystate_gff_13_SFF_3_n8,
         key3FF_keystate_gff_13_SFF_3_n7, key3FF_keystate_gff_14_SFF_0_n11,
         key3FF_keystate_gff_14_SFF_0_n10, key3FF_keystate_gff_14_SFF_0_n8,
         key3FF_keystate_gff_14_SFF_0_n7, key3FF_keystate_gff_14_SFF_1_n11,
         key3FF_keystate_gff_14_SFF_1_n10, key3FF_keystate_gff_14_SFF_1_n8,
         key3FF_keystate_gff_14_SFF_1_n7, key3FF_keystate_gff_14_SFF_2_n11,
         key3FF_keystate_gff_14_SFF_2_n10, key3FF_keystate_gff_14_SFF_2_n8,
         key3FF_keystate_gff_14_SFF_2_n7, key3FF_keystate_gff_14_SFF_3_n11,
         key3FF_keystate_gff_14_SFF_3_n10, key3FF_keystate_gff_14_SFF_3_n8,
         key3FF_keystate_gff_14_SFF_3_n7, key3FF_keystate_gff_15_SFF_0_n11,
         key3FF_keystate_gff_15_SFF_0_n10, key3FF_keystate_gff_15_SFF_0_n8,
         key3FF_keystate_gff_15_SFF_0_n7, key3FF_keystate_gff_15_SFF_1_n11,
         key3FF_keystate_gff_15_SFF_1_n10, key3FF_keystate_gff_15_SFF_1_n8,
         key3FF_keystate_gff_15_SFF_1_n7, key3FF_keystate_gff_15_SFF_2_n11,
         key3FF_keystate_gff_15_SFF_2_n10, key3FF_keystate_gff_15_SFF_2_n9,
         key3FF_keystate_gff_15_SFF_2_n7, key3FF_keystate_gff_15_SFF_2_n6,
         key3FF_keystate_gff_15_SFF_3_n11, key3FF_keystate_gff_15_SFF_3_n10,
         key3FF_keystate_gff_15_SFF_3_n9, key3FF_keystate_gff_15_SFF_3_n7,
         key3FF_keystate_gff_15_SFF_3_n6, key3FF_keystate_gff_16_SFF_0_n11,
         key3FF_keystate_gff_16_SFF_0_n10, key3FF_keystate_gff_16_SFF_0_n9,
         key3FF_keystate_gff_16_SFF_0_n7, key3FF_keystate_gff_16_SFF_0_n6,
         key3FF_keystate_gff_16_SFF_1_n11, key3FF_keystate_gff_16_SFF_1_n10,
         key3FF_keystate_gff_16_SFF_1_n9, key3FF_keystate_gff_16_SFF_1_n7,
         key3FF_keystate_gff_16_SFF_1_n6, key3FF_keystate_gff_16_SFF_2_n10,
         key3FF_keystate_gff_16_SFF_2_n9, key3FF_keystate_gff_16_SFF_2_n7,
         key3FF_keystate_gff_16_SFF_2_n6, key3FF_keystate_gff_16_SFF_3_n10,
         key3FF_keystate_gff_16_SFF_3_n9, key3FF_keystate_gff_16_SFF_3_n7,
         key3FF_keystate_gff_16_SFF_3_n6, key3FF_keystate_gff_17_SFF_0_n12,
         key3FF_keystate_gff_17_SFF_0_n11, key3FF_keystate_gff_17_SFF_0_n10,
         key3FF_keystate_gff_17_SFF_0_n8, key3FF_keystate_gff_17_SFF_0_n7,
         key3FF_keystate_gff_17_SFF_1_n12, key3FF_keystate_gff_17_SFF_1_n11,
         key3FF_keystate_gff_17_SFF_1_n10, key3FF_keystate_gff_17_SFF_1_n8,
         key3FF_keystate_gff_17_SFF_1_n7, key3FF_keystate_gff_17_SFF_2_n11,
         key3FF_keystate_gff_17_SFF_2_n10, key3FF_keystate_gff_17_SFF_2_n8,
         key3FF_keystate_gff_17_SFF_2_n7, key3FF_keystate_gff_17_SFF_3_n11,
         key3FF_keystate_gff_17_SFF_3_n10, key3FF_keystate_gff_17_SFF_3_n8,
         key3FF_keystate_gff_17_SFF_3_n7, key3FF_keystate_gff_18_SFF_0_n11,
         key3FF_keystate_gff_18_SFF_0_n10, key3FF_keystate_gff_18_SFF_0_n8,
         key3FF_keystate_gff_18_SFF_0_n7, key3FF_keystate_gff_18_SFF_1_n11,
         key3FF_keystate_gff_18_SFF_1_n10, key3FF_keystate_gff_18_SFF_1_n8,
         key3FF_keystate_gff_18_SFF_1_n7, key3FF_keystate_gff_18_SFF_2_n11,
         key3FF_keystate_gff_18_SFF_2_n10, key3FF_keystate_gff_18_SFF_2_n8,
         key3FF_keystate_gff_18_SFF_2_n7, key3FF_keystate_gff_18_SFF_3_n11,
         key3FF_keystate_gff_18_SFF_3_n10, key3FF_keystate_gff_18_SFF_3_n8,
         key3FF_keystate_gff_18_SFF_3_n7, key3FF_keystate_gff_19_SFF_0_n11,
         key3FF_keystate_gff_19_SFF_0_n10, key3FF_keystate_gff_19_SFF_0_n8,
         key3FF_keystate_gff_19_SFF_0_n7, key3FF_keystate_gff_19_SFF_1_n11,
         key3FF_keystate_gff_19_SFF_1_n10, key3FF_keystate_gff_19_SFF_1_n8,
         key3FF_keystate_gff_19_SFF_1_n7, key3FF_keystate_gff_19_SFF_2_n11,
         key3FF_keystate_gff_19_SFF_2_n10, key3FF_keystate_gff_19_SFF_2_n9,
         key3FF_keystate_gff_19_SFF_2_n7, key3FF_keystate_gff_19_SFF_2_n6,
         key3FF_keystate_gff_19_SFF_3_n11, key3FF_keystate_gff_19_SFF_3_n10,
         key3FF_keystate_gff_19_SFF_3_n9, key3FF_keystate_gff_19_SFF_3_n7,
         key3FF_keystate_gff_19_SFF_3_n6, key3FF_keystate_gff_20_SFF_0_n10,
         key3FF_keystate_gff_20_SFF_0_n9, key3FF_keystate_gff_20_SFF_0_n7,
         key3FF_keystate_gff_20_SFF_0_n6, key3FF_keystate_gff_20_SFF_1_n10,
         key3FF_keystate_gff_20_SFF_1_n9, key3FF_keystate_gff_20_SFF_1_n7,
         key3FF_keystate_gff_20_SFF_1_n6, key3FF_keystate_gff_20_SFF_2_n10,
         key3FF_keystate_gff_20_SFF_2_n9, key3FF_keystate_gff_20_SFF_2_n7,
         key3FF_keystate_gff_20_SFF_2_n6, key3FF_keystate_gff_20_SFF_3_n10,
         key3FF_keystate_gff_20_SFF_3_n9, key3FF_keystate_gff_20_SFF_3_n7,
         key3FF_keystate_gff_20_SFF_3_n6, sbox_F_in3_3_, sbox_F_in2_3_,
         sbox_F_in1_3_, sbox_F_n4, sbox_F_n3, sbox_F_n2, sbox_F_n1,
         sbox_F_Inst_1__CF_Inst_n1, sbox_F_Inst_3__CF_Inst_n1,
         sbox_F_Inst_4__CF_Inst_n2, sbox_F_Inst_5__CF_Inst_n2,
         sbox_F_Inst_6__CF_Inst_n2, sbox_F_Inst_7__CF_Inst_n2,
         sbox_F_Inst_8__CF_Inst_n2, sbox_F_Inst_8__CF_Inst_n1,
         sbox_F_Inst_9__CF_Inst_n2, sbox_F_Inst_10__CF_Inst_n2,
         sbox_F_Inst_10__CF_Inst_n1, sbox_F_Inst_11__CF_Inst_n2,
         sbox_F_Inst_12__CF_Inst_n2, sbox_F_Inst_12__CF_Inst_n1,
         sbox_F_Inst_13__CF_Inst_n2, sbox_F_Inst_14__CF_Inst_n2,
         sbox_F_Inst_15__CF_Inst_n2, sbox_F_Inst_16__CF_Inst_n2,
         sbox_F_Inst_17__CF_Inst_n2, sbox_F_Inst_18__CF_Inst_n1,
         sbox_F_Inst_19__CF_Inst_n2, sbox_F_Inst_19__CF_Inst_n1,
         sbox_F_Inst_20__CF_Inst_n2, sbox_F_Inst_20__CF_Inst_n1,
         sbox_F_Inst_22__CF_Inst_n1, sbox_F_Inst_23__CF_Inst_n1,
         sbox_F_Inst_24__CF_Inst_n1, sbox_F_Inst_26__CF_Inst_n1,
         sbox_F_Inst_27__CF_Inst_n3, sbox_F_Inst_27__CF_Inst_n2,
         sbox_F_Inst_28__CF_Inst_n2, sbox_F_Inst_28__CF_Inst_n1,
         sbox_F_Inst_29__CF_Inst_n2, sbox_F_Inst_29__CF_Inst_n1,
         sbox_F_Inst_30__CF_Inst_n2, sbox_F_Inst_30__CF_Inst_n1,
         sbox_F_Inst_31__CF_Inst_n1, sbox_F_Inst_32__CF_Inst_n1,
         sbox_F_Inst_33__CF_Inst_n5, sbox_F_Inst_33__CF_Inst_n4,
         sbox_F_Inst_33__CF_Inst_n3, sbox_F_Inst_35__CF_Inst_n2,
         sbox_F_Inst_35__CF_Inst_n1, sbox_F_InstXOR_0__Compression1_n3,
         sbox_F_InstXOR_0__Compression2_n3, sbox_F_InstXOR_0__Compression3_n3,
         sbox_F_InstXOR_1__Compression1_n3, sbox_F_InstXOR_1__Compression2_n3,
         sbox_F_InstXOR_1__Compression3_n3, sbox_F_InstXOR_2__Compression1_n3,
         sbox_F_InstXOR_2__Compression2_n3, sbox_F_InstXOR_2__Compression3_n3,
         sbox_F_InstXOR_3__Compression1_n3, sbox_F_InstXOR_3__Compression2_n3,
         sbox_F_InstXOR_3__Compression3_n3, sbox_G_n1, sbox_G_N3, sbox_G_N2,
         sbox_G_Inst_1__CF_Inst_n2, sbox_G_Inst_2__CF_Inst_n2,
         sbox_G_Inst_2__CF_Inst_n1, sbox_G_Inst_3__CF_Inst_n2,
         sbox_G_Inst_5__CF_Inst_n2, sbox_G_Inst_5__CF_Inst_n1,
         sbox_G_Inst_6__CF_Inst_n1, sbox_G_Inst_8__CF_Inst_n2,
         sbox_G_Inst_9__CF_Inst_n2, sbox_G_Inst_9__CF_Inst_n1,
         sbox_G_Inst_11__CF_Inst_n2, sbox_G_Inst_11__CF_Inst_n1,
         sbox_G_Inst_12__CF_Inst_n2, sbox_G_Inst_12__CF_Inst_n1,
         sbox_G_Inst_14__CF_Inst_n1, sbox_G_Inst_15__CF_Inst_n2,
         sbox_G_Inst_15__CF_Inst_n1, sbox_G_Inst_17__CF_Inst_n2,
         sbox_G_Inst_18__CF_Inst_n2, sbox_G_Inst_19__CF_Inst_n2,
         sbox_G_Inst_20__CF_Inst_n2, sbox_G_Inst_20__CF_Inst_n1,
         sbox_G_Inst_23__CF_Inst_n2, sbox_G_Inst_23__CF_Inst_n1,
         sbox_G_Inst_24__CF_Inst_n1, sbox_G_InstXOR_0__Compression1_n3,
         sbox_G_InstXOR_0__Compression2_n3, sbox_G_InstXOR_0__Compression3_n3,
         sbox_G_InstXOR_1__Compression1_n3, sbox_G_InstXOR_1__Compression2_n3,
         sbox_G_InstXOR_1__Compression3_n3, sbox_G_InstXOR_2__Compression1_n3,
         sbox_G_InstXOR_2__Compression2_n3, sbox_G_InstXOR_2__Compression3_n3;
  wire   [4:0] counter;
  wire   [3:0] sboxOut1;
  wire   [3:0] sboxOut2;
  wire   [3:0] sboxOut3;
  wire   [3:0] roundkey1;
  wire   [3:1] keyRegKS1;
  wire   [3:0] roundkey2;
  wire   [3:1] keyRegKS2;
  wire   [3:0] roundkey3;
  wire   [3:1] keyRegKS3;
  wire   [3:0] AddKeyOut1;
  wire   [3:0] AddKeyOut2;
  wire   [3:0] AddKeyOut3;
  wire   [63:0] state1FF_inputPar;
  wire   [63:0] state2FF_inputPar;
  wire   [63:0] state3FF_inputPar;
  wire   [4:0] key1FF_counterAdd;
  wire   [75:3] key1FF_outputPar;
  wire   [4:0] key2FF_counterAdd;
  wire   [75:3] key2FF_outputPar;
  wire   [4:0] key3FF_counterAdd;
  wire   [75:3] key3FF_outputPar;
  wire   [3:0] sbox_F_in3_reg;
  wire   [3:0] sbox_F_in2_reg;
  wire   [3:0] sbox_F_in1_reg;
  wire   [3:0] sbox_q3;
  wire   [3:0] sbox_Rq3;
  wire   [3:0] sbox_q2;
  wire   [3:0] sbox_Rq2;
  wire   [3:0] sbox_q1;
  wire   [3:0] sbox_Rq1;
  wire   [3:0] sbox_F_q3;
  wire   [3:0] sbox_F_q2;
  wire   [3:0] sbox_F_q1;
  wire   [35:0] sbox_F_CF_Reg;
  wire   [35:0] sbox_F_CF_Out;
  wire   [26:0] sbox_G_CF_Reg;
  wire   [26:0] sbox_G_CF_Out;

  BUF_X2 U26 ( .A(selInit), .Z(n4) );
  XOR2_X1 U27 ( .A(state1FF_inputPar[15]), .B(roundkey1[0]), .Z(AddKeyOut1[0])
         );
  XOR2_X1 U28 ( .A(state1FF_inputPar[31]), .B(roundkey1[1]), .Z(AddKeyOut1[1])
         );
  XOR2_X1 U29 ( .A(state1FF_inputPar[47]), .B(roundkey1[2]), .Z(AddKeyOut1[2])
         );
  XOR2_X1 U30 ( .A(state1FF_inputPar[63]), .B(roundkey1[3]), .Z(AddKeyOut1[3])
         );
  XOR2_X1 U31 ( .A(state2FF_inputPar[15]), .B(roundkey2[0]), .Z(AddKeyOut2[0])
         );
  XOR2_X1 U32 ( .A(state2FF_inputPar[31]), .B(roundkey2[1]), .Z(AddKeyOut2[1])
         );
  XOR2_X1 U33 ( .A(state2FF_inputPar[47]), .B(roundkey2[2]), .Z(AddKeyOut2[2])
         );
  XOR2_X1 U34 ( .A(state2FF_inputPar[63]), .B(roundkey2[3]), .Z(AddKeyOut2[3])
         );
  XOR2_X1 U35 ( .A(state3FF_inputPar[15]), .B(roundkey3[0]), .Z(AddKeyOut3[0])
         );
  XOR2_X1 U36 ( .A(state3FF_inputPar[31]), .B(roundkey3[1]), .Z(AddKeyOut3[1])
         );
  XOR2_X1 U37 ( .A(state3FF_inputPar[47]), .B(roundkey3[2]), .Z(AddKeyOut3[2])
         );
  XOR2_X1 U38 ( .A(state3FF_inputPar[63]), .B(roundkey3[3]), .Z(AddKeyOut3[3])
         );
  NAND2_X1 fsm_U33 ( .A1(fsm_en_countSerial), .A2(fsm_n31), .ZN(selSbox) );
  OAI21_X1 fsm_U32 ( .B1(fsm_n30), .B2(fsm_n29), .A(fsm_n28), .ZN(fsm_n23) );
  AOI21_X1 fsm_U31 ( .B1(fsm_n27), .B2(fsm_n26), .A(fsm_n25), .ZN(fsm_n30) );
  AOI221_X1 fsm_U30 ( .B1(fsm_n24), .B2(fsm_n20), .C1(fsm_n19), .C2(fsm_n20), 
        .A(fsm_n29), .ZN(fsm_n22) );
  OR3_X1 fsm_U29 ( .A1(enData), .A2(fsm_ps_state_0_), .A3(fsm_ps_state_1_), 
        .ZN(fsm_n20) );
  OAI21_X1 fsm_U28 ( .B1(fsm_n18), .B2(fsm_n29), .A(fsm_n28), .ZN(fsm_n21) );
  NAND3_X1 fsm_U27 ( .A1(nReset), .A2(done), .A3(fsm_n19), .ZN(fsm_n28) );
  NAND4_X1 fsm_U26 ( .A1(fsm_n17), .A2(fsm_countSerial_3_), .A3(
        fsm_countSerial_2_), .A4(fsm_n16), .ZN(fsm_n19) );
  AND2_X1 fsm_U25 ( .A1(fsm_countSerial_0_), .A2(fsm_countSerial_1_), .ZN(
        fsm_n17) );
  AOI21_X1 fsm_U24 ( .B1(fsm_n15), .B2(counter[2]), .A(fsm_en_countRound), 
        .ZN(fsm_n18) );
  NOR2_X1 fsm_U23 ( .A1(fsm_n14), .A2(fsm_n13), .ZN(fsm_n15) );
  NAND4_X1 fsm_U22 ( .A1(counter[1]), .A2(counter[3]), .A3(counter[0]), .A4(
        counter[4]), .ZN(fsm_n13) );
  NOR2_X1 fsm_U21 ( .A1(fsm_n12), .A2(fsm_n26), .ZN(fsm_en_countRound) );
  NAND4_X1 fsm_U20 ( .A1(fsm_countSerial_4_), .A2(fsm_countSerial_0_), .A3(
        fsm_countSerial_1_), .A4(fsm_n11), .ZN(fsm_n26) );
  NOR2_X1 fsm_U19 ( .A1(fsm_countSerial_3_), .A2(fsm_countSerial_2_), .ZN(
        fsm_n11) );
  INV_X1 fsm_U18 ( .A(fsm_n27), .ZN(fsm_n12) );
  NOR2_X1 fsm_U17 ( .A1(fsm_n10), .A2(fsm_ps_state_1_), .ZN(fsm_n27) );
  INV_X1 fsm_U16 ( .A(fsm_n24), .ZN(done) );
  NAND2_X1 fsm_U15 ( .A1(fsm_en_countSerial), .A2(fsm_ps_state_1_), .ZN(
        fsm_n24) );
  NOR2_X1 fsm_U14 ( .A1(fsm_rst_countSerial), .A2(fsm_ps_state_1_), .ZN(
        selInit) );
  INV_X1 fsm_U13 ( .A(selInit), .ZN(fsm_n9) );
  NAND2_X1 fsm_U12 ( .A1(enData), .A2(fsm_ps_state_0_), .ZN(fsm_n10) );
  INV_X1 fsm_U11 ( .A(fsm_countSerial_4_), .ZN(fsm_n16) );
  INV_X1 fsm_U10 ( .A(fsm_n10), .ZN(fsm_en_countSerial) );
  OAI21_X1 fsm_U9 ( .B1(fsm_ps_state_1_), .B2(fsm_n16), .A(fsm_en_countSerial), 
        .ZN(fsm_n31) );
  NOR2_X1 fsm_U8 ( .A1(fsm_ps_state_2_), .A2(fsm_ps_state_0_), .ZN(fsm_n25) );
  INV_X1 fsm_U7 ( .A(fsm_n25), .ZN(fsm_rst_countSerial) );
  NAND2_X1 fsm_U6 ( .A1(fsm_n31), .A2(fsm_rst_countSerial), .ZN(enKey) );
  NAND2_X1 fsm_U5 ( .A1(fsm_ps_state_1_), .A2(fsm_n25), .ZN(fsm_n14) );
  INV_X1 fsm_U4 ( .A(nReset), .ZN(fsm_n29) );
  INV_X1 fsm_U3 ( .A(fsm_n14), .ZN(selP) );
  DFF_X1 fsm_ps_state_reg_2_ ( .D(fsm_n22), .CK(clk), .Q(fsm_ps_state_2_), 
        .QN(enData) );
  DFF_X1 fsm_ps_state_reg_1_ ( .D(fsm_n21), .CK(clk), .Q(fsm_ps_state_1_), 
        .QN() );
  DFF_X1 fsm_ps_state_reg_0_ ( .D(fsm_n23), .CK(clk), .Q(fsm_ps_state_0_), 
        .QN() );
  OAI22_X1 fsm_cnt_rnd_U18 ( .A1(fsm_cnt_rnd_n25), .A2(fsm_cnt_rnd_n38), .B1(
        fsm_cnt_rnd_n20), .B2(fsm_cnt_rnd_n37), .ZN(fsm_cnt_rnd_n2) );
  OR2_X1 fsm_cnt_rnd_U17 ( .A1(fsm_cnt_rnd_n36), .A2(counter[1]), .ZN(
        fsm_cnt_rnd_n37) );
  AOI21_X1 fsm_cnt_rnd_U16 ( .B1(fsm_cnt_rnd_n35), .B2(fsm_cnt_rnd_n20), .A(
        fsm_cnt_rnd_n38), .ZN(fsm_cnt_rnd_n19) );
  OAI22_X1 fsm_cnt_rnd_U15 ( .A1(fsm_cnt_rnd_n26), .A2(fsm_cnt_rnd_n33), .B1(
        fsm_cnt_rnd_n32), .B2(counter[2]), .ZN(fsm_cnt_rnd_n34) );
  OAI21_X1 fsm_cnt_rnd_U14 ( .B1(fsm_cnt_rnd_n36), .B2(counter[1]), .A(
        fsm_cnt_rnd_n38), .ZN(fsm_cnt_rnd_n33) );
  OAI21_X1 fsm_cnt_rnd_U13 ( .B1(fsm_cnt_rnd_n35), .B2(fsm_cnt_rnd_n20), .A(
        fsm_n9), .ZN(fsm_cnt_rnd_n38) );
  INV_X1 fsm_cnt_rnd_U12 ( .A(fsm_en_countRound), .ZN(fsm_cnt_rnd_n35) );
  AOI22_X1 fsm_cnt_rnd_U11 ( .A1(counter[3]), .A2(fsm_cnt_rnd_n31), .B1(
        fsm_cnt_rnd_n30), .B2(fsm_cnt_rnd_n24), .ZN(fsm_cnt_rnd_n21) );
  NAND2_X1 fsm_cnt_rnd_U10 ( .A1(counter[2]), .A2(fsm_cnt_rnd_n32), .ZN(
        fsm_cnt_rnd_n30) );
  NOR3_X1 fsm_cnt_rnd_U9 ( .A1(fsm_cnt_rnd_n25), .A2(fsm_cnt_rnd_n20), .A3(
        fsm_cnt_rnd_n36), .ZN(fsm_cnt_rnd_n32) );
  OAI21_X1 fsm_cnt_rnd_U8 ( .B1(fsm_cnt_rnd_n36), .B2(counter[3]), .A(
        fsm_cnt_rnd_n31), .ZN(fsm_cnt_rnd_n29) );
  NAND2_X1 fsm_cnt_rnd_U7 ( .A1(fsm_n9), .A2(fsm_cnt_rnd_n28), .ZN(
        fsm_cnt_rnd_n31) );
  NAND4_X1 fsm_cnt_rnd_U6 ( .A1(counter[1]), .A2(fsm_en_countRound), .A3(
        counter[0]), .A4(counter[2]), .ZN(fsm_cnt_rnd_n28) );
  NAND2_X1 fsm_cnt_rnd_U5 ( .A1(fsm_n9), .A2(fsm_en_countRound), .ZN(
        fsm_cnt_rnd_n36) );
  MUX2_X1 fsm_cnt_rnd_U4 ( .A(fsm_cnt_rnd_n29), .B(fsm_cnt_rnd_n27), .S(
        fsm_cnt_rnd_n23), .Z(fsm_cnt_rnd_n22) );
  NOR2_X1 fsm_cnt_rnd_U3 ( .A1(fsm_cnt_rnd_n24), .A2(fsm_cnt_rnd_n30), .ZN(
        fsm_cnt_rnd_n27) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_4_ ( .D(fsm_cnt_rnd_n22), .CK(clk), .Q(
        counter[4]), .QN(fsm_cnt_rnd_n23) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_3_ ( .D(fsm_cnt_rnd_n21), .CK(clk), .Q(
        counter[3]), .QN(fsm_cnt_rnd_n24) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_2_ ( .D(fsm_cnt_rnd_n34), .CK(clk), .Q(
        fsm_cnt_rnd_n26), .QN(counter[2]) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_1_ ( .D(fsm_cnt_rnd_n2), .CK(clk), .Q(
        counter[1]), .QN(fsm_cnt_rnd_n25) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_0_ ( .D(fsm_cnt_rnd_n19), .CK(clk), .Q(
        counter[0]), .QN(fsm_cnt_rnd_n20) );
  AOI22_X1 fsm_cnt_ser_U22 ( .A1(fsm_countSerial_0_), .A2(fsm_cnt_ser_n43), 
        .B1(fsm_cnt_ser_n42), .B2(fsm_cnt_ser_n29), .ZN(fsm_cnt_ser_n5) );
  OR2_X1 fsm_cnt_ser_U21 ( .A1(fsm_cnt_ser_n41), .A2(fsm_en_countSerial), .ZN(
        fsm_cnt_ser_n43) );
  OAI21_X1 fsm_cnt_ser_U20 ( .B1(fsm_cnt_ser_n40), .B2(fsm_countSerial_4_), 
        .A(fsm_cnt_ser_n39), .ZN(fsm_cnt_ser_n20) );
  OAI21_X1 fsm_cnt_ser_U19 ( .B1(fsm_cnt_ser_n38), .B2(fsm_cnt_ser_n37), .A(
        fsm_countSerial_4_), .ZN(fsm_cnt_ser_n39) );
  NAND3_X1 fsm_cnt_ser_U18 ( .A1(fsm_cnt_ser_n36), .A2(fsm_countSerial_3_), 
        .A3(fsm_cnt_ser_n35), .ZN(fsm_cnt_ser_n40) );
  AOI22_X1 fsm_cnt_ser_U17 ( .A1(fsm_countSerial_3_), .A2(fsm_cnt_ser_n38), 
        .B1(fsm_cnt_ser_n37), .B2(fsm_cnt_ser_n35), .ZN(fsm_cnt_ser_n34) );
  NOR2_X1 fsm_cnt_ser_U16 ( .A1(fsm_countSerial_3_), .A2(fsm_cnt_ser_n42), 
        .ZN(fsm_cnt_ser_n37) );
  AOI21_X1 fsm_cnt_ser_U15 ( .B1(fsm_en_countSerial), .B2(fsm_cnt_ser_n35), 
        .A(fsm_cnt_ser_n41), .ZN(fsm_cnt_ser_n38) );
  NOR3_X1 fsm_cnt_ser_U14 ( .A1(fsm_cnt_ser_n29), .A2(fsm_cnt_ser_n30), .A3(
        fsm_cnt_ser_n28), .ZN(fsm_cnt_ser_n35) );
  AOI22_X1 fsm_cnt_ser_U13 ( .A1(fsm_countSerial_1_), .A2(fsm_cnt_ser_n31), 
        .B1(fsm_cnt_ser_n33), .B2(fsm_cnt_ser_n28), .ZN(fsm_cnt_ser_n23) );
  NAND2_X1 fsm_cnt_ser_U12 ( .A1(fsm_cnt_ser_n36), .A2(fsm_countSerial_0_), 
        .ZN(fsm_cnt_ser_n33) );
  INV_X1 fsm_cnt_ser_U11 ( .A(fsm_cnt_ser_n42), .ZN(fsm_cnt_ser_n36) );
  NAND2_X1 fsm_cnt_ser_U10 ( .A1(fsm_en_countSerial), .A2(fsm_rst_countSerial), 
        .ZN(fsm_cnt_ser_n42) );
  INV_X1 fsm_cnt_ser_U9 ( .A(fsm_cnt_ser_n32), .ZN(fsm_cnt_ser_n31) );
  AOI21_X1 fsm_cnt_ser_U8 ( .B1(fsm_en_countSerial), .B2(fsm_countSerial_0_), 
        .A(fsm_cnt_ser_n41), .ZN(fsm_cnt_ser_n32) );
  INV_X1 fsm_cnt_ser_U7 ( .A(fsm_rst_countSerial), .ZN(fsm_cnt_ser_n41) );
  INV_X1 fsm_cnt_ser_U5 ( .A(fsm_cnt_ser_n30), .ZN(fsm_cnt_ser_n26) );
  AOI21_X1 fsm_cnt_ser_U4 ( .B1(fsm_cnt_ser_n28), .B2(fsm_cnt_ser_n36), .A(
        fsm_cnt_ser_n32), .ZN(fsm_cnt_ser_n25) );
  OAI33_X1 fsm_cnt_ser_U3 ( .A1(1'b0), .A2(fsm_cnt_ser_n30), .A3(
        fsm_cnt_ser_n25), .B1(fsm_cnt_ser_n26), .B2(fsm_cnt_ser_n28), .B3(
        fsm_cnt_ser_n33), .ZN(fsm_cnt_ser_n22) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_3_ ( .D(fsm_cnt_ser_n34), .CK(clk), .Q(), 
        .QN(fsm_countSerial_3_) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_0_ ( .D(fsm_cnt_ser_n5), .CK(clk), .Q(
        fsm_countSerial_0_), .QN(fsm_cnt_ser_n29) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_1_ ( .D(fsm_cnt_ser_n23), .CK(clk), .Q(
        fsm_countSerial_1_), .QN(fsm_cnt_ser_n28) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_2_ ( .D(fsm_cnt_ser_n22), .CK(clk), .Q(
        fsm_countSerial_2_), .QN(fsm_cnt_ser_n30) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_4_ ( .D(fsm_cnt_ser_n20), .CK(clk), .Q(
        fsm_countSerial_4_), .QN() );
  MUX2_X1 state1FF_U5 ( .A(sboxOut1[0]), .B(dataIn1[0]), .S(n4), .Z(
        state1FF_n1) );
  MUX2_X1 state1FF_U4 ( .A(sboxOut1[2]), .B(dataIn1[2]), .S(n4), .Z(
        state1FF_n2) );
  MUX2_X1 state1FF_U3 ( .A(sboxOut1[1]), .B(dataIn1[1]), .S(n4), .Z(
        state1FF_n3) );
  MUX2_X1 state1FF_U2 ( .A(sboxOut1[3]), .B(dataIn1[3]), .S(n4), .Z(
        state1FF_n4) );
  BUF_X1 state1FF_state_U8 ( .A(selP), .Z(state1FF_state_n11) );
  BUF_X1 state1FF_state_U7 ( .A(selP), .Z(state1FF_state_n10) );
  BUF_X1 state1FF_state_U6 ( .A(selP), .Z(state1FF_state_n13) );
  BUF_X1 state1FF_state_U5 ( .A(selP), .Z(state1FF_state_n12) );
  BUF_X2 state1FF_state_U4 ( .A(enData), .Z(state1FF_state_n6) );
  BUF_X2 state1FF_state_U3 ( .A(enData), .Z(state1FF_state_n9) );
  BUF_X2 state1FF_state_U2 ( .A(enData), .Z(state1FF_state_n8) );
  BUF_X2 state1FF_state_U1 ( .A(enData), .Z(state1FF_state_n7) );
  OAI21_X1 state1FF_state_gff_1_SFF_0_U4 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_1_SFF_0_n7), .A(state1FF_state_gff_1_SFF_0_n10), 
        .ZN(state1FF_state_gff_1_SFF_0_n6) );
  OAI221_X1 state1FF_state_gff_1_SFF_0_U3 ( .B1(state1FF_state_n13), .B2(
        state1FF_n1), .C1(state1FF_state_gff_1_SFF_0_n9), .C2(
        state1FF_inputPar[0]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_1_SFF_0_n10) );
  INV_X1 state1FF_state_gff_1_SFF_0_U2 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_1_SFF_0_n9) );
  DFF_X1 state1FF_state_gff_1_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_1_SFF_0_n6), .CK(clk), .Q(state1FF_inputPar[0]), 
        .QN(state1FF_state_gff_1_SFF_0_n7) );
  OAI21_X1 state1FF_state_gff_1_SFF_1_U4 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_1_SFF_1_n8), .A(state1FF_state_gff_1_SFF_1_n11), 
        .ZN(state1FF_state_gff_1_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_1_SFF_1_U3 ( .B1(state1FF_state_n13), .B2(
        state1FF_n3), .C1(state1FF_state_gff_1_SFF_1_n10), .C2(
        state1FF_inputPar[1]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_1_SFF_1_n11) );
  INV_X1 state1FF_state_gff_1_SFF_1_U2 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_1_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_1_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_1_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[16]), 
        .QN(state1FF_state_gff_1_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_1_SFF_2_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_1_SFF_2_n8), .A(state1FF_state_gff_1_SFF_2_n12), 
        .ZN(state1FF_state_gff_1_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_1_SFF_2_U4 ( .B1(state1FF_state_gff_1_SFF_2_n10), .B2(state1FF_n2), .C1(state1FF_state_gff_1_SFF_2_n11), .C2(
        state1FF_inputPar[2]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_1_SFF_2_n12) );
  INV_X1 state1FF_state_gff_1_SFF_2_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_1_SFF_2_n11) );
  INV_X1 state1FF_state_gff_1_SFF_2_U2 ( .A(state1FF_state_gff_1_SFF_2_n11), 
        .ZN(state1FF_state_gff_1_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_1_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_1_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[32]), 
        .QN(state1FF_state_gff_1_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_1_SFF_3_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_1_SFF_3_n8), .A(state1FF_state_gff_1_SFF_3_n12), 
        .ZN(state1FF_state_gff_1_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_1_SFF_3_U4 ( .B1(state1FF_state_gff_1_SFF_3_n10), .B2(state1FF_n4), .C1(state1FF_state_gff_1_SFF_3_n11), .C2(
        state1FF_inputPar[3]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_1_SFF_3_n12) );
  INV_X1 state1FF_state_gff_1_SFF_3_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_1_SFF_3_n11) );
  INV_X1 state1FF_state_gff_1_SFF_3_U2 ( .A(state1FF_state_gff_1_SFF_3_n11), 
        .ZN(state1FF_state_gff_1_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_1_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_1_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[48]), 
        .QN(state1FF_state_gff_1_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_2_SFF_0_U5 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_2_SFF_0_n8), .A(state1FF_state_gff_2_SFF_0_n12), 
        .ZN(state1FF_state_gff_2_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_2_SFF_0_U4 ( .B1(state1FF_state_gff_2_SFF_0_n10), .B2(state1FF_inputPar[0]), .C1(state1FF_state_gff_2_SFF_0_n11), .C2(
        state1FF_inputPar[4]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_2_SFF_0_n12) );
  INV_X1 state1FF_state_gff_2_SFF_0_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_2_SFF_0_n11) );
  INV_X1 state1FF_state_gff_2_SFF_0_U2 ( .A(state1FF_state_gff_2_SFF_0_n11), 
        .ZN(state1FF_state_gff_2_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_2_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_2_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[1]), 
        .QN(state1FF_state_gff_2_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_2_SFF_1_U5 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_2_SFF_1_n8), .A(state1FF_state_gff_2_SFF_1_n12), 
        .ZN(state1FF_state_gff_2_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_2_SFF_1_U4 ( .B1(state1FF_state_gff_2_SFF_1_n10), .B2(state1FF_inputPar[16]), .C1(state1FF_state_gff_2_SFF_1_n11), .C2(
        state1FF_inputPar[5]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_2_SFF_1_n12) );
  INV_X1 state1FF_state_gff_2_SFF_1_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_2_SFF_1_n11) );
  INV_X1 state1FF_state_gff_2_SFF_1_U2 ( .A(state1FF_state_gff_2_SFF_1_n11), 
        .ZN(state1FF_state_gff_2_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_2_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_2_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[17]), 
        .QN(state1FF_state_gff_2_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_2_SFF_2_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_2_SFF_2_n8), .A(state1FF_state_gff_2_SFF_2_n11), 
        .ZN(state1FF_state_gff_2_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_2_SFF_2_U3 ( .B1(state1FF_state_n13), .B2(
        state1FF_inputPar[32]), .C1(state1FF_state_gff_2_SFF_2_n10), .C2(
        state1FF_inputPar[6]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_2_SFF_2_n11) );
  INV_X1 state1FF_state_gff_2_SFF_2_U2 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_2_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_2_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_2_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[33]), 
        .QN(state1FF_state_gff_2_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_2_SFF_3_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_2_SFF_3_n8), .A(state1FF_state_gff_2_SFF_3_n11), 
        .ZN(state1FF_state_gff_2_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_2_SFF_3_U3 ( .B1(state1FF_state_n13), .B2(
        state1FF_inputPar[48]), .C1(state1FF_state_gff_2_SFF_3_n10), .C2(
        state1FF_inputPar[7]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_2_SFF_3_n11) );
  INV_X1 state1FF_state_gff_2_SFF_3_U2 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_2_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_2_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_2_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[49]), 
        .QN(state1FF_state_gff_2_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_3_SFF_0_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_3_SFF_0_n8), .A(state1FF_state_gff_3_SFF_0_n12), 
        .ZN(state1FF_state_gff_3_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_3_SFF_0_U4 ( .B1(state1FF_state_gff_3_SFF_0_n10), .B2(state1FF_inputPar[1]), .C1(state1FF_state_gff_3_SFF_0_n11), .C2(
        state1FF_inputPar[8]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_3_SFF_0_n12) );
  INV_X1 state1FF_state_gff_3_SFF_0_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_3_SFF_0_n11) );
  INV_X1 state1FF_state_gff_3_SFF_0_U2 ( .A(state1FF_state_gff_3_SFF_0_n11), 
        .ZN(state1FF_state_gff_3_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_3_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_3_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[2]), 
        .QN(state1FF_state_gff_3_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_3_SFF_1_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_3_SFF_1_n8), .A(state1FF_state_gff_3_SFF_1_n12), 
        .ZN(state1FF_state_gff_3_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_3_SFF_1_U4 ( .B1(state1FF_state_gff_3_SFF_1_n10), .B2(state1FF_inputPar[17]), .C1(state1FF_state_gff_3_SFF_1_n11), .C2(
        state1FF_inputPar[9]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_3_SFF_1_n12) );
  INV_X1 state1FF_state_gff_3_SFF_1_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_3_SFF_1_n11) );
  INV_X1 state1FF_state_gff_3_SFF_1_U2 ( .A(state1FF_state_gff_3_SFF_1_n11), 
        .ZN(state1FF_state_gff_3_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_3_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_3_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[18]), 
        .QN(state1FF_state_gff_3_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_3_SFF_2_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_3_SFF_2_n8), .A(state1FF_state_gff_3_SFF_2_n12), 
        .ZN(state1FF_state_gff_3_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_3_SFF_2_U4 ( .B1(state1FF_state_gff_3_SFF_2_n10), .B2(state1FF_inputPar[33]), .C1(state1FF_state_gff_3_SFF_2_n11), .C2(
        state1FF_inputPar[10]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_3_SFF_2_n12) );
  INV_X1 state1FF_state_gff_3_SFF_2_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_3_SFF_2_n11) );
  INV_X1 state1FF_state_gff_3_SFF_2_U2 ( .A(state1FF_state_gff_3_SFF_2_n11), 
        .ZN(state1FF_state_gff_3_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_3_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_3_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[34]), 
        .QN(state1FF_state_gff_3_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_3_SFF_3_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_3_SFF_3_n8), .A(state1FF_state_gff_3_SFF_3_n12), 
        .ZN(state1FF_state_gff_3_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_3_SFF_3_U4 ( .B1(state1FF_state_gff_3_SFF_3_n10), .B2(state1FF_inputPar[49]), .C1(state1FF_state_gff_3_SFF_3_n11), .C2(
        state1FF_inputPar[11]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_3_SFF_3_n12) );
  INV_X1 state1FF_state_gff_3_SFF_3_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_3_SFF_3_n11) );
  INV_X1 state1FF_state_gff_3_SFF_3_U2 ( .A(state1FF_state_gff_3_SFF_3_n11), 
        .ZN(state1FF_state_gff_3_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_3_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_3_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[50]), 
        .QN(state1FF_state_gff_3_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_4_SFF_0_U4 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_4_SFF_0_n8), .A(state1FF_state_gff_4_SFF_0_n11), 
        .ZN(state1FF_state_gff_4_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_4_SFF_0_U3 ( .B1(state1FF_state_n13), .B2(
        state1FF_inputPar[2]), .C1(state1FF_state_gff_4_SFF_0_n10), .C2(
        state1FF_inputPar[12]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_4_SFF_0_n11) );
  INV_X1 state1FF_state_gff_4_SFF_0_U2 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_4_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_4_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_4_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[3]), 
        .QN(state1FF_state_gff_4_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_4_SFF_1_U4 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_4_SFF_1_n8), .A(state1FF_state_gff_4_SFF_1_n11), 
        .ZN(state1FF_state_gff_4_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_4_SFF_1_U3 ( .B1(state1FF_state_n13), .B2(
        state1FF_inputPar[18]), .C1(state1FF_state_gff_4_SFF_1_n10), .C2(
        state1FF_inputPar[13]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_4_SFF_1_n11) );
  INV_X1 state1FF_state_gff_4_SFF_1_U2 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_4_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_4_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_4_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[19]), 
        .QN(state1FF_state_gff_4_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_4_SFF_2_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_4_SFF_2_n7), .A(state1FF_state_gff_4_SFF_2_n11), 
        .ZN(state1FF_state_gff_4_SFF_2_n6) );
  OAI221_X1 state1FF_state_gff_4_SFF_2_U4 ( .B1(state1FF_state_gff_4_SFF_2_n9), 
        .B2(state1FF_inputPar[34]), .C1(state1FF_state_gff_4_SFF_2_n10), .C2(
        state1FF_inputPar[14]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_4_SFF_2_n11) );
  INV_X1 state1FF_state_gff_4_SFF_2_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_4_SFF_2_n10) );
  INV_X1 state1FF_state_gff_4_SFF_2_U2 ( .A(state1FF_state_gff_4_SFF_2_n10), 
        .ZN(state1FF_state_gff_4_SFF_2_n9) );
  DFF_X1 state1FF_state_gff_4_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_4_SFF_2_n6), .CK(clk), .Q(state1FF_inputPar[35]), 
        .QN(state1FF_state_gff_4_SFF_2_n7) );
  OAI21_X1 state1FF_state_gff_4_SFF_3_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_4_SFF_3_n7), .A(state1FF_state_gff_4_SFF_3_n11), 
        .ZN(state1FF_state_gff_4_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_4_SFF_3_U4 ( .B1(state1FF_state_gff_4_SFF_3_n9), 
        .B2(state1FF_inputPar[50]), .C1(state1FF_state_gff_4_SFF_3_n10), .C2(
        state1FF_inputPar[15]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_4_SFF_3_n11) );
  INV_X1 state1FF_state_gff_4_SFF_3_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_4_SFF_3_n10) );
  INV_X1 state1FF_state_gff_4_SFF_3_U2 ( .A(state1FF_state_gff_4_SFF_3_n10), 
        .ZN(state1FF_state_gff_4_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_4_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_4_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[51]), 
        .QN(state1FF_state_gff_4_SFF_3_n7) );
  OAI21_X1 state1FF_state_gff_5_SFF_0_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_5_SFF_0_n7), .A(state1FF_state_gff_5_SFF_0_n11), 
        .ZN(state1FF_state_gff_5_SFF_0_n6) );
  OAI221_X1 state1FF_state_gff_5_SFF_0_U4 ( .B1(state1FF_state_gff_5_SFF_0_n9), 
        .B2(state1FF_inputPar[3]), .C1(state1FF_state_gff_5_SFF_0_n10), .C2(
        state1FF_inputPar[16]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_5_SFF_0_n11) );
  INV_X1 state1FF_state_gff_5_SFF_0_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_5_SFF_0_n10) );
  INV_X1 state1FF_state_gff_5_SFF_0_U2 ( .A(state1FF_state_gff_5_SFF_0_n10), 
        .ZN(state1FF_state_gff_5_SFF_0_n9) );
  DFF_X1 state1FF_state_gff_5_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_5_SFF_0_n6), .CK(clk), .Q(state1FF_inputPar[4]), 
        .QN(state1FF_state_gff_5_SFF_0_n7) );
  OAI21_X1 state1FF_state_gff_5_SFF_1_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_5_SFF_1_n7), .A(state1FF_state_gff_5_SFF_1_n11), 
        .ZN(state1FF_state_gff_5_SFF_1_n6) );
  OAI221_X1 state1FF_state_gff_5_SFF_1_U4 ( .B1(state1FF_state_gff_5_SFF_1_n9), 
        .B2(state1FF_inputPar[19]), .C1(state1FF_state_gff_5_SFF_1_n10), .C2(
        state1FF_inputPar[17]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_5_SFF_1_n11) );
  INV_X1 state1FF_state_gff_5_SFF_1_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_5_SFF_1_n10) );
  INV_X1 state1FF_state_gff_5_SFF_1_U2 ( .A(state1FF_state_gff_5_SFF_1_n10), 
        .ZN(state1FF_state_gff_5_SFF_1_n9) );
  DFF_X1 state1FF_state_gff_5_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_5_SFF_1_n6), .CK(clk), .Q(state1FF_inputPar[20]), 
        .QN(state1FF_state_gff_5_SFF_1_n7) );
  OAI21_X1 state1FF_state_gff_5_SFF_2_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_5_SFF_2_n7), .A(state1FF_state_gff_5_SFF_2_n11), 
        .ZN(state1FF_state_gff_5_SFF_2_n6) );
  OAI221_X1 state1FF_state_gff_5_SFF_2_U4 ( .B1(state1FF_state_gff_5_SFF_2_n9), 
        .B2(state1FF_inputPar[35]), .C1(state1FF_state_gff_5_SFF_2_n10), .C2(
        state1FF_inputPar[18]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_5_SFF_2_n11) );
  INV_X1 state1FF_state_gff_5_SFF_2_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_5_SFF_2_n10) );
  INV_X1 state1FF_state_gff_5_SFF_2_U2 ( .A(state1FF_state_gff_5_SFF_2_n10), 
        .ZN(state1FF_state_gff_5_SFF_2_n9) );
  DFF_X1 state1FF_state_gff_5_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_5_SFF_2_n6), .CK(clk), .Q(state1FF_inputPar[36]), 
        .QN(state1FF_state_gff_5_SFF_2_n7) );
  OAI21_X1 state1FF_state_gff_5_SFF_3_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_5_SFF_3_n7), .A(state1FF_state_gff_5_SFF_3_n11), 
        .ZN(state1FF_state_gff_5_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_5_SFF_3_U4 ( .B1(state1FF_state_gff_5_SFF_3_n9), 
        .B2(state1FF_inputPar[51]), .C1(state1FF_state_gff_5_SFF_3_n10), .C2(
        state1FF_inputPar[19]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_5_SFF_3_n11) );
  INV_X1 state1FF_state_gff_5_SFF_3_U3 ( .A(state1FF_state_n13), .ZN(
        state1FF_state_gff_5_SFF_3_n10) );
  INV_X1 state1FF_state_gff_5_SFF_3_U2 ( .A(state1FF_state_gff_5_SFF_3_n10), 
        .ZN(state1FF_state_gff_5_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_5_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_5_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[52]), 
        .QN(state1FF_state_gff_5_SFF_3_n7) );
  OAI21_X1 state1FF_state_gff_6_SFF_0_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_6_SFF_0_n8), .A(state1FF_state_gff_6_SFF_0_n12), 
        .ZN(state1FF_state_gff_6_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_6_SFF_0_U4 ( .B1(state1FF_state_gff_6_SFF_0_n10), .B2(state1FF_inputPar[4]), .C1(state1FF_state_gff_6_SFF_0_n11), .C2(
        state1FF_inputPar[20]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_6_SFF_0_n12) );
  INV_X1 state1FF_state_gff_6_SFF_0_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_6_SFF_0_n11) );
  INV_X1 state1FF_state_gff_6_SFF_0_U2 ( .A(state1FF_state_gff_6_SFF_0_n11), 
        .ZN(state1FF_state_gff_6_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_6_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_6_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[5]), 
        .QN(state1FF_state_gff_6_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_6_SFF_1_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_6_SFF_1_n8), .A(state1FF_state_gff_6_SFF_1_n12), 
        .ZN(state1FF_state_gff_6_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_6_SFF_1_U4 ( .B1(state1FF_state_gff_6_SFF_1_n10), .B2(state1FF_inputPar[20]), .C1(state1FF_state_gff_6_SFF_1_n11), .C2(
        state1FF_inputPar[21]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_6_SFF_1_n12) );
  INV_X1 state1FF_state_gff_6_SFF_1_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_6_SFF_1_n11) );
  INV_X1 state1FF_state_gff_6_SFF_1_U2 ( .A(state1FF_state_gff_6_SFF_1_n11), 
        .ZN(state1FF_state_gff_6_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_6_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_6_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[21]), 
        .QN(state1FF_state_gff_6_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_6_SFF_2_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_6_SFF_2_n8), .A(state1FF_state_gff_6_SFF_2_n12), 
        .ZN(state1FF_state_gff_6_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_6_SFF_2_U4 ( .B1(state1FF_state_gff_6_SFF_2_n10), .B2(state1FF_inputPar[36]), .C1(state1FF_state_gff_6_SFF_2_n11), .C2(
        state1FF_inputPar[22]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_6_SFF_2_n12) );
  INV_X1 state1FF_state_gff_6_SFF_2_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_6_SFF_2_n11) );
  INV_X1 state1FF_state_gff_6_SFF_2_U2 ( .A(state1FF_state_gff_6_SFF_2_n11), 
        .ZN(state1FF_state_gff_6_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_6_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_6_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[37]), 
        .QN(state1FF_state_gff_6_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_6_SFF_3_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_6_SFF_3_n8), .A(state1FF_state_gff_6_SFF_3_n12), 
        .ZN(state1FF_state_gff_6_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_6_SFF_3_U4 ( .B1(state1FF_state_gff_6_SFF_3_n10), .B2(state1FF_inputPar[52]), .C1(state1FF_state_gff_6_SFF_3_n11), .C2(
        state1FF_inputPar[23]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_6_SFF_3_n12) );
  INV_X1 state1FF_state_gff_6_SFF_3_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_6_SFF_3_n11) );
  INV_X1 state1FF_state_gff_6_SFF_3_U2 ( .A(state1FF_state_gff_6_SFF_3_n11), 
        .ZN(state1FF_state_gff_6_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_6_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_6_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[53]), 
        .QN(state1FF_state_gff_6_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_7_SFF_0_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_7_SFF_0_n8), .A(state1FF_state_gff_7_SFF_0_n12), 
        .ZN(state1FF_state_gff_7_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_7_SFF_0_U4 ( .B1(state1FF_state_gff_7_SFF_0_n10), .B2(state1FF_inputPar[5]), .C1(state1FF_state_gff_7_SFF_0_n11), .C2(
        state1FF_inputPar[24]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_7_SFF_0_n12) );
  INV_X1 state1FF_state_gff_7_SFF_0_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_7_SFF_0_n11) );
  INV_X1 state1FF_state_gff_7_SFF_0_U2 ( .A(state1FF_state_gff_7_SFF_0_n11), 
        .ZN(state1FF_state_gff_7_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_7_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_7_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[6]), 
        .QN(state1FF_state_gff_7_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_7_SFF_1_U5 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_7_SFF_1_n8), .A(state1FF_state_gff_7_SFF_1_n12), 
        .ZN(state1FF_state_gff_7_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_7_SFF_1_U4 ( .B1(state1FF_state_gff_7_SFF_1_n10), .B2(state1FF_inputPar[21]), .C1(state1FF_state_gff_7_SFF_1_n11), .C2(
        state1FF_inputPar[25]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_7_SFF_1_n12) );
  INV_X1 state1FF_state_gff_7_SFF_1_U3 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_7_SFF_1_n11) );
  INV_X1 state1FF_state_gff_7_SFF_1_U2 ( .A(state1FF_state_gff_7_SFF_1_n11), 
        .ZN(state1FF_state_gff_7_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_7_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_7_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[22]), 
        .QN(state1FF_state_gff_7_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_7_SFF_2_U4 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_7_SFF_2_n8), .A(state1FF_state_gff_7_SFF_2_n11), 
        .ZN(state1FF_state_gff_7_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_7_SFF_2_U3 ( .B1(state1FF_state_n10), .B2(
        state1FF_inputPar[37]), .C1(state1FF_state_gff_7_SFF_2_n10), .C2(
        state1FF_inputPar[26]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_7_SFF_2_n11) );
  INV_X1 state1FF_state_gff_7_SFF_2_U2 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_7_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_7_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_7_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[38]), 
        .QN(state1FF_state_gff_7_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_7_SFF_3_U4 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_7_SFF_3_n8), .A(state1FF_state_gff_7_SFF_3_n11), 
        .ZN(state1FF_state_gff_7_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_7_SFF_3_U3 ( .B1(state1FF_state_n10), .B2(
        state1FF_inputPar[53]), .C1(state1FF_state_gff_7_SFF_3_n10), .C2(
        state1FF_inputPar[27]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_7_SFF_3_n11) );
  INV_X1 state1FF_state_gff_7_SFF_3_U2 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_7_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_7_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_7_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[54]), 
        .QN(state1FF_state_gff_7_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_8_SFF_0_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_8_SFF_0_n8), .A(state1FF_state_gff_8_SFF_0_n12), 
        .ZN(state1FF_state_gff_8_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_8_SFF_0_U4 ( .B1(state1FF_state_gff_8_SFF_0_n10), .B2(state1FF_inputPar[6]), .C1(state1FF_state_gff_8_SFF_0_n11), .C2(
        state1FF_inputPar[28]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_8_SFF_0_n12) );
  INV_X1 state1FF_state_gff_8_SFF_0_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_8_SFF_0_n11) );
  INV_X1 state1FF_state_gff_8_SFF_0_U2 ( .A(state1FF_state_gff_8_SFF_0_n11), 
        .ZN(state1FF_state_gff_8_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_8_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_8_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[7]), 
        .QN(state1FF_state_gff_8_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_8_SFF_1_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_8_SFF_1_n8), .A(state1FF_state_gff_8_SFF_1_n12), 
        .ZN(state1FF_state_gff_8_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_8_SFF_1_U4 ( .B1(state1FF_state_gff_8_SFF_1_n10), .B2(state1FF_inputPar[22]), .C1(state1FF_state_gff_8_SFF_1_n11), .C2(
        state1FF_inputPar[29]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_8_SFF_1_n12) );
  INV_X1 state1FF_state_gff_8_SFF_1_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_8_SFF_1_n11) );
  INV_X1 state1FF_state_gff_8_SFF_1_U2 ( .A(state1FF_state_gff_8_SFF_1_n11), 
        .ZN(state1FF_state_gff_8_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_8_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_8_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[23]), 
        .QN(state1FF_state_gff_8_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_8_SFF_2_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_8_SFF_2_n7), .A(state1FF_state_gff_8_SFF_2_n11), 
        .ZN(state1FF_state_gff_8_SFF_2_n6) );
  OAI221_X1 state1FF_state_gff_8_SFF_2_U4 ( .B1(state1FF_state_gff_8_SFF_2_n9), 
        .B2(state1FF_inputPar[38]), .C1(state1FF_state_gff_8_SFF_2_n10), .C2(
        state1FF_inputPar[30]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_8_SFF_2_n11) );
  INV_X1 state1FF_state_gff_8_SFF_2_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_8_SFF_2_n10) );
  INV_X1 state1FF_state_gff_8_SFF_2_U2 ( .A(state1FF_state_gff_8_SFF_2_n10), 
        .ZN(state1FF_state_gff_8_SFF_2_n9) );
  DFF_X1 state1FF_state_gff_8_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_8_SFF_2_n6), .CK(clk), .Q(state1FF_inputPar[39]), 
        .QN(state1FF_state_gff_8_SFF_2_n7) );
  OAI21_X1 state1FF_state_gff_8_SFF_3_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_8_SFF_3_n7), .A(state1FF_state_gff_8_SFF_3_n11), 
        .ZN(state1FF_state_gff_8_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_8_SFF_3_U4 ( .B1(state1FF_state_gff_8_SFF_3_n9), 
        .B2(state1FF_inputPar[54]), .C1(state1FF_state_gff_8_SFF_3_n10), .C2(
        state1FF_inputPar[31]), .A(state1FF_state_n6), .ZN(
        state1FF_state_gff_8_SFF_3_n11) );
  INV_X1 state1FF_state_gff_8_SFF_3_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_8_SFF_3_n10) );
  INV_X1 state1FF_state_gff_8_SFF_3_U2 ( .A(state1FF_state_gff_8_SFF_3_n10), 
        .ZN(state1FF_state_gff_8_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_8_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_8_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[55]), 
        .QN(state1FF_state_gff_8_SFF_3_n7) );
  OAI21_X1 state1FF_state_gff_9_SFF_0_U5 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_9_SFF_0_n7), .A(state1FF_state_gff_9_SFF_0_n11), 
        .ZN(state1FF_state_gff_9_SFF_0_n6) );
  OAI221_X1 state1FF_state_gff_9_SFF_0_U4 ( .B1(state1FF_state_gff_9_SFF_0_n9), 
        .B2(state1FF_inputPar[7]), .C1(state1FF_state_gff_9_SFF_0_n10), .C2(
        state1FF_inputPar[32]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_9_SFF_0_n11) );
  INV_X1 state1FF_state_gff_9_SFF_0_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_9_SFF_0_n10) );
  INV_X1 state1FF_state_gff_9_SFF_0_U2 ( .A(state1FF_state_gff_9_SFF_0_n10), 
        .ZN(state1FF_state_gff_9_SFF_0_n9) );
  DFF_X1 state1FF_state_gff_9_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_9_SFF_0_n6), .CK(clk), .Q(state1FF_inputPar[8]), 
        .QN(state1FF_state_gff_9_SFF_0_n7) );
  OAI21_X1 state1FF_state_gff_9_SFF_1_U5 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_9_SFF_1_n7), .A(state1FF_state_gff_9_SFF_1_n11), 
        .ZN(state1FF_state_gff_9_SFF_1_n6) );
  OAI221_X1 state1FF_state_gff_9_SFF_1_U4 ( .B1(state1FF_state_gff_9_SFF_1_n9), 
        .B2(state1FF_inputPar[23]), .C1(state1FF_state_gff_9_SFF_1_n10), .C2(
        state1FF_inputPar[33]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_9_SFF_1_n11) );
  INV_X1 state1FF_state_gff_9_SFF_1_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_9_SFF_1_n10) );
  INV_X1 state1FF_state_gff_9_SFF_1_U2 ( .A(state1FF_state_gff_9_SFF_1_n10), 
        .ZN(state1FF_state_gff_9_SFF_1_n9) );
  DFF_X1 state1FF_state_gff_9_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_9_SFF_1_n6), .CK(clk), .Q(state1FF_inputPar[24]), 
        .QN(state1FF_state_gff_9_SFF_1_n7) );
  OAI21_X1 state1FF_state_gff_9_SFF_2_U5 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_9_SFF_2_n7), .A(state1FF_state_gff_9_SFF_2_n11), 
        .ZN(state1FF_state_gff_9_SFF_2_n6) );
  OAI221_X1 state1FF_state_gff_9_SFF_2_U4 ( .B1(state1FF_state_gff_9_SFF_2_n9), 
        .B2(state1FF_inputPar[39]), .C1(state1FF_state_gff_9_SFF_2_n10), .C2(
        state1FF_inputPar[34]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_9_SFF_2_n11) );
  INV_X1 state1FF_state_gff_9_SFF_2_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_9_SFF_2_n10) );
  INV_X1 state1FF_state_gff_9_SFF_2_U2 ( .A(state1FF_state_gff_9_SFF_2_n10), 
        .ZN(state1FF_state_gff_9_SFF_2_n9) );
  DFF_X1 state1FF_state_gff_9_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_9_SFF_2_n6), .CK(clk), .Q(state1FF_inputPar[40]), 
        .QN(state1FF_state_gff_9_SFF_2_n7) );
  OAI21_X1 state1FF_state_gff_9_SFF_3_U5 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_9_SFF_3_n7), .A(state1FF_state_gff_9_SFF_3_n11), 
        .ZN(state1FF_state_gff_9_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_9_SFF_3_U4 ( .B1(state1FF_state_gff_9_SFF_3_n9), 
        .B2(state1FF_inputPar[55]), .C1(state1FF_state_gff_9_SFF_3_n10), .C2(
        state1FF_inputPar[35]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_9_SFF_3_n11) );
  INV_X1 state1FF_state_gff_9_SFF_3_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_9_SFF_3_n10) );
  INV_X1 state1FF_state_gff_9_SFF_3_U2 ( .A(state1FF_state_gff_9_SFF_3_n10), 
        .ZN(state1FF_state_gff_9_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_9_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_9_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[56]), 
        .QN(state1FF_state_gff_9_SFF_3_n7) );
  OAI21_X1 state1FF_state_gff_10_SFF_0_U4 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_10_SFF_0_n8), .A(state1FF_state_gff_10_SFF_0_n11), 
        .ZN(state1FF_state_gff_10_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_10_SFF_0_U3 ( .B1(state1FF_state_n10), .B2(
        state1FF_inputPar[8]), .C1(state1FF_state_gff_10_SFF_0_n10), .C2(
        state1FF_inputPar[36]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_10_SFF_0_n11) );
  INV_X1 state1FF_state_gff_10_SFF_0_U2 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_10_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_10_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_10_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[9]), 
        .QN(state1FF_state_gff_10_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_10_SFF_1_U4 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_10_SFF_1_n8), .A(state1FF_state_gff_10_SFF_1_n11), 
        .ZN(state1FF_state_gff_10_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_10_SFF_1_U3 ( .B1(state1FF_state_n10), .B2(
        state1FF_inputPar[24]), .C1(state1FF_state_gff_10_SFF_1_n10), .C2(
        state1FF_inputPar[37]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_10_SFF_1_n11) );
  INV_X1 state1FF_state_gff_10_SFF_1_U2 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_10_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_10_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_10_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[25]), 
        .QN(state1FF_state_gff_10_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_10_SFF_2_U4 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_10_SFF_2_n8), .A(state1FF_state_gff_10_SFF_2_n11), 
        .ZN(state1FF_state_gff_10_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_10_SFF_2_U3 ( .B1(state1FF_state_n10), .B2(
        state1FF_inputPar[40]), .C1(state1FF_state_gff_10_SFF_2_n10), .C2(
        state1FF_inputPar[38]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_10_SFF_2_n11) );
  INV_X1 state1FF_state_gff_10_SFF_2_U2 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_10_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_10_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_10_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[41]), 
        .QN(state1FF_state_gff_10_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_10_SFF_3_U4 ( .B1(state1FF_state_n7), .B2(
        state1FF_state_gff_10_SFF_3_n8), .A(state1FF_state_gff_10_SFF_3_n11), 
        .ZN(state1FF_state_gff_10_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_10_SFF_3_U3 ( .B1(state1FF_state_n10), .B2(
        state1FF_inputPar[56]), .C1(state1FF_state_gff_10_SFF_3_n10), .C2(
        state1FF_inputPar[39]), .A(state1FF_state_n7), .ZN(
        state1FF_state_gff_10_SFF_3_n11) );
  INV_X1 state1FF_state_gff_10_SFF_3_U2 ( .A(state1FF_state_n10), .ZN(
        state1FF_state_gff_10_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_10_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_10_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[57]), 
        .QN(state1FF_state_gff_10_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_11_SFF_0_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_11_SFF_0_n8), .A(state1FF_state_gff_11_SFF_0_n12), 
        .ZN(state1FF_state_gff_11_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_11_SFF_0_U4 ( .B1(
        state1FF_state_gff_11_SFF_0_n10), .B2(state1FF_inputPar[9]), .C1(
        state1FF_state_gff_11_SFF_0_n11), .C2(state1FF_inputPar[40]), .A(
        state1FF_state_n8), .ZN(state1FF_state_gff_11_SFF_0_n12) );
  INV_X1 state1FF_state_gff_11_SFF_0_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_11_SFF_0_n11) );
  INV_X1 state1FF_state_gff_11_SFF_0_U2 ( .A(state1FF_state_gff_11_SFF_0_n11), 
        .ZN(state1FF_state_gff_11_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_11_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_11_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[10]), 
        .QN(state1FF_state_gff_11_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_11_SFF_1_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_11_SFF_1_n8), .A(state1FF_state_gff_11_SFF_1_n12), 
        .ZN(state1FF_state_gff_11_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_11_SFF_1_U4 ( .B1(
        state1FF_state_gff_11_SFF_1_n10), .B2(state1FF_inputPar[25]), .C1(
        state1FF_state_gff_11_SFF_1_n11), .C2(state1FF_inputPar[41]), .A(
        state1FF_state_n8), .ZN(state1FF_state_gff_11_SFF_1_n12) );
  INV_X1 state1FF_state_gff_11_SFF_1_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_11_SFF_1_n11) );
  INV_X1 state1FF_state_gff_11_SFF_1_U2 ( .A(state1FF_state_gff_11_SFF_1_n11), 
        .ZN(state1FF_state_gff_11_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_11_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_11_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[26]), 
        .QN(state1FF_state_gff_11_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_11_SFF_2_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_11_SFF_2_n8), .A(state1FF_state_gff_11_SFF_2_n12), 
        .ZN(state1FF_state_gff_11_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_11_SFF_2_U4 ( .B1(
        state1FF_state_gff_11_SFF_2_n10), .B2(state1FF_inputPar[41]), .C1(
        state1FF_state_gff_11_SFF_2_n11), .C2(state1FF_inputPar[42]), .A(
        state1FF_state_n8), .ZN(state1FF_state_gff_11_SFF_2_n12) );
  INV_X1 state1FF_state_gff_11_SFF_2_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_11_SFF_2_n11) );
  INV_X1 state1FF_state_gff_11_SFF_2_U2 ( .A(state1FF_state_gff_11_SFF_2_n11), 
        .ZN(state1FF_state_gff_11_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_11_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_11_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[42]), 
        .QN(state1FF_state_gff_11_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_11_SFF_3_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_11_SFF_3_n8), .A(state1FF_state_gff_11_SFF_3_n12), 
        .ZN(state1FF_state_gff_11_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_11_SFF_3_U4 ( .B1(
        state1FF_state_gff_11_SFF_3_n10), .B2(state1FF_inputPar[57]), .C1(
        state1FF_state_gff_11_SFF_3_n11), .C2(state1FF_inputPar[43]), .A(
        state1FF_state_n8), .ZN(state1FF_state_gff_11_SFF_3_n12) );
  INV_X1 state1FF_state_gff_11_SFF_3_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_11_SFF_3_n11) );
  INV_X1 state1FF_state_gff_11_SFF_3_U2 ( .A(state1FF_state_gff_11_SFF_3_n11), 
        .ZN(state1FF_state_gff_11_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_11_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_11_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[58]), 
        .QN(state1FF_state_gff_11_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_12_SFF_0_U4 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_12_SFF_0_n8), .A(state1FF_state_gff_12_SFF_0_n11), 
        .ZN(state1FF_state_gff_12_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_12_SFF_0_U3 ( .B1(state1FF_state_n11), .B2(
        state1FF_inputPar[10]), .C1(state1FF_state_gff_12_SFF_0_n10), .C2(
        state1FF_inputPar[44]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_12_SFF_0_n11) );
  INV_X1 state1FF_state_gff_12_SFF_0_U2 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_12_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_12_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_12_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[11]), 
        .QN(state1FF_state_gff_12_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_12_SFF_1_U4 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_12_SFF_1_n8), .A(state1FF_state_gff_12_SFF_1_n11), 
        .ZN(state1FF_state_gff_12_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_12_SFF_1_U3 ( .B1(state1FF_state_n11), .B2(
        state1FF_inputPar[26]), .C1(state1FF_state_gff_12_SFF_1_n10), .C2(
        state1FF_inputPar[45]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_12_SFF_1_n11) );
  INV_X1 state1FF_state_gff_12_SFF_1_U2 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_12_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_12_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_12_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[27]), 
        .QN(state1FF_state_gff_12_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_12_SFF_2_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_12_SFF_2_n7), .A(state1FF_state_gff_12_SFF_2_n11), 
        .ZN(state1FF_state_gff_12_SFF_2_n6) );
  OAI221_X1 state1FF_state_gff_12_SFF_2_U4 ( .B1(
        state1FF_state_gff_12_SFF_2_n9), .B2(state1FF_inputPar[42]), .C1(
        state1FF_state_gff_12_SFF_2_n10), .C2(state1FF_inputPar[46]), .A(
        state1FF_state_n8), .ZN(state1FF_state_gff_12_SFF_2_n11) );
  INV_X1 state1FF_state_gff_12_SFF_2_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_12_SFF_2_n10) );
  INV_X1 state1FF_state_gff_12_SFF_2_U2 ( .A(state1FF_state_gff_12_SFF_2_n10), 
        .ZN(state1FF_state_gff_12_SFF_2_n9) );
  DFF_X1 state1FF_state_gff_12_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_12_SFF_2_n6), .CK(clk), .Q(state1FF_inputPar[43]), 
        .QN(state1FF_state_gff_12_SFF_2_n7) );
  OAI21_X1 state1FF_state_gff_12_SFF_3_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_12_SFF_3_n7), .A(state1FF_state_gff_12_SFF_3_n11), 
        .ZN(state1FF_state_gff_12_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_12_SFF_3_U4 ( .B1(
        state1FF_state_gff_12_SFF_3_n9), .B2(state1FF_inputPar[58]), .C1(
        state1FF_state_gff_12_SFF_3_n10), .C2(state1FF_inputPar[47]), .A(
        state1FF_state_n8), .ZN(state1FF_state_gff_12_SFF_3_n11) );
  INV_X1 state1FF_state_gff_12_SFF_3_U3 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_12_SFF_3_n10) );
  INV_X1 state1FF_state_gff_12_SFF_3_U2 ( .A(state1FF_state_gff_12_SFF_3_n10), 
        .ZN(state1FF_state_gff_12_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_12_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_12_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[59]), 
        .QN(state1FF_state_gff_12_SFF_3_n7) );
  OAI21_X1 state1FF_state_gff_13_SFF_0_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_13_SFF_0_n7), .A(state1FF_state_gff_13_SFF_0_n11), 
        .ZN(state1FF_state_gff_13_SFF_0_n6) );
  OAI221_X1 state1FF_state_gff_13_SFF_0_U4 ( .B1(
        state1FF_state_gff_13_SFF_0_n9), .B2(state1FF_inputPar[11]), .C1(
        state1FF_state_gff_13_SFF_0_n10), .C2(state1FF_inputPar[48]), .A(
        state1FF_state_n6), .ZN(state1FF_state_gff_13_SFF_0_n11) );
  INV_X1 state1FF_state_gff_13_SFF_0_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_13_SFF_0_n10) );
  INV_X1 state1FF_state_gff_13_SFF_0_U2 ( .A(state1FF_state_gff_13_SFF_0_n10), 
        .ZN(state1FF_state_gff_13_SFF_0_n9) );
  DFF_X1 state1FF_state_gff_13_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_13_SFF_0_n6), .CK(clk), .Q(state1FF_inputPar[12]), 
        .QN(state1FF_state_gff_13_SFF_0_n7) );
  OAI21_X1 state1FF_state_gff_13_SFF_1_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_13_SFF_1_n7), .A(state1FF_state_gff_13_SFF_1_n11), 
        .ZN(state1FF_state_gff_13_SFF_1_n6) );
  OAI221_X1 state1FF_state_gff_13_SFF_1_U4 ( .B1(
        state1FF_state_gff_13_SFF_1_n9), .B2(state1FF_inputPar[27]), .C1(
        state1FF_state_gff_13_SFF_1_n10), .C2(state1FF_inputPar[49]), .A(
        state1FF_state_n6), .ZN(state1FF_state_gff_13_SFF_1_n11) );
  INV_X1 state1FF_state_gff_13_SFF_1_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_13_SFF_1_n10) );
  INV_X1 state1FF_state_gff_13_SFF_1_U2 ( .A(state1FF_state_gff_13_SFF_1_n10), 
        .ZN(state1FF_state_gff_13_SFF_1_n9) );
  DFF_X1 state1FF_state_gff_13_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_13_SFF_1_n6), .CK(clk), .Q(state1FF_inputPar[28]), 
        .QN(state1FF_state_gff_13_SFF_1_n7) );
  OAI21_X1 state1FF_state_gff_13_SFF_2_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_13_SFF_2_n7), .A(state1FF_state_gff_13_SFF_2_n11), 
        .ZN(state1FF_state_gff_13_SFF_2_n6) );
  OAI221_X1 state1FF_state_gff_13_SFF_2_U4 ( .B1(
        state1FF_state_gff_13_SFF_2_n9), .B2(state1FF_inputPar[43]), .C1(
        state1FF_state_gff_13_SFF_2_n10), .C2(state1FF_inputPar[50]), .A(
        state1FF_state_n6), .ZN(state1FF_state_gff_13_SFF_2_n11) );
  INV_X1 state1FF_state_gff_13_SFF_2_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_13_SFF_2_n10) );
  INV_X1 state1FF_state_gff_13_SFF_2_U2 ( .A(state1FF_state_gff_13_SFF_2_n10), 
        .ZN(state1FF_state_gff_13_SFF_2_n9) );
  DFF_X1 state1FF_state_gff_13_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_13_SFF_2_n6), .CK(clk), .Q(state1FF_inputPar[44]), 
        .QN(state1FF_state_gff_13_SFF_2_n7) );
  OAI21_X1 state1FF_state_gff_13_SFF_3_U5 ( .B1(state1FF_state_n6), .B2(
        state1FF_state_gff_13_SFF_3_n7), .A(state1FF_state_gff_13_SFF_3_n11), 
        .ZN(state1FF_state_gff_13_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_13_SFF_3_U4 ( .B1(
        state1FF_state_gff_13_SFF_3_n9), .B2(state1FF_inputPar[59]), .C1(
        state1FF_state_gff_13_SFF_3_n10), .C2(state1FF_inputPar[51]), .A(
        state1FF_state_n6), .ZN(state1FF_state_gff_13_SFF_3_n11) );
  INV_X1 state1FF_state_gff_13_SFF_3_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_13_SFF_3_n10) );
  INV_X1 state1FF_state_gff_13_SFF_3_U2 ( .A(state1FF_state_gff_13_SFF_3_n10), 
        .ZN(state1FF_state_gff_13_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_13_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_13_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[60]), 
        .QN(state1FF_state_gff_13_SFF_3_n7) );
  OAI21_X1 state1FF_state_gff_14_SFF_0_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_14_SFF_0_n8), .A(state1FF_state_gff_14_SFF_0_n11), 
        .ZN(state1FF_state_gff_14_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_14_SFF_0_U3 ( .B1(state1FF_state_n11), .B2(
        state1FF_inputPar[12]), .C1(state1FF_state_gff_14_SFF_0_n10), .C2(
        state1FF_inputPar[52]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_14_SFF_0_n11) );
  INV_X1 state1FF_state_gff_14_SFF_0_U2 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_14_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_14_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_14_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[13]), 
        .QN(state1FF_state_gff_14_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_14_SFF_1_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_14_SFF_1_n8), .A(state1FF_state_gff_14_SFF_1_n11), 
        .ZN(state1FF_state_gff_14_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_14_SFF_1_U3 ( .B1(state1FF_state_n11), .B2(
        state1FF_inputPar[28]), .C1(state1FF_state_gff_14_SFF_1_n10), .C2(
        state1FF_inputPar[53]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_14_SFF_1_n11) );
  INV_X1 state1FF_state_gff_14_SFF_1_U2 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_14_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_14_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_14_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[29]), 
        .QN(state1FF_state_gff_14_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_14_SFF_2_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_14_SFF_2_n8), .A(state1FF_state_gff_14_SFF_2_n11), 
        .ZN(state1FF_state_gff_14_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_14_SFF_2_U3 ( .B1(state1FF_state_n11), .B2(
        state1FF_inputPar[44]), .C1(state1FF_state_gff_14_SFF_2_n10), .C2(
        state1FF_inputPar[54]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_14_SFF_2_n11) );
  INV_X1 state1FF_state_gff_14_SFF_2_U2 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_14_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_14_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_14_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[45]), 
        .QN(state1FF_state_gff_14_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_14_SFF_3_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_14_SFF_3_n8), .A(state1FF_state_gff_14_SFF_3_n11), 
        .ZN(state1FF_state_gff_14_SFF_3_n7) );
  OAI221_X1 state1FF_state_gff_14_SFF_3_U3 ( .B1(state1FF_state_n11), .B2(
        state1FF_inputPar[60]), .C1(state1FF_state_gff_14_SFF_3_n10), .C2(
        state1FF_inputPar[55]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_14_SFF_3_n11) );
  INV_X1 state1FF_state_gff_14_SFF_3_U2 ( .A(state1FF_state_n11), .ZN(
        state1FF_state_gff_14_SFF_3_n10) );
  DFF_X1 state1FF_state_gff_14_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_14_SFF_3_n7), .CK(clk), .Q(state1FF_inputPar[61]), 
        .QN(state1FF_state_gff_14_SFF_3_n8) );
  OAI21_X1 state1FF_state_gff_15_SFF_0_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_15_SFF_0_n8), .A(state1FF_state_gff_15_SFF_0_n11), 
        .ZN(state1FF_state_gff_15_SFF_0_n7) );
  OAI221_X1 state1FF_state_gff_15_SFF_0_U3 ( .B1(state1FF_state_n12), .B2(
        state1FF_inputPar[13]), .C1(state1FF_state_gff_15_SFF_0_n10), .C2(
        state1FF_inputPar[56]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_15_SFF_0_n11) );
  INV_X1 state1FF_state_gff_15_SFF_0_U2 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_15_SFF_0_n10) );
  DFF_X1 state1FF_state_gff_15_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_15_SFF_0_n7), .CK(clk), .Q(state1FF_inputPar[14]), 
        .QN(state1FF_state_gff_15_SFF_0_n8) );
  OAI21_X1 state1FF_state_gff_15_SFF_1_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_15_SFF_1_n8), .A(state1FF_state_gff_15_SFF_1_n11), 
        .ZN(state1FF_state_gff_15_SFF_1_n7) );
  OAI221_X1 state1FF_state_gff_15_SFF_1_U3 ( .B1(state1FF_state_n12), .B2(
        state1FF_inputPar[29]), .C1(state1FF_state_gff_15_SFF_1_n10), .C2(
        state1FF_inputPar[57]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_15_SFF_1_n11) );
  INV_X1 state1FF_state_gff_15_SFF_1_U2 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_15_SFF_1_n10) );
  DFF_X1 state1FF_state_gff_15_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_15_SFF_1_n7), .CK(clk), .Q(state1FF_inputPar[30]), 
        .QN(state1FF_state_gff_15_SFF_1_n8) );
  OAI21_X1 state1FF_state_gff_15_SFF_2_U4 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_15_SFF_2_n8), .A(state1FF_state_gff_15_SFF_2_n11), 
        .ZN(state1FF_state_gff_15_SFF_2_n7) );
  OAI221_X1 state1FF_state_gff_15_SFF_2_U3 ( .B1(state1FF_state_n12), .B2(
        state1FF_inputPar[45]), .C1(state1FF_state_gff_15_SFF_2_n10), .C2(
        state1FF_inputPar[58]), .A(state1FF_state_n9), .ZN(
        state1FF_state_gff_15_SFF_2_n11) );
  INV_X1 state1FF_state_gff_15_SFF_2_U2 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_15_SFF_2_n10) );
  DFF_X1 state1FF_state_gff_15_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_15_SFF_2_n7), .CK(clk), .Q(state1FF_inputPar[46]), 
        .QN(state1FF_state_gff_15_SFF_2_n8) );
  OAI21_X1 state1FF_state_gff_15_SFF_3_U5 ( .B1(state1FF_state_n9), .B2(
        state1FF_state_gff_15_SFF_3_n7), .A(state1FF_state_gff_15_SFF_3_n11), 
        .ZN(state1FF_state_gff_15_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_15_SFF_3_U4 ( .B1(
        state1FF_state_gff_15_SFF_3_n9), .B2(state1FF_inputPar[61]), .C1(
        state1FF_state_gff_15_SFF_3_n10), .C2(state1FF_inputPar[59]), .A(
        state1FF_state_n9), .ZN(state1FF_state_gff_15_SFF_3_n11) );
  INV_X1 state1FF_state_gff_15_SFF_3_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_15_SFF_3_n10) );
  INV_X1 state1FF_state_gff_15_SFF_3_U2 ( .A(state1FF_state_gff_15_SFF_3_n10), 
        .ZN(state1FF_state_gff_15_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_15_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_15_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[62]), 
        .QN(state1FF_state_gff_15_SFF_3_n7) );
  OAI21_X1 state1FF_state_gff_16_SFF_0_U5 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_16_SFF_0_n7), .A(state1FF_state_gff_16_SFF_0_n11), 
        .ZN(state1FF_state_gff_16_SFF_0_n6) );
  OAI221_X1 state1FF_state_gff_16_SFF_0_U4 ( .B1(
        state1FF_state_gff_16_SFF_0_n9), .B2(state1FF_inputPar[14]), .C1(
        state1FF_state_gff_16_SFF_0_n10), .C2(state1FF_inputPar[60]), .A(
        state1FF_state_n8), .ZN(state1FF_state_gff_16_SFF_0_n11) );
  INV_X1 state1FF_state_gff_16_SFF_0_U3 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_16_SFF_0_n10) );
  INV_X1 state1FF_state_gff_16_SFF_0_U2 ( .A(state1FF_state_gff_16_SFF_0_n10), 
        .ZN(state1FF_state_gff_16_SFF_0_n9) );
  DFF_X1 state1FF_state_gff_16_SFF_0_Cell_reg ( .D(
        state1FF_state_gff_16_SFF_0_n6), .CK(clk), .Q(state1FF_inputPar[15]), 
        .QN(state1FF_state_gff_16_SFF_0_n7) );
  OAI21_X1 state1FF_state_gff_16_SFF_1_U4 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_16_SFF_1_n7), .A(state1FF_state_gff_16_SFF_1_n10), 
        .ZN(state1FF_state_gff_16_SFF_1_n6) );
  OAI221_X1 state1FF_state_gff_16_SFF_1_U3 ( .B1(state1FF_state_n12), .B2(
        state1FF_inputPar[30]), .C1(state1FF_state_gff_16_SFF_1_n9), .C2(
        state1FF_inputPar[61]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_16_SFF_1_n10) );
  INV_X1 state1FF_state_gff_16_SFF_1_U2 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_16_SFF_1_n9) );
  DFF_X1 state1FF_state_gff_16_SFF_1_Cell_reg ( .D(
        state1FF_state_gff_16_SFF_1_n6), .CK(clk), .Q(state1FF_inputPar[31]), 
        .QN(state1FF_state_gff_16_SFF_1_n7) );
  OAI21_X1 state1FF_state_gff_16_SFF_2_U4 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_16_SFF_2_n7), .A(state1FF_state_gff_16_SFF_2_n10), 
        .ZN(state1FF_state_gff_16_SFF_2_n6) );
  OAI221_X1 state1FF_state_gff_16_SFF_2_U3 ( .B1(state1FF_state_n12), .B2(
        state1FF_inputPar[46]), .C1(state1FF_state_gff_16_SFF_2_n9), .C2(
        state1FF_inputPar[62]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_16_SFF_2_n10) );
  INV_X1 state1FF_state_gff_16_SFF_2_U2 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_16_SFF_2_n9) );
  DFF_X1 state1FF_state_gff_16_SFF_2_Cell_reg ( .D(
        state1FF_state_gff_16_SFF_2_n6), .CK(clk), .Q(state1FF_inputPar[47]), 
        .QN(state1FF_state_gff_16_SFF_2_n7) );
  OAI21_X1 state1FF_state_gff_16_SFF_3_U4 ( .B1(state1FF_state_n8), .B2(
        state1FF_state_gff_16_SFF_3_n7), .A(state1FF_state_gff_16_SFF_3_n10), 
        .ZN(state1FF_state_gff_16_SFF_3_n6) );
  OAI221_X1 state1FF_state_gff_16_SFF_3_U3 ( .B1(state1FF_state_n12), .B2(
        state1FF_inputPar[62]), .C1(state1FF_state_gff_16_SFF_3_n9), .C2(
        state1FF_inputPar[63]), .A(state1FF_state_n8), .ZN(
        state1FF_state_gff_16_SFF_3_n10) );
  INV_X1 state1FF_state_gff_16_SFF_3_U2 ( .A(state1FF_state_n12), .ZN(
        state1FF_state_gff_16_SFF_3_n9) );
  DFF_X1 state1FF_state_gff_16_SFF_3_Cell_reg ( .D(
        state1FF_state_gff_16_SFF_3_n6), .CK(clk), .Q(state1FF_inputPar[63]), 
        .QN(state1FF_state_gff_16_SFF_3_n7) );
  MUX2_X1 state2FF_U5 ( .A(sboxOut2[2]), .B(dataIn2[2]), .S(n4), .Z(
        state2FF_n1) );
  MUX2_X1 state2FF_U4 ( .A(sboxOut2[1]), .B(dataIn2[1]), .S(n4), .Z(
        state2FF_n2) );
  MUX2_X1 state2FF_U3 ( .A(sboxOut2[0]), .B(dataIn2[0]), .S(n4), .Z(
        state2FF_n3) );
  MUX2_X1 state2FF_U2 ( .A(sboxOut2[3]), .B(dataIn2[3]), .S(n4), .Z(
        state2FF_n4) );
  BUF_X1 state2FF_state_U8 ( .A(selP), .Z(state2FF_state_n12) );
  BUF_X1 state2FF_state_U7 ( .A(selP), .Z(state2FF_state_n10) );
  BUF_X1 state2FF_state_U6 ( .A(selP), .Z(state2FF_state_n13) );
  BUF_X1 state2FF_state_U5 ( .A(selP), .Z(state2FF_state_n11) );
  BUF_X2 state2FF_state_U4 ( .A(enData), .Z(state2FF_state_n9) );
  BUF_X2 state2FF_state_U3 ( .A(enData), .Z(state2FF_state_n6) );
  BUF_X2 state2FF_state_U2 ( .A(enData), .Z(state2FF_state_n7) );
  BUF_X2 state2FF_state_U1 ( .A(enData), .Z(state2FF_state_n8) );
  OAI21_X1 state2FF_state_gff_1_SFF_0_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_1_SFF_0_n8), .A(state2FF_state_gff_1_SFF_0_n12), 
        .ZN(state2FF_state_gff_1_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_1_SFF_0_U4 ( .B1(state2FF_state_gff_1_SFF_0_n10), .B2(state2FF_n3), .C1(state2FF_state_gff_1_SFF_0_n11), .C2(
        state2FF_inputPar[0]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_1_SFF_0_n12) );
  INV_X1 state2FF_state_gff_1_SFF_0_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_1_SFF_0_n11) );
  INV_X1 state2FF_state_gff_1_SFF_0_U2 ( .A(state2FF_state_gff_1_SFF_0_n11), 
        .ZN(state2FF_state_gff_1_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_1_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_1_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[0]), 
        .QN(state2FF_state_gff_1_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_1_SFF_1_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_1_SFF_1_n8), .A(state2FF_state_gff_1_SFF_1_n12), 
        .ZN(state2FF_state_gff_1_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_1_SFF_1_U4 ( .B1(state2FF_state_gff_1_SFF_1_n10), .B2(state2FF_n2), .C1(state2FF_state_gff_1_SFF_1_n11), .C2(
        state2FF_inputPar[1]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_1_SFF_1_n12) );
  INV_X1 state2FF_state_gff_1_SFF_1_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_1_SFF_1_n11) );
  INV_X1 state2FF_state_gff_1_SFF_1_U2 ( .A(state2FF_state_gff_1_SFF_1_n11), 
        .ZN(state2FF_state_gff_1_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_1_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_1_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[16]), 
        .QN(state2FF_state_gff_1_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_1_SFF_2_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_1_SFF_2_n8), .A(state2FF_state_gff_1_SFF_2_n12), 
        .ZN(state2FF_state_gff_1_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_1_SFF_2_U4 ( .B1(state2FF_state_gff_1_SFF_2_n10), .B2(state2FF_n1), .C1(state2FF_state_gff_1_SFF_2_n11), .C2(
        state2FF_inputPar[2]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_1_SFF_2_n12) );
  INV_X1 state2FF_state_gff_1_SFF_2_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_1_SFF_2_n11) );
  INV_X1 state2FF_state_gff_1_SFF_2_U2 ( .A(state2FF_state_gff_1_SFF_2_n11), 
        .ZN(state2FF_state_gff_1_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_1_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_1_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[32]), 
        .QN(state2FF_state_gff_1_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_1_SFF_3_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_1_SFF_3_n8), .A(state2FF_state_gff_1_SFF_3_n12), 
        .ZN(state2FF_state_gff_1_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_1_SFF_3_U4 ( .B1(state2FF_state_gff_1_SFF_3_n10), .B2(state2FF_n4), .C1(state2FF_state_gff_1_SFF_3_n11), .C2(
        state2FF_inputPar[3]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_1_SFF_3_n12) );
  INV_X1 state2FF_state_gff_1_SFF_3_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_1_SFF_3_n11) );
  INV_X1 state2FF_state_gff_1_SFF_3_U2 ( .A(state2FF_state_gff_1_SFF_3_n11), 
        .ZN(state2FF_state_gff_1_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_1_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_1_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[48]), 
        .QN(state2FF_state_gff_1_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_2_SFF_0_U5 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_2_SFF_0_n8), .A(state2FF_state_gff_2_SFF_0_n12), 
        .ZN(state2FF_state_gff_2_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_2_SFF_0_U4 ( .B1(state2FF_state_gff_2_SFF_0_n10), .B2(state2FF_inputPar[0]), .C1(state2FF_state_gff_2_SFF_0_n11), .C2(
        state2FF_inputPar[4]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_2_SFF_0_n12) );
  INV_X1 state2FF_state_gff_2_SFF_0_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_2_SFF_0_n11) );
  INV_X1 state2FF_state_gff_2_SFF_0_U2 ( .A(state2FF_state_gff_2_SFF_0_n11), 
        .ZN(state2FF_state_gff_2_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_2_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_2_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[1]), 
        .QN(state2FF_state_gff_2_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_2_SFF_1_U5 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_2_SFF_1_n8), .A(state2FF_state_gff_2_SFF_1_n12), 
        .ZN(state2FF_state_gff_2_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_2_SFF_1_U4 ( .B1(state2FF_state_gff_2_SFF_1_n10), .B2(state2FF_inputPar[16]), .C1(state2FF_state_gff_2_SFF_1_n11), .C2(
        state2FF_inputPar[5]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_2_SFF_1_n12) );
  INV_X1 state2FF_state_gff_2_SFF_1_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_2_SFF_1_n11) );
  INV_X1 state2FF_state_gff_2_SFF_1_U2 ( .A(state2FF_state_gff_2_SFF_1_n11), 
        .ZN(state2FF_state_gff_2_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_2_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_2_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[17]), 
        .QN(state2FF_state_gff_2_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_2_SFF_2_U5 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_2_SFF_2_n8), .A(state2FF_state_gff_2_SFF_2_n12), 
        .ZN(state2FF_state_gff_2_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_2_SFF_2_U4 ( .B1(state2FF_state_gff_2_SFF_2_n10), .B2(state2FF_inputPar[32]), .C1(state2FF_state_gff_2_SFF_2_n11), .C2(
        state2FF_inputPar[6]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_2_SFF_2_n12) );
  INV_X1 state2FF_state_gff_2_SFF_2_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_2_SFF_2_n11) );
  INV_X1 state2FF_state_gff_2_SFF_2_U2 ( .A(state2FF_state_gff_2_SFF_2_n11), 
        .ZN(state2FF_state_gff_2_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_2_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_2_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[33]), 
        .QN(state2FF_state_gff_2_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_2_SFF_3_U5 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_2_SFF_3_n8), .A(state2FF_state_gff_2_SFF_3_n12), 
        .ZN(state2FF_state_gff_2_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_2_SFF_3_U4 ( .B1(state2FF_state_gff_2_SFF_3_n10), .B2(state2FF_inputPar[48]), .C1(state2FF_state_gff_2_SFF_3_n11), .C2(
        state2FF_inputPar[7]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_2_SFF_3_n12) );
  INV_X1 state2FF_state_gff_2_SFF_3_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_2_SFF_3_n11) );
  INV_X1 state2FF_state_gff_2_SFF_3_U2 ( .A(state2FF_state_gff_2_SFF_3_n11), 
        .ZN(state2FF_state_gff_2_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_2_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_2_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[49]), 
        .QN(state2FF_state_gff_2_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_3_SFF_0_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_3_SFF_0_n8), .A(state2FF_state_gff_3_SFF_0_n12), 
        .ZN(state2FF_state_gff_3_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_3_SFF_0_U4 ( .B1(state2FF_state_gff_3_SFF_0_n10), .B2(state2FF_inputPar[1]), .C1(state2FF_state_gff_3_SFF_0_n11), .C2(
        state2FF_inputPar[8]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_3_SFF_0_n12) );
  INV_X1 state2FF_state_gff_3_SFF_0_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_3_SFF_0_n11) );
  INV_X1 state2FF_state_gff_3_SFF_0_U2 ( .A(state2FF_state_gff_3_SFF_0_n11), 
        .ZN(state2FF_state_gff_3_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_3_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_3_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[2]), 
        .QN(state2FF_state_gff_3_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_3_SFF_1_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_3_SFF_1_n8), .A(state2FF_state_gff_3_SFF_1_n12), 
        .ZN(state2FF_state_gff_3_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_3_SFF_1_U4 ( .B1(state2FF_state_gff_3_SFF_1_n10), .B2(state2FF_inputPar[17]), .C1(state2FF_state_gff_3_SFF_1_n11), .C2(
        state2FF_inputPar[9]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_3_SFF_1_n12) );
  INV_X1 state2FF_state_gff_3_SFF_1_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_3_SFF_1_n11) );
  INV_X1 state2FF_state_gff_3_SFF_1_U2 ( .A(state2FF_state_gff_3_SFF_1_n11), 
        .ZN(state2FF_state_gff_3_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_3_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_3_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[18]), 
        .QN(state2FF_state_gff_3_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_3_SFF_2_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_3_SFF_2_n7), .A(state2FF_state_gff_3_SFF_2_n11), 
        .ZN(state2FF_state_gff_3_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_3_SFF_2_U4 ( .B1(state2FF_state_gff_3_SFF_2_n9), 
        .B2(state2FF_inputPar[33]), .C1(state2FF_state_gff_3_SFF_2_n10), .C2(
        state2FF_inputPar[10]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_3_SFF_2_n11) );
  INV_X1 state2FF_state_gff_3_SFF_2_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_3_SFF_2_n10) );
  INV_X1 state2FF_state_gff_3_SFF_2_U2 ( .A(state2FF_state_gff_3_SFF_2_n10), 
        .ZN(state2FF_state_gff_3_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_3_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_3_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[34]), 
        .QN(state2FF_state_gff_3_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_3_SFF_3_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_3_SFF_3_n7), .A(state2FF_state_gff_3_SFF_3_n11), 
        .ZN(state2FF_state_gff_3_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_3_SFF_3_U4 ( .B1(state2FF_state_gff_3_SFF_3_n9), 
        .B2(state2FF_inputPar[49]), .C1(state2FF_state_gff_3_SFF_3_n10), .C2(
        state2FF_inputPar[11]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_3_SFF_3_n11) );
  INV_X1 state2FF_state_gff_3_SFF_3_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_3_SFF_3_n10) );
  INV_X1 state2FF_state_gff_3_SFF_3_U2 ( .A(state2FF_state_gff_3_SFF_3_n10), 
        .ZN(state2FF_state_gff_3_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_3_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_3_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[50]), 
        .QN(state2FF_state_gff_3_SFF_3_n7) );
  OAI21_X1 state2FF_state_gff_4_SFF_0_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_4_SFF_0_n7), .A(state2FF_state_gff_4_SFF_0_n11), 
        .ZN(state2FF_state_gff_4_SFF_0_n6) );
  OAI221_X1 state2FF_state_gff_4_SFF_0_U4 ( .B1(state2FF_state_gff_4_SFF_0_n9), 
        .B2(state2FF_inputPar[2]), .C1(state2FF_state_gff_4_SFF_0_n10), .C2(
        state2FF_inputPar[12]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_4_SFF_0_n11) );
  INV_X1 state2FF_state_gff_4_SFF_0_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_4_SFF_0_n10) );
  INV_X1 state2FF_state_gff_4_SFF_0_U2 ( .A(state2FF_state_gff_4_SFF_0_n10), 
        .ZN(state2FF_state_gff_4_SFF_0_n9) );
  DFF_X1 state2FF_state_gff_4_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_4_SFF_0_n6), .CK(clk), .Q(state2FF_inputPar[3]), 
        .QN(state2FF_state_gff_4_SFF_0_n7) );
  OAI21_X1 state2FF_state_gff_4_SFF_1_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_4_SFF_1_n7), .A(state2FF_state_gff_4_SFF_1_n11), 
        .ZN(state2FF_state_gff_4_SFF_1_n6) );
  OAI221_X1 state2FF_state_gff_4_SFF_1_U4 ( .B1(state2FF_state_gff_4_SFF_1_n9), 
        .B2(state2FF_inputPar[18]), .C1(state2FF_state_gff_4_SFF_1_n10), .C2(
        state2FF_inputPar[13]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_4_SFF_1_n11) );
  INV_X1 state2FF_state_gff_4_SFF_1_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_4_SFF_1_n10) );
  INV_X1 state2FF_state_gff_4_SFF_1_U2 ( .A(state2FF_state_gff_4_SFF_1_n10), 
        .ZN(state2FF_state_gff_4_SFF_1_n9) );
  DFF_X1 state2FF_state_gff_4_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_4_SFF_1_n6), .CK(clk), .Q(state2FF_inputPar[19]), 
        .QN(state2FF_state_gff_4_SFF_1_n7) );
  OAI21_X1 state2FF_state_gff_4_SFF_2_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_4_SFF_2_n7), .A(state2FF_state_gff_4_SFF_2_n11), 
        .ZN(state2FF_state_gff_4_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_4_SFF_2_U4 ( .B1(state2FF_state_gff_4_SFF_2_n9), 
        .B2(state2FF_inputPar[34]), .C1(state2FF_state_gff_4_SFF_2_n10), .C2(
        state2FF_inputPar[14]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_4_SFF_2_n11) );
  INV_X1 state2FF_state_gff_4_SFF_2_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_4_SFF_2_n10) );
  INV_X1 state2FF_state_gff_4_SFF_2_U2 ( .A(state2FF_state_gff_4_SFF_2_n10), 
        .ZN(state2FF_state_gff_4_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_4_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_4_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[35]), 
        .QN(state2FF_state_gff_4_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_4_SFF_3_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_4_SFF_3_n7), .A(state2FF_state_gff_4_SFF_3_n11), 
        .ZN(state2FF_state_gff_4_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_4_SFF_3_U4 ( .B1(state2FF_state_gff_4_SFF_3_n9), 
        .B2(state2FF_inputPar[50]), .C1(state2FF_state_gff_4_SFF_3_n10), .C2(
        state2FF_inputPar[15]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_4_SFF_3_n11) );
  INV_X1 state2FF_state_gff_4_SFF_3_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_4_SFF_3_n10) );
  INV_X1 state2FF_state_gff_4_SFF_3_U2 ( .A(state2FF_state_gff_4_SFF_3_n10), 
        .ZN(state2FF_state_gff_4_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_4_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_4_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[51]), 
        .QN(state2FF_state_gff_4_SFF_3_n7) );
  OAI21_X1 state2FF_state_gff_5_SFF_0_U5 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_5_SFF_0_n8), .A(state2FF_state_gff_5_SFF_0_n12), 
        .ZN(state2FF_state_gff_5_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_5_SFF_0_U4 ( .B1(state2FF_state_gff_5_SFF_0_n10), .B2(state2FF_inputPar[3]), .C1(state2FF_state_gff_5_SFF_0_n11), .C2(
        state2FF_inputPar[16]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_5_SFF_0_n12) );
  INV_X1 state2FF_state_gff_5_SFF_0_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_5_SFF_0_n11) );
  INV_X1 state2FF_state_gff_5_SFF_0_U2 ( .A(state2FF_state_gff_5_SFF_0_n11), 
        .ZN(state2FF_state_gff_5_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_5_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_5_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[4]), 
        .QN(state2FF_state_gff_5_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_5_SFF_1_U5 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_5_SFF_1_n8), .A(state2FF_state_gff_5_SFF_1_n12), 
        .ZN(state2FF_state_gff_5_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_5_SFF_1_U4 ( .B1(state2FF_state_gff_5_SFF_1_n10), .B2(state2FF_inputPar[19]), .C1(state2FF_state_gff_5_SFF_1_n11), .C2(
        state2FF_inputPar[17]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_5_SFF_1_n12) );
  INV_X1 state2FF_state_gff_5_SFF_1_U3 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_5_SFF_1_n11) );
  INV_X1 state2FF_state_gff_5_SFF_1_U2 ( .A(state2FF_state_gff_5_SFF_1_n11), 
        .ZN(state2FF_state_gff_5_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_5_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_5_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[20]), 
        .QN(state2FF_state_gff_5_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_5_SFF_2_U4 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_5_SFF_2_n8), .A(state2FF_state_gff_5_SFF_2_n11), 
        .ZN(state2FF_state_gff_5_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_5_SFF_2_U3 ( .B1(state2FF_state_n10), .B2(
        state2FF_inputPar[35]), .C1(state2FF_state_gff_5_SFF_2_n10), .C2(
        state2FF_inputPar[18]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_5_SFF_2_n11) );
  INV_X1 state2FF_state_gff_5_SFF_2_U2 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_5_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_5_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_5_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[36]), 
        .QN(state2FF_state_gff_5_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_5_SFF_3_U4 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_5_SFF_3_n8), .A(state2FF_state_gff_5_SFF_3_n11), 
        .ZN(state2FF_state_gff_5_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_5_SFF_3_U3 ( .B1(state2FF_state_n10), .B2(
        state2FF_inputPar[51]), .C1(state2FF_state_gff_5_SFF_3_n10), .C2(
        state2FF_inputPar[19]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_5_SFF_3_n11) );
  INV_X1 state2FF_state_gff_5_SFF_3_U2 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_5_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_5_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_5_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[52]), 
        .QN(state2FF_state_gff_5_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_6_SFF_0_U4 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_6_SFF_0_n8), .A(state2FF_state_gff_6_SFF_0_n11), 
        .ZN(state2FF_state_gff_6_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_6_SFF_0_U3 ( .B1(state2FF_state_n10), .B2(
        state2FF_inputPar[4]), .C1(state2FF_state_gff_6_SFF_0_n10), .C2(
        state2FF_inputPar[20]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_6_SFF_0_n11) );
  INV_X1 state2FF_state_gff_6_SFF_0_U2 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_6_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_6_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_6_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[5]), 
        .QN(state2FF_state_gff_6_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_6_SFF_1_U4 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_6_SFF_1_n8), .A(state2FF_state_gff_6_SFF_1_n11), 
        .ZN(state2FF_state_gff_6_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_6_SFF_1_U3 ( .B1(state2FF_state_n10), .B2(
        state2FF_inputPar[20]), .C1(state2FF_state_gff_6_SFF_1_n10), .C2(
        state2FF_inputPar[21]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_6_SFF_1_n11) );
  INV_X1 state2FF_state_gff_6_SFF_1_U2 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_6_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_6_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_6_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[21]), 
        .QN(state2FF_state_gff_6_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_6_SFF_2_U4 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_6_SFF_2_n8), .A(state2FF_state_gff_6_SFF_2_n11), 
        .ZN(state2FF_state_gff_6_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_6_SFF_2_U3 ( .B1(state2FF_state_n10), .B2(
        state2FF_inputPar[36]), .C1(state2FF_state_gff_6_SFF_2_n10), .C2(
        state2FF_inputPar[22]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_6_SFF_2_n11) );
  INV_X1 state2FF_state_gff_6_SFF_2_U2 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_6_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_6_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_6_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[37]), 
        .QN(state2FF_state_gff_6_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_6_SFF_3_U4 ( .B1(state2FF_state_n8), .B2(
        state2FF_state_gff_6_SFF_3_n8), .A(state2FF_state_gff_6_SFF_3_n11), 
        .ZN(state2FF_state_gff_6_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_6_SFF_3_U3 ( .B1(state2FF_state_n10), .B2(
        state2FF_inputPar[52]), .C1(state2FF_state_gff_6_SFF_3_n10), .C2(
        state2FF_inputPar[23]), .A(state2FF_state_n8), .ZN(
        state2FF_state_gff_6_SFF_3_n11) );
  INV_X1 state2FF_state_gff_6_SFF_3_U2 ( .A(state2FF_state_n10), .ZN(
        state2FF_state_gff_6_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_6_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_6_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[53]), 
        .QN(state2FF_state_gff_6_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_7_SFF_0_U4 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_7_SFF_0_n8), .A(state2FF_state_gff_7_SFF_0_n11), 
        .ZN(state2FF_state_gff_7_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_7_SFF_0_U3 ( .B1(state2FF_state_n12), .B2(
        state2FF_inputPar[5]), .C1(state2FF_state_gff_7_SFF_0_n10), .C2(
        state2FF_inputPar[24]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_7_SFF_0_n11) );
  INV_X1 state2FF_state_gff_7_SFF_0_U2 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_7_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_7_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_7_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[6]), 
        .QN(state2FF_state_gff_7_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_7_SFF_1_U4 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_7_SFF_1_n8), .A(state2FF_state_gff_7_SFF_1_n11), 
        .ZN(state2FF_state_gff_7_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_7_SFF_1_U3 ( .B1(state2FF_state_n12), .B2(
        state2FF_inputPar[21]), .C1(state2FF_state_gff_7_SFF_1_n10), .C2(
        state2FF_inputPar[25]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_7_SFF_1_n11) );
  INV_X1 state2FF_state_gff_7_SFF_1_U2 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_7_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_7_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_7_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[22]), 
        .QN(state2FF_state_gff_7_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_7_SFF_2_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_7_SFF_2_n7), .A(state2FF_state_gff_7_SFF_2_n11), 
        .ZN(state2FF_state_gff_7_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_7_SFF_2_U4 ( .B1(state2FF_state_gff_7_SFF_2_n9), 
        .B2(state2FF_inputPar[37]), .C1(state2FF_state_gff_7_SFF_2_n10), .C2(
        state2FF_inputPar[26]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_7_SFF_2_n11) );
  INV_X1 state2FF_state_gff_7_SFF_2_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_7_SFF_2_n10) );
  INV_X1 state2FF_state_gff_7_SFF_2_U2 ( .A(state2FF_state_gff_7_SFF_2_n10), 
        .ZN(state2FF_state_gff_7_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_7_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_7_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[38]), 
        .QN(state2FF_state_gff_7_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_7_SFF_3_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_7_SFF_3_n7), .A(state2FF_state_gff_7_SFF_3_n11), 
        .ZN(state2FF_state_gff_7_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_7_SFF_3_U4 ( .B1(state2FF_state_gff_7_SFF_3_n9), 
        .B2(state2FF_inputPar[53]), .C1(state2FF_state_gff_7_SFF_3_n10), .C2(
        state2FF_inputPar[27]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_7_SFF_3_n11) );
  INV_X1 state2FF_state_gff_7_SFF_3_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_7_SFF_3_n10) );
  INV_X1 state2FF_state_gff_7_SFF_3_U2 ( .A(state2FF_state_gff_7_SFF_3_n10), 
        .ZN(state2FF_state_gff_7_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_7_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_7_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[54]), 
        .QN(state2FF_state_gff_7_SFF_3_n7) );
  OAI21_X1 state2FF_state_gff_8_SFF_0_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_8_SFF_0_n7), .A(state2FF_state_gff_8_SFF_0_n11), 
        .ZN(state2FF_state_gff_8_SFF_0_n6) );
  OAI221_X1 state2FF_state_gff_8_SFF_0_U4 ( .B1(state2FF_state_gff_8_SFF_0_n9), 
        .B2(state2FF_inputPar[6]), .C1(state2FF_state_gff_8_SFF_0_n10), .C2(
        state2FF_inputPar[28]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_8_SFF_0_n11) );
  INV_X1 state2FF_state_gff_8_SFF_0_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_8_SFF_0_n10) );
  INV_X1 state2FF_state_gff_8_SFF_0_U2 ( .A(state2FF_state_gff_8_SFF_0_n10), 
        .ZN(state2FF_state_gff_8_SFF_0_n9) );
  DFF_X1 state2FF_state_gff_8_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_8_SFF_0_n6), .CK(clk), .Q(state2FF_inputPar[7]), 
        .QN(state2FF_state_gff_8_SFF_0_n7) );
  OAI21_X1 state2FF_state_gff_8_SFF_1_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_8_SFF_1_n7), .A(state2FF_state_gff_8_SFF_1_n11), 
        .ZN(state2FF_state_gff_8_SFF_1_n6) );
  OAI221_X1 state2FF_state_gff_8_SFF_1_U4 ( .B1(state2FF_state_gff_8_SFF_1_n9), 
        .B2(state2FF_inputPar[22]), .C1(state2FF_state_gff_8_SFF_1_n10), .C2(
        state2FF_inputPar[29]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_8_SFF_1_n11) );
  INV_X1 state2FF_state_gff_8_SFF_1_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_8_SFF_1_n10) );
  INV_X1 state2FF_state_gff_8_SFF_1_U2 ( .A(state2FF_state_gff_8_SFF_1_n10), 
        .ZN(state2FF_state_gff_8_SFF_1_n9) );
  DFF_X1 state2FF_state_gff_8_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_8_SFF_1_n6), .CK(clk), .Q(state2FF_inputPar[23]), 
        .QN(state2FF_state_gff_8_SFF_1_n7) );
  OAI21_X1 state2FF_state_gff_8_SFF_2_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_8_SFF_2_n7), .A(state2FF_state_gff_8_SFF_2_n11), 
        .ZN(state2FF_state_gff_8_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_8_SFF_2_U4 ( .B1(state2FF_state_gff_8_SFF_2_n9), 
        .B2(state2FF_inputPar[38]), .C1(state2FF_state_gff_8_SFF_2_n10), .C2(
        state2FF_inputPar[30]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_8_SFF_2_n11) );
  INV_X1 state2FF_state_gff_8_SFF_2_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_8_SFF_2_n10) );
  INV_X1 state2FF_state_gff_8_SFF_2_U2 ( .A(state2FF_state_gff_8_SFF_2_n10), 
        .ZN(state2FF_state_gff_8_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_8_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_8_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[39]), 
        .QN(state2FF_state_gff_8_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_8_SFF_3_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_8_SFF_3_n7), .A(state2FF_state_gff_8_SFF_3_n11), 
        .ZN(state2FF_state_gff_8_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_8_SFF_3_U4 ( .B1(state2FF_state_gff_8_SFF_3_n9), 
        .B2(state2FF_inputPar[54]), .C1(state2FF_state_gff_8_SFF_3_n10), .C2(
        state2FF_inputPar[31]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_8_SFF_3_n11) );
  INV_X1 state2FF_state_gff_8_SFF_3_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_8_SFF_3_n10) );
  INV_X1 state2FF_state_gff_8_SFF_3_U2 ( .A(state2FF_state_gff_8_SFF_3_n10), 
        .ZN(state2FF_state_gff_8_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_8_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_8_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[55]), 
        .QN(state2FF_state_gff_8_SFF_3_n7) );
  OAI21_X1 state2FF_state_gff_9_SFF_0_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_9_SFF_0_n8), .A(state2FF_state_gff_9_SFF_0_n12), 
        .ZN(state2FF_state_gff_9_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_9_SFF_0_U4 ( .B1(state2FF_state_gff_9_SFF_0_n10), .B2(state2FF_inputPar[7]), .C1(state2FF_state_gff_9_SFF_0_n11), .C2(
        state2FF_inputPar[32]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_9_SFF_0_n12) );
  INV_X1 state2FF_state_gff_9_SFF_0_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_9_SFF_0_n11) );
  INV_X1 state2FF_state_gff_9_SFF_0_U2 ( .A(state2FF_state_gff_9_SFF_0_n11), 
        .ZN(state2FF_state_gff_9_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_9_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_9_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[8]), 
        .QN(state2FF_state_gff_9_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_9_SFF_1_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_9_SFF_1_n8), .A(state2FF_state_gff_9_SFF_1_n12), 
        .ZN(state2FF_state_gff_9_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_9_SFF_1_U4 ( .B1(state2FF_state_gff_9_SFF_1_n10), .B2(state2FF_inputPar[23]), .C1(state2FF_state_gff_9_SFF_1_n11), .C2(
        state2FF_inputPar[33]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_9_SFF_1_n12) );
  INV_X1 state2FF_state_gff_9_SFF_1_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_9_SFF_1_n11) );
  INV_X1 state2FF_state_gff_9_SFF_1_U2 ( .A(state2FF_state_gff_9_SFF_1_n11), 
        .ZN(state2FF_state_gff_9_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_9_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_9_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[24]), 
        .QN(state2FF_state_gff_9_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_9_SFF_2_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_9_SFF_2_n8), .A(state2FF_state_gff_9_SFF_2_n12), 
        .ZN(state2FF_state_gff_9_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_9_SFF_2_U4 ( .B1(state2FF_state_gff_9_SFF_2_n10), .B2(state2FF_inputPar[39]), .C1(state2FF_state_gff_9_SFF_2_n11), .C2(
        state2FF_inputPar[34]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_9_SFF_2_n12) );
  INV_X1 state2FF_state_gff_9_SFF_2_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_9_SFF_2_n11) );
  INV_X1 state2FF_state_gff_9_SFF_2_U2 ( .A(state2FF_state_gff_9_SFF_2_n11), 
        .ZN(state2FF_state_gff_9_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_9_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_9_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[40]), 
        .QN(state2FF_state_gff_9_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_9_SFF_3_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_9_SFF_3_n8), .A(state2FF_state_gff_9_SFF_3_n12), 
        .ZN(state2FF_state_gff_9_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_9_SFF_3_U4 ( .B1(state2FF_state_gff_9_SFF_3_n10), .B2(state2FF_inputPar[55]), .C1(state2FF_state_gff_9_SFF_3_n11), .C2(
        state2FF_inputPar[35]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_9_SFF_3_n12) );
  INV_X1 state2FF_state_gff_9_SFF_3_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_9_SFF_3_n11) );
  INV_X1 state2FF_state_gff_9_SFF_3_U2 ( .A(state2FF_state_gff_9_SFF_3_n11), 
        .ZN(state2FF_state_gff_9_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_9_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_9_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[56]), 
        .QN(state2FF_state_gff_9_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_10_SFF_0_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_10_SFF_0_n8), .A(state2FF_state_gff_10_SFF_0_n12), 
        .ZN(state2FF_state_gff_10_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_10_SFF_0_U4 ( .B1(
        state2FF_state_gff_10_SFF_0_n10), .B2(state2FF_inputPar[8]), .C1(
        state2FF_state_gff_10_SFF_0_n11), .C2(state2FF_inputPar[36]), .A(
        state2FF_state_n7), .ZN(state2FF_state_gff_10_SFF_0_n12) );
  INV_X1 state2FF_state_gff_10_SFF_0_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_10_SFF_0_n11) );
  INV_X1 state2FF_state_gff_10_SFF_0_U2 ( .A(state2FF_state_gff_10_SFF_0_n11), 
        .ZN(state2FF_state_gff_10_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_10_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_10_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[9]), 
        .QN(state2FF_state_gff_10_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_10_SFF_1_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_10_SFF_1_n8), .A(state2FF_state_gff_10_SFF_1_n12), 
        .ZN(state2FF_state_gff_10_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_10_SFF_1_U4 ( .B1(
        state2FF_state_gff_10_SFF_1_n10), .B2(state2FF_inputPar[24]), .C1(
        state2FF_state_gff_10_SFF_1_n11), .C2(state2FF_inputPar[37]), .A(
        state2FF_state_n7), .ZN(state2FF_state_gff_10_SFF_1_n12) );
  INV_X1 state2FF_state_gff_10_SFF_1_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_10_SFF_1_n11) );
  INV_X1 state2FF_state_gff_10_SFF_1_U2 ( .A(state2FF_state_gff_10_SFF_1_n11), 
        .ZN(state2FF_state_gff_10_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_10_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_10_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[25]), 
        .QN(state2FF_state_gff_10_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_10_SFF_2_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_10_SFF_2_n8), .A(state2FF_state_gff_10_SFF_2_n12), 
        .ZN(state2FF_state_gff_10_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_10_SFF_2_U4 ( .B1(
        state2FF_state_gff_10_SFF_2_n10), .B2(state2FF_inputPar[40]), .C1(
        state2FF_state_gff_10_SFF_2_n11), .C2(state2FF_inputPar[38]), .A(
        state2FF_state_n7), .ZN(state2FF_state_gff_10_SFF_2_n12) );
  INV_X1 state2FF_state_gff_10_SFF_2_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_10_SFF_2_n11) );
  INV_X1 state2FF_state_gff_10_SFF_2_U2 ( .A(state2FF_state_gff_10_SFF_2_n11), 
        .ZN(state2FF_state_gff_10_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_10_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_10_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[41]), 
        .QN(state2FF_state_gff_10_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_10_SFF_3_U5 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_10_SFF_3_n8), .A(state2FF_state_gff_10_SFF_3_n12), 
        .ZN(state2FF_state_gff_10_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_10_SFF_3_U4 ( .B1(
        state2FF_state_gff_10_SFF_3_n10), .B2(state2FF_inputPar[56]), .C1(
        state2FF_state_gff_10_SFF_3_n11), .C2(state2FF_inputPar[39]), .A(
        state2FF_state_n7), .ZN(state2FF_state_gff_10_SFF_3_n12) );
  INV_X1 state2FF_state_gff_10_SFF_3_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_10_SFF_3_n11) );
  INV_X1 state2FF_state_gff_10_SFF_3_U2 ( .A(state2FF_state_gff_10_SFF_3_n11), 
        .ZN(state2FF_state_gff_10_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_10_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_10_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[57]), 
        .QN(state2FF_state_gff_10_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_11_SFF_0_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_11_SFF_0_n8), .A(state2FF_state_gff_11_SFF_0_n11), 
        .ZN(state2FF_state_gff_11_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_11_SFF_0_U3 ( .B1(state2FF_state_n12), .B2(
        state2FF_inputPar[9]), .C1(state2FF_state_gff_11_SFF_0_n10), .C2(
        state2FF_inputPar[40]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_11_SFF_0_n11) );
  INV_X1 state2FF_state_gff_11_SFF_0_U2 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_11_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_11_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_11_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[10]), 
        .QN(state2FF_state_gff_11_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_11_SFF_1_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_11_SFF_1_n8), .A(state2FF_state_gff_11_SFF_1_n11), 
        .ZN(state2FF_state_gff_11_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_11_SFF_1_U3 ( .B1(state2FF_state_n12), .B2(
        state2FF_inputPar[25]), .C1(state2FF_state_gff_11_SFF_1_n10), .C2(
        state2FF_inputPar[41]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_11_SFF_1_n11) );
  INV_X1 state2FF_state_gff_11_SFF_1_U2 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_11_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_11_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_11_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[26]), 
        .QN(state2FF_state_gff_11_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_11_SFF_2_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_11_SFF_2_n7), .A(state2FF_state_gff_11_SFF_2_n11), 
        .ZN(state2FF_state_gff_11_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_11_SFF_2_U4 ( .B1(
        state2FF_state_gff_11_SFF_2_n9), .B2(state2FF_inputPar[41]), .C1(
        state2FF_state_gff_11_SFF_2_n10), .C2(state2FF_inputPar[42]), .A(
        state2FF_state_n9), .ZN(state2FF_state_gff_11_SFF_2_n11) );
  INV_X1 state2FF_state_gff_11_SFF_2_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_11_SFF_2_n10) );
  INV_X1 state2FF_state_gff_11_SFF_2_U2 ( .A(state2FF_state_gff_11_SFF_2_n10), 
        .ZN(state2FF_state_gff_11_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_11_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_11_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[42]), 
        .QN(state2FF_state_gff_11_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_11_SFF_3_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_11_SFF_3_n7), .A(state2FF_state_gff_11_SFF_3_n11), 
        .ZN(state2FF_state_gff_11_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_11_SFF_3_U4 ( .B1(
        state2FF_state_gff_11_SFF_3_n9), .B2(state2FF_inputPar[57]), .C1(
        state2FF_state_gff_11_SFF_3_n10), .C2(state2FF_inputPar[43]), .A(
        state2FF_state_n9), .ZN(state2FF_state_gff_11_SFF_3_n11) );
  INV_X1 state2FF_state_gff_11_SFF_3_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_11_SFF_3_n10) );
  INV_X1 state2FF_state_gff_11_SFF_3_U2 ( .A(state2FF_state_gff_11_SFF_3_n10), 
        .ZN(state2FF_state_gff_11_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_11_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_11_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[58]), 
        .QN(state2FF_state_gff_11_SFF_3_n7) );
  OAI21_X1 state2FF_state_gff_12_SFF_0_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_12_SFF_0_n7), .A(state2FF_state_gff_12_SFF_0_n11), 
        .ZN(state2FF_state_gff_12_SFF_0_n6) );
  OAI221_X1 state2FF_state_gff_12_SFF_0_U4 ( .B1(
        state2FF_state_gff_12_SFF_0_n9), .B2(state2FF_inputPar[10]), .C1(
        state2FF_state_gff_12_SFF_0_n10), .C2(state2FF_inputPar[44]), .A(
        state2FF_state_n6), .ZN(state2FF_state_gff_12_SFF_0_n11) );
  INV_X1 state2FF_state_gff_12_SFF_0_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_12_SFF_0_n10) );
  INV_X1 state2FF_state_gff_12_SFF_0_U2 ( .A(state2FF_state_gff_12_SFF_0_n10), 
        .ZN(state2FF_state_gff_12_SFF_0_n9) );
  DFF_X1 state2FF_state_gff_12_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_12_SFF_0_n6), .CK(clk), .Q(state2FF_inputPar[11]), 
        .QN(state2FF_state_gff_12_SFF_0_n7) );
  OAI21_X1 state2FF_state_gff_12_SFF_1_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_12_SFF_1_n7), .A(state2FF_state_gff_12_SFF_1_n11), 
        .ZN(state2FF_state_gff_12_SFF_1_n6) );
  OAI221_X1 state2FF_state_gff_12_SFF_1_U4 ( .B1(
        state2FF_state_gff_12_SFF_1_n9), .B2(state2FF_inputPar[26]), .C1(
        state2FF_state_gff_12_SFF_1_n10), .C2(state2FF_inputPar[45]), .A(
        state2FF_state_n6), .ZN(state2FF_state_gff_12_SFF_1_n11) );
  INV_X1 state2FF_state_gff_12_SFF_1_U3 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_12_SFF_1_n10) );
  INV_X1 state2FF_state_gff_12_SFF_1_U2 ( .A(state2FF_state_gff_12_SFF_1_n10), 
        .ZN(state2FF_state_gff_12_SFF_1_n9) );
  DFF_X1 state2FF_state_gff_12_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_12_SFF_1_n6), .CK(clk), .Q(state2FF_inputPar[27]), 
        .QN(state2FF_state_gff_12_SFF_1_n7) );
  OAI21_X1 state2FF_state_gff_12_SFF_2_U4 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_12_SFF_2_n7), .A(state2FF_state_gff_12_SFF_2_n10), 
        .ZN(state2FF_state_gff_12_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_12_SFF_2_U3 ( .B1(state2FF_state_n13), .B2(
        state2FF_inputPar[42]), .C1(state2FF_state_gff_12_SFF_2_n9), .C2(
        state2FF_inputPar[46]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_12_SFF_2_n10) );
  INV_X1 state2FF_state_gff_12_SFF_2_U2 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_12_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_12_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_12_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[43]), 
        .QN(state2FF_state_gff_12_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_12_SFF_3_U4 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_12_SFF_3_n7), .A(state2FF_state_gff_12_SFF_3_n10), 
        .ZN(state2FF_state_gff_12_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_12_SFF_3_U3 ( .B1(state2FF_state_n13), .B2(
        state2FF_inputPar[58]), .C1(state2FF_state_gff_12_SFF_3_n9), .C2(
        state2FF_inputPar[47]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_12_SFF_3_n10) );
  INV_X1 state2FF_state_gff_12_SFF_3_U2 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_12_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_12_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_12_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[59]), 
        .QN(state2FF_state_gff_12_SFF_3_n7) );
  OAI21_X1 state2FF_state_gff_13_SFF_0_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_13_SFF_0_n8), .A(state2FF_state_gff_13_SFF_0_n12), 
        .ZN(state2FF_state_gff_13_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_13_SFF_0_U4 ( .B1(
        state2FF_state_gff_13_SFF_0_n10), .B2(state2FF_inputPar[11]), .C1(
        state2FF_state_gff_13_SFF_0_n11), .C2(state2FF_inputPar[48]), .A(
        state2FF_state_n6), .ZN(state2FF_state_gff_13_SFF_0_n12) );
  INV_X1 state2FF_state_gff_13_SFF_0_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_13_SFF_0_n11) );
  INV_X1 state2FF_state_gff_13_SFF_0_U2 ( .A(state2FF_state_gff_13_SFF_0_n11), 
        .ZN(state2FF_state_gff_13_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_13_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_13_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[12]), 
        .QN(state2FF_state_gff_13_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_13_SFF_1_U5 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_13_SFF_1_n8), .A(state2FF_state_gff_13_SFF_1_n12), 
        .ZN(state2FF_state_gff_13_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_13_SFF_1_U4 ( .B1(
        state2FF_state_gff_13_SFF_1_n10), .B2(state2FF_inputPar[27]), .C1(
        state2FF_state_gff_13_SFF_1_n11), .C2(state2FF_inputPar[49]), .A(
        state2FF_state_n6), .ZN(state2FF_state_gff_13_SFF_1_n12) );
  INV_X1 state2FF_state_gff_13_SFF_1_U3 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_13_SFF_1_n11) );
  INV_X1 state2FF_state_gff_13_SFF_1_U2 ( .A(state2FF_state_gff_13_SFF_1_n11), 
        .ZN(state2FF_state_gff_13_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_13_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_13_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[28]), 
        .QN(state2FF_state_gff_13_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_13_SFF_2_U4 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_13_SFF_2_n8), .A(state2FF_state_gff_13_SFF_2_n11), 
        .ZN(state2FF_state_gff_13_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_13_SFF_2_U3 ( .B1(state2FF_state_n11), .B2(
        state2FF_inputPar[43]), .C1(state2FF_state_gff_13_SFF_2_n10), .C2(
        state2FF_inputPar[50]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_13_SFF_2_n11) );
  INV_X1 state2FF_state_gff_13_SFF_2_U2 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_13_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_13_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_13_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[44]), 
        .QN(state2FF_state_gff_13_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_13_SFF_3_U4 ( .B1(state2FF_state_n6), .B2(
        state2FF_state_gff_13_SFF_3_n8), .A(state2FF_state_gff_13_SFF_3_n11), 
        .ZN(state2FF_state_gff_13_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_13_SFF_3_U3 ( .B1(state2FF_state_n11), .B2(
        state2FF_inputPar[59]), .C1(state2FF_state_gff_13_SFF_3_n10), .C2(
        state2FF_inputPar[51]), .A(state2FF_state_n6), .ZN(
        state2FF_state_gff_13_SFF_3_n11) );
  INV_X1 state2FF_state_gff_13_SFF_3_U2 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_13_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_13_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_13_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[60]), 
        .QN(state2FF_state_gff_13_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_14_SFF_0_U4 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_14_SFF_0_n8), .A(state2FF_state_gff_14_SFF_0_n11), 
        .ZN(state2FF_state_gff_14_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_14_SFF_0_U3 ( .B1(state2FF_state_n11), .B2(
        state2FF_inputPar[12]), .C1(state2FF_state_gff_14_SFF_0_n10), .C2(
        state2FF_inputPar[52]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_14_SFF_0_n11) );
  INV_X1 state2FF_state_gff_14_SFF_0_U2 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_14_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_14_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_14_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[13]), 
        .QN(state2FF_state_gff_14_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_14_SFF_1_U4 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_14_SFF_1_n8), .A(state2FF_state_gff_14_SFF_1_n11), 
        .ZN(state2FF_state_gff_14_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_14_SFF_1_U3 ( .B1(state2FF_state_n11), .B2(
        state2FF_inputPar[28]), .C1(state2FF_state_gff_14_SFF_1_n10), .C2(
        state2FF_inputPar[53]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_14_SFF_1_n11) );
  INV_X1 state2FF_state_gff_14_SFF_1_U2 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_14_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_14_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_14_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[29]), 
        .QN(state2FF_state_gff_14_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_14_SFF_2_U4 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_14_SFF_2_n8), .A(state2FF_state_gff_14_SFF_2_n11), 
        .ZN(state2FF_state_gff_14_SFF_2_n7) );
  OAI221_X1 state2FF_state_gff_14_SFF_2_U3 ( .B1(state2FF_state_n11), .B2(
        state2FF_inputPar[44]), .C1(state2FF_state_gff_14_SFF_2_n10), .C2(
        state2FF_inputPar[54]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_14_SFF_2_n11) );
  INV_X1 state2FF_state_gff_14_SFF_2_U2 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_14_SFF_2_n10) );
  DFF_X1 state2FF_state_gff_14_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_14_SFF_2_n7), .CK(clk), .Q(state2FF_inputPar[45]), 
        .QN(state2FF_state_gff_14_SFF_2_n8) );
  OAI21_X1 state2FF_state_gff_14_SFF_3_U4 ( .B1(state2FF_state_n7), .B2(
        state2FF_state_gff_14_SFF_3_n8), .A(state2FF_state_gff_14_SFF_3_n11), 
        .ZN(state2FF_state_gff_14_SFF_3_n7) );
  OAI221_X1 state2FF_state_gff_14_SFF_3_U3 ( .B1(state2FF_state_n11), .B2(
        state2FF_inputPar[60]), .C1(state2FF_state_gff_14_SFF_3_n10), .C2(
        state2FF_inputPar[55]), .A(state2FF_state_n7), .ZN(
        state2FF_state_gff_14_SFF_3_n11) );
  INV_X1 state2FF_state_gff_14_SFF_3_U2 ( .A(state2FF_state_n11), .ZN(
        state2FF_state_gff_14_SFF_3_n10) );
  DFF_X1 state2FF_state_gff_14_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_14_SFF_3_n7), .CK(clk), .Q(state2FF_inputPar[61]), 
        .QN(state2FF_state_gff_14_SFF_3_n8) );
  OAI21_X1 state2FF_state_gff_15_SFF_0_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_15_SFF_0_n8), .A(state2FF_state_gff_15_SFF_0_n11), 
        .ZN(state2FF_state_gff_15_SFF_0_n7) );
  OAI221_X1 state2FF_state_gff_15_SFF_0_U3 ( .B1(state2FF_state_n12), .B2(
        state2FF_inputPar[13]), .C1(state2FF_state_gff_15_SFF_0_n10), .C2(
        state2FF_inputPar[56]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_15_SFF_0_n11) );
  INV_X1 state2FF_state_gff_15_SFF_0_U2 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_15_SFF_0_n10) );
  DFF_X1 state2FF_state_gff_15_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_15_SFF_0_n7), .CK(clk), .Q(state2FF_inputPar[14]), 
        .QN(state2FF_state_gff_15_SFF_0_n8) );
  OAI21_X1 state2FF_state_gff_15_SFF_1_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_15_SFF_1_n8), .A(state2FF_state_gff_15_SFF_1_n11), 
        .ZN(state2FF_state_gff_15_SFF_1_n7) );
  OAI221_X1 state2FF_state_gff_15_SFF_1_U3 ( .B1(state2FF_state_n12), .B2(
        state2FF_inputPar[29]), .C1(state2FF_state_gff_15_SFF_1_n10), .C2(
        state2FF_inputPar[57]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_15_SFF_1_n11) );
  INV_X1 state2FF_state_gff_15_SFF_1_U2 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_15_SFF_1_n10) );
  DFF_X1 state2FF_state_gff_15_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_15_SFF_1_n7), .CK(clk), .Q(state2FF_inputPar[30]), 
        .QN(state2FF_state_gff_15_SFF_1_n8) );
  OAI21_X1 state2FF_state_gff_15_SFF_2_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_15_SFF_2_n7), .A(state2FF_state_gff_15_SFF_2_n11), 
        .ZN(state2FF_state_gff_15_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_15_SFF_2_U4 ( .B1(
        state2FF_state_gff_15_SFF_2_n9), .B2(state2FF_inputPar[45]), .C1(
        state2FF_state_gff_15_SFF_2_n10), .C2(state2FF_inputPar[58]), .A(
        state2FF_state_n9), .ZN(state2FF_state_gff_15_SFF_2_n11) );
  INV_X1 state2FF_state_gff_15_SFF_2_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_15_SFF_2_n10) );
  INV_X1 state2FF_state_gff_15_SFF_2_U2 ( .A(state2FF_state_gff_15_SFF_2_n10), 
        .ZN(state2FF_state_gff_15_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_15_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_15_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[46]), 
        .QN(state2FF_state_gff_15_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_15_SFF_3_U5 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_15_SFF_3_n7), .A(state2FF_state_gff_15_SFF_3_n11), 
        .ZN(state2FF_state_gff_15_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_15_SFF_3_U4 ( .B1(
        state2FF_state_gff_15_SFF_3_n9), .B2(state2FF_inputPar[61]), .C1(
        state2FF_state_gff_15_SFF_3_n10), .C2(state2FF_inputPar[59]), .A(
        state2FF_state_n9), .ZN(state2FF_state_gff_15_SFF_3_n11) );
  INV_X1 state2FF_state_gff_15_SFF_3_U3 ( .A(state2FF_state_n12), .ZN(
        state2FF_state_gff_15_SFF_3_n10) );
  INV_X1 state2FF_state_gff_15_SFF_3_U2 ( .A(state2FF_state_gff_15_SFF_3_n10), 
        .ZN(state2FF_state_gff_15_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_15_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_15_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[62]), 
        .QN(state2FF_state_gff_15_SFF_3_n7) );
  OAI21_X1 state2FF_state_gff_16_SFF_0_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_16_SFF_0_n7), .A(state2FF_state_gff_16_SFF_0_n10), 
        .ZN(state2FF_state_gff_16_SFF_0_n6) );
  OAI221_X1 state2FF_state_gff_16_SFF_0_U3 ( .B1(state2FF_state_n13), .B2(
        state2FF_inputPar[14]), .C1(state2FF_state_gff_16_SFF_0_n9), .C2(
        state2FF_inputPar[60]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_16_SFF_0_n10) );
  INV_X1 state2FF_state_gff_16_SFF_0_U2 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_16_SFF_0_n9) );
  DFF_X1 state2FF_state_gff_16_SFF_0_Cell_reg ( .D(
        state2FF_state_gff_16_SFF_0_n6), .CK(clk), .Q(state2FF_inputPar[15]), 
        .QN(state2FF_state_gff_16_SFF_0_n7) );
  OAI21_X1 state2FF_state_gff_16_SFF_1_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_16_SFF_1_n7), .A(state2FF_state_gff_16_SFF_1_n10), 
        .ZN(state2FF_state_gff_16_SFF_1_n6) );
  OAI221_X1 state2FF_state_gff_16_SFF_1_U3 ( .B1(state2FF_state_n13), .B2(
        state2FF_inputPar[30]), .C1(state2FF_state_gff_16_SFF_1_n9), .C2(
        state2FF_inputPar[61]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_16_SFF_1_n10) );
  INV_X1 state2FF_state_gff_16_SFF_1_U2 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_16_SFF_1_n9) );
  DFF_X1 state2FF_state_gff_16_SFF_1_Cell_reg ( .D(
        state2FF_state_gff_16_SFF_1_n6), .CK(clk), .Q(state2FF_inputPar[31]), 
        .QN(state2FF_state_gff_16_SFF_1_n7) );
  OAI21_X1 state2FF_state_gff_16_SFF_2_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_16_SFF_2_n7), .A(state2FF_state_gff_16_SFF_2_n10), 
        .ZN(state2FF_state_gff_16_SFF_2_n6) );
  OAI221_X1 state2FF_state_gff_16_SFF_2_U3 ( .B1(state2FF_state_n13), .B2(
        state2FF_inputPar[46]), .C1(state2FF_state_gff_16_SFF_2_n9), .C2(
        state2FF_inputPar[62]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_16_SFF_2_n10) );
  INV_X1 state2FF_state_gff_16_SFF_2_U2 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_16_SFF_2_n9) );
  DFF_X1 state2FF_state_gff_16_SFF_2_Cell_reg ( .D(
        state2FF_state_gff_16_SFF_2_n6), .CK(clk), .Q(state2FF_inputPar[47]), 
        .QN(state2FF_state_gff_16_SFF_2_n7) );
  OAI21_X1 state2FF_state_gff_16_SFF_3_U4 ( .B1(state2FF_state_n9), .B2(
        state2FF_state_gff_16_SFF_3_n7), .A(state2FF_state_gff_16_SFF_3_n10), 
        .ZN(state2FF_state_gff_16_SFF_3_n6) );
  OAI221_X1 state2FF_state_gff_16_SFF_3_U3 ( .B1(state2FF_state_n13), .B2(
        state2FF_inputPar[62]), .C1(state2FF_state_gff_16_SFF_3_n9), .C2(
        state2FF_inputPar[63]), .A(state2FF_state_n9), .ZN(
        state2FF_state_gff_16_SFF_3_n10) );
  INV_X1 state2FF_state_gff_16_SFF_3_U2 ( .A(state2FF_state_n13), .ZN(
        state2FF_state_gff_16_SFF_3_n9) );
  DFF_X1 state2FF_state_gff_16_SFF_3_Cell_reg ( .D(
        state2FF_state_gff_16_SFF_3_n6), .CK(clk), .Q(state2FF_inputPar[63]), 
        .QN(state2FF_state_gff_16_SFF_3_n7) );
  MUX2_X1 state3FF_U5 ( .A(sboxOut3[2]), .B(dataIn3[2]), .S(n4), .Z(
        state3FF_n1) );
  MUX2_X1 state3FF_U4 ( .A(sboxOut3[1]), .B(dataIn3[1]), .S(n4), .Z(
        state3FF_n2) );
  MUX2_X1 state3FF_U3 ( .A(sboxOut3[0]), .B(dataIn3[0]), .S(n4), .Z(
        state3FF_n3) );
  MUX2_X1 state3FF_U2 ( .A(sboxOut3[3]), .B(dataIn3[3]), .S(n4), .Z(
        state3FF_n4) );
  BUF_X2 state3FF_state_U7 ( .A(enData), .Z(state3FF_state_n7) );
  BUF_X2 state3FF_state_U6 ( .A(enData), .Z(state3FF_state_n8) );
  BUF_X2 state3FF_state_U5 ( .A(enData), .Z(state3FF_state_n6) );
  BUF_X1 state3FF_state_U4 ( .A(selP), .Z(state3FF_state_n11) );
  BUF_X1 state3FF_state_U3 ( .A(selP), .Z(state3FF_state_n12) );
  BUF_X1 state3FF_state_U2 ( .A(selP), .Z(state3FF_state_n9) );
  BUF_X1 state3FF_state_U1 ( .A(selP), .Z(state3FF_state_n10) );
  OAI21_X1 state3FF_state_gff_1_SFF_0_U5 ( .B1(enData), .B2(
        state3FF_state_gff_1_SFF_0_n8), .A(state3FF_state_gff_1_SFF_0_n12), 
        .ZN(state3FF_state_gff_1_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_1_SFF_0_U4 ( .B1(state3FF_state_gff_1_SFF_0_n10), .B2(state3FF_n3), .C1(state3FF_state_gff_1_SFF_0_n11), .C2(
        state3FF_inputPar[0]), .A(enData), .ZN(state3FF_state_gff_1_SFF_0_n12)
         );
  INV_X1 state3FF_state_gff_1_SFF_0_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_1_SFF_0_n11) );
  INV_X1 state3FF_state_gff_1_SFF_0_U2 ( .A(state3FF_state_gff_1_SFF_0_n11), 
        .ZN(state3FF_state_gff_1_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_1_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_1_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[0]), 
        .QN(state3FF_state_gff_1_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_1_SFF_1_U5 ( .B1(enData), .B2(
        state3FF_state_gff_1_SFF_1_n8), .A(state3FF_state_gff_1_SFF_1_n12), 
        .ZN(state3FF_state_gff_1_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_1_SFF_1_U4 ( .B1(state3FF_state_gff_1_SFF_1_n10), .B2(state3FF_n2), .C1(state3FF_state_gff_1_SFF_1_n11), .C2(
        state3FF_inputPar[1]), .A(enData), .ZN(state3FF_state_gff_1_SFF_1_n12)
         );
  INV_X1 state3FF_state_gff_1_SFF_1_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_1_SFF_1_n11) );
  INV_X1 state3FF_state_gff_1_SFF_1_U2 ( .A(state3FF_state_gff_1_SFF_1_n11), 
        .ZN(state3FF_state_gff_1_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_1_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_1_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[16]), 
        .QN(state3FF_state_gff_1_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_1_SFF_2_U5 ( .B1(enData), .B2(
        state3FF_state_gff_1_SFF_2_n8), .A(state3FF_state_gff_1_SFF_2_n12), 
        .ZN(state3FF_state_gff_1_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_1_SFF_2_U4 ( .B1(state3FF_state_gff_1_SFF_2_n10), .B2(state3FF_n1), .C1(state3FF_state_gff_1_SFF_2_n11), .C2(
        state3FF_inputPar[2]), .A(enData), .ZN(state3FF_state_gff_1_SFF_2_n12)
         );
  INV_X1 state3FF_state_gff_1_SFF_2_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_1_SFF_2_n11) );
  INV_X1 state3FF_state_gff_1_SFF_2_U2 ( .A(state3FF_state_gff_1_SFF_2_n11), 
        .ZN(state3FF_state_gff_1_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_1_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_1_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[32]), 
        .QN(state3FF_state_gff_1_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_1_SFF_3_U5 ( .B1(enData), .B2(
        state3FF_state_gff_1_SFF_3_n8), .A(state3FF_state_gff_1_SFF_3_n12), 
        .ZN(state3FF_state_gff_1_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_1_SFF_3_U4 ( .B1(state3FF_state_gff_1_SFF_3_n10), .B2(state3FF_n4), .C1(state3FF_state_gff_1_SFF_3_n11), .C2(
        state3FF_inputPar[3]), .A(enData), .ZN(state3FF_state_gff_1_SFF_3_n12)
         );
  INV_X1 state3FF_state_gff_1_SFF_3_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_1_SFF_3_n11) );
  INV_X1 state3FF_state_gff_1_SFF_3_U2 ( .A(state3FF_state_gff_1_SFF_3_n11), 
        .ZN(state3FF_state_gff_1_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_1_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_1_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[48]), 
        .QN(state3FF_state_gff_1_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_2_SFF_0_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_2_SFF_0_n8), .A(state3FF_state_gff_2_SFF_0_n12), 
        .ZN(state3FF_state_gff_2_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_2_SFF_0_U4 ( .B1(state3FF_state_gff_2_SFF_0_n10), .B2(state3FF_inputPar[0]), .C1(state3FF_state_gff_2_SFF_0_n11), .C2(
        state3FF_inputPar[4]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_2_SFF_0_n12) );
  INV_X1 state3FF_state_gff_2_SFF_0_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_2_SFF_0_n11) );
  INV_X1 state3FF_state_gff_2_SFF_0_U2 ( .A(state3FF_state_gff_2_SFF_0_n11), 
        .ZN(state3FF_state_gff_2_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_2_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_2_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[1]), 
        .QN(state3FF_state_gff_2_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_2_SFF_1_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_2_SFF_1_n8), .A(state3FF_state_gff_2_SFF_1_n12), 
        .ZN(state3FF_state_gff_2_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_2_SFF_1_U4 ( .B1(state3FF_state_gff_2_SFF_1_n10), .B2(state3FF_inputPar[16]), .C1(state3FF_state_gff_2_SFF_1_n11), .C2(
        state3FF_inputPar[5]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_2_SFF_1_n12) );
  INV_X1 state3FF_state_gff_2_SFF_1_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_2_SFF_1_n11) );
  INV_X1 state3FF_state_gff_2_SFF_1_U2 ( .A(state3FF_state_gff_2_SFF_1_n11), 
        .ZN(state3FF_state_gff_2_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_2_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_2_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[17]), 
        .QN(state3FF_state_gff_2_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_2_SFF_2_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_2_SFF_2_n8), .A(state3FF_state_gff_2_SFF_2_n12), 
        .ZN(state3FF_state_gff_2_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_2_SFF_2_U4 ( .B1(state3FF_state_gff_2_SFF_2_n10), .B2(state3FF_inputPar[32]), .C1(state3FF_state_gff_2_SFF_2_n11), .C2(
        state3FF_inputPar[6]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_2_SFF_2_n12) );
  INV_X1 state3FF_state_gff_2_SFF_2_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_2_SFF_2_n11) );
  INV_X1 state3FF_state_gff_2_SFF_2_U2 ( .A(state3FF_state_gff_2_SFF_2_n11), 
        .ZN(state3FF_state_gff_2_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_2_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_2_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[33]), 
        .QN(state3FF_state_gff_2_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_2_SFF_3_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_2_SFF_3_n8), .A(state3FF_state_gff_2_SFF_3_n12), 
        .ZN(state3FF_state_gff_2_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_2_SFF_3_U4 ( .B1(state3FF_state_gff_2_SFF_3_n10), .B2(state3FF_inputPar[48]), .C1(state3FF_state_gff_2_SFF_3_n11), .C2(
        state3FF_inputPar[7]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_2_SFF_3_n12) );
  INV_X1 state3FF_state_gff_2_SFF_3_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_2_SFF_3_n11) );
  INV_X1 state3FF_state_gff_2_SFF_3_U2 ( .A(state3FF_state_gff_2_SFF_3_n11), 
        .ZN(state3FF_state_gff_2_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_2_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_2_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[49]), 
        .QN(state3FF_state_gff_2_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_3_SFF_0_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_3_SFF_0_n8), .A(state3FF_state_gff_3_SFF_0_n12), 
        .ZN(state3FF_state_gff_3_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_3_SFF_0_U4 ( .B1(state3FF_state_gff_3_SFF_0_n10), .B2(state3FF_inputPar[1]), .C1(state3FF_state_gff_3_SFF_0_n11), .C2(
        state3FF_inputPar[8]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_3_SFF_0_n12) );
  INV_X1 state3FF_state_gff_3_SFF_0_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_3_SFF_0_n11) );
  INV_X1 state3FF_state_gff_3_SFF_0_U2 ( .A(state3FF_state_gff_3_SFF_0_n11), 
        .ZN(state3FF_state_gff_3_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_3_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_3_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[2]), 
        .QN(state3FF_state_gff_3_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_3_SFF_1_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_3_SFF_1_n8), .A(state3FF_state_gff_3_SFF_1_n12), 
        .ZN(state3FF_state_gff_3_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_3_SFF_1_U4 ( .B1(state3FF_state_gff_3_SFF_1_n10), .B2(state3FF_inputPar[17]), .C1(state3FF_state_gff_3_SFF_1_n11), .C2(
        state3FF_inputPar[9]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_3_SFF_1_n12) );
  INV_X1 state3FF_state_gff_3_SFF_1_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_3_SFF_1_n11) );
  INV_X1 state3FF_state_gff_3_SFF_1_U2 ( .A(state3FF_state_gff_3_SFF_1_n11), 
        .ZN(state3FF_state_gff_3_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_3_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_3_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[18]), 
        .QN(state3FF_state_gff_3_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_3_SFF_2_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_3_SFF_2_n7), .A(state3FF_state_gff_3_SFF_2_n11), 
        .ZN(state3FF_state_gff_3_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_3_SFF_2_U4 ( .B1(state3FF_state_gff_3_SFF_2_n9), 
        .B2(state3FF_inputPar[33]), .C1(state3FF_state_gff_3_SFF_2_n10), .C2(
        state3FF_inputPar[10]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_3_SFF_2_n11) );
  INV_X1 state3FF_state_gff_3_SFF_2_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_3_SFF_2_n10) );
  INV_X1 state3FF_state_gff_3_SFF_2_U2 ( .A(state3FF_state_gff_3_SFF_2_n10), 
        .ZN(state3FF_state_gff_3_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_3_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_3_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[34]), 
        .QN(state3FF_state_gff_3_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_3_SFF_3_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_3_SFF_3_n7), .A(state3FF_state_gff_3_SFF_3_n11), 
        .ZN(state3FF_state_gff_3_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_3_SFF_3_U4 ( .B1(state3FF_state_gff_3_SFF_3_n9), 
        .B2(state3FF_inputPar[49]), .C1(state3FF_state_gff_3_SFF_3_n10), .C2(
        state3FF_inputPar[11]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_3_SFF_3_n11) );
  INV_X1 state3FF_state_gff_3_SFF_3_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_3_SFF_3_n10) );
  INV_X1 state3FF_state_gff_3_SFF_3_U2 ( .A(state3FF_state_gff_3_SFF_3_n10), 
        .ZN(state3FF_state_gff_3_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_3_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_3_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[50]), 
        .QN(state3FF_state_gff_3_SFF_3_n7) );
  OAI21_X1 state3FF_state_gff_4_SFF_0_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_4_SFF_0_n7), .A(state3FF_state_gff_4_SFF_0_n11), 
        .ZN(state3FF_state_gff_4_SFF_0_n6) );
  OAI221_X1 state3FF_state_gff_4_SFF_0_U4 ( .B1(state3FF_state_gff_4_SFF_0_n9), 
        .B2(state3FF_inputPar[2]), .C1(state3FF_state_gff_4_SFF_0_n10), .C2(
        state3FF_inputPar[12]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_4_SFF_0_n11) );
  INV_X1 state3FF_state_gff_4_SFF_0_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_4_SFF_0_n10) );
  INV_X1 state3FF_state_gff_4_SFF_0_U2 ( .A(state3FF_state_gff_4_SFF_0_n10), 
        .ZN(state3FF_state_gff_4_SFF_0_n9) );
  DFF_X1 state3FF_state_gff_4_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_4_SFF_0_n6), .CK(clk), .Q(state3FF_inputPar[3]), 
        .QN(state3FF_state_gff_4_SFF_0_n7) );
  OAI21_X1 state3FF_state_gff_4_SFF_1_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_4_SFF_1_n7), .A(state3FF_state_gff_4_SFF_1_n11), 
        .ZN(state3FF_state_gff_4_SFF_1_n6) );
  OAI221_X1 state3FF_state_gff_4_SFF_1_U4 ( .B1(state3FF_state_gff_4_SFF_1_n9), 
        .B2(state3FF_inputPar[18]), .C1(state3FF_state_gff_4_SFF_1_n10), .C2(
        state3FF_inputPar[13]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_4_SFF_1_n11) );
  INV_X1 state3FF_state_gff_4_SFF_1_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_4_SFF_1_n10) );
  INV_X1 state3FF_state_gff_4_SFF_1_U2 ( .A(state3FF_state_gff_4_SFF_1_n10), 
        .ZN(state3FF_state_gff_4_SFF_1_n9) );
  DFF_X1 state3FF_state_gff_4_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_4_SFF_1_n6), .CK(clk), .Q(state3FF_inputPar[19]), 
        .QN(state3FF_state_gff_4_SFF_1_n7) );
  OAI21_X1 state3FF_state_gff_4_SFF_2_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_4_SFF_2_n7), .A(state3FF_state_gff_4_SFF_2_n11), 
        .ZN(state3FF_state_gff_4_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_4_SFF_2_U4 ( .B1(state3FF_state_gff_4_SFF_2_n9), 
        .B2(state3FF_inputPar[34]), .C1(state3FF_state_gff_4_SFF_2_n10), .C2(
        state3FF_inputPar[14]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_4_SFF_2_n11) );
  INV_X1 state3FF_state_gff_4_SFF_2_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_4_SFF_2_n10) );
  INV_X1 state3FF_state_gff_4_SFF_2_U2 ( .A(state3FF_state_gff_4_SFF_2_n10), 
        .ZN(state3FF_state_gff_4_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_4_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_4_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[35]), 
        .QN(state3FF_state_gff_4_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_4_SFF_3_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_4_SFF_3_n7), .A(state3FF_state_gff_4_SFF_3_n11), 
        .ZN(state3FF_state_gff_4_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_4_SFF_3_U4 ( .B1(state3FF_state_gff_4_SFF_3_n9), 
        .B2(state3FF_inputPar[50]), .C1(state3FF_state_gff_4_SFF_3_n10), .C2(
        state3FF_inputPar[15]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_4_SFF_3_n11) );
  INV_X1 state3FF_state_gff_4_SFF_3_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_4_SFF_3_n10) );
  INV_X1 state3FF_state_gff_4_SFF_3_U2 ( .A(state3FF_state_gff_4_SFF_3_n10), 
        .ZN(state3FF_state_gff_4_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_4_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_4_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[51]), 
        .QN(state3FF_state_gff_4_SFF_3_n7) );
  OAI21_X1 state3FF_state_gff_5_SFF_0_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_5_SFF_0_n8), .A(state3FF_state_gff_5_SFF_0_n12), 
        .ZN(state3FF_state_gff_5_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_5_SFF_0_U4 ( .B1(state3FF_state_gff_5_SFF_0_n10), .B2(state3FF_inputPar[3]), .C1(state3FF_state_gff_5_SFF_0_n11), .C2(
        state3FF_inputPar[16]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_5_SFF_0_n12) );
  INV_X1 state3FF_state_gff_5_SFF_0_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_5_SFF_0_n11) );
  INV_X1 state3FF_state_gff_5_SFF_0_U2 ( .A(state3FF_state_gff_5_SFF_0_n11), 
        .ZN(state3FF_state_gff_5_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_5_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_5_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[4]), 
        .QN(state3FF_state_gff_5_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_5_SFF_1_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_5_SFF_1_n8), .A(state3FF_state_gff_5_SFF_1_n12), 
        .ZN(state3FF_state_gff_5_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_5_SFF_1_U4 ( .B1(state3FF_state_gff_5_SFF_1_n10), .B2(state3FF_inputPar[19]), .C1(state3FF_state_gff_5_SFF_1_n11), .C2(
        state3FF_inputPar[17]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_5_SFF_1_n12) );
  INV_X1 state3FF_state_gff_5_SFF_1_U3 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_5_SFF_1_n11) );
  INV_X1 state3FF_state_gff_5_SFF_1_U2 ( .A(state3FF_state_gff_5_SFF_1_n11), 
        .ZN(state3FF_state_gff_5_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_5_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_5_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[20]), 
        .QN(state3FF_state_gff_5_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_5_SFF_2_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_5_SFF_2_n8), .A(state3FF_state_gff_5_SFF_2_n11), 
        .ZN(state3FF_state_gff_5_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_5_SFF_2_U3 ( .B1(state3FF_state_n9), .B2(
        state3FF_inputPar[35]), .C1(state3FF_state_gff_5_SFF_2_n10), .C2(
        state3FF_inputPar[18]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_5_SFF_2_n11) );
  INV_X1 state3FF_state_gff_5_SFF_2_U2 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_5_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_5_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_5_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[36]), 
        .QN(state3FF_state_gff_5_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_5_SFF_3_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_5_SFF_3_n8), .A(state3FF_state_gff_5_SFF_3_n11), 
        .ZN(state3FF_state_gff_5_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_5_SFF_3_U3 ( .B1(state3FF_state_n9), .B2(
        state3FF_inputPar[51]), .C1(state3FF_state_gff_5_SFF_3_n10), .C2(
        state3FF_inputPar[19]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_5_SFF_3_n11) );
  INV_X1 state3FF_state_gff_5_SFF_3_U2 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_5_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_5_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_5_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[52]), 
        .QN(state3FF_state_gff_5_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_6_SFF_0_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_6_SFF_0_n8), .A(state3FF_state_gff_6_SFF_0_n11), 
        .ZN(state3FF_state_gff_6_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_6_SFF_0_U3 ( .B1(state3FF_state_n9), .B2(
        state3FF_inputPar[4]), .C1(state3FF_state_gff_6_SFF_0_n10), .C2(
        state3FF_inputPar[20]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_6_SFF_0_n11) );
  INV_X1 state3FF_state_gff_6_SFF_0_U2 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_6_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_6_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_6_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[5]), 
        .QN(state3FF_state_gff_6_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_6_SFF_1_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_6_SFF_1_n8), .A(state3FF_state_gff_6_SFF_1_n11), 
        .ZN(state3FF_state_gff_6_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_6_SFF_1_U3 ( .B1(state3FF_state_n9), .B2(
        state3FF_inputPar[20]), .C1(state3FF_state_gff_6_SFF_1_n10), .C2(
        state3FF_inputPar[21]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_6_SFF_1_n11) );
  INV_X1 state3FF_state_gff_6_SFF_1_U2 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_6_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_6_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_6_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[21]), 
        .QN(state3FF_state_gff_6_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_6_SFF_2_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_6_SFF_2_n8), .A(state3FF_state_gff_6_SFF_2_n11), 
        .ZN(state3FF_state_gff_6_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_6_SFF_2_U3 ( .B1(state3FF_state_n9), .B2(
        state3FF_inputPar[36]), .C1(state3FF_state_gff_6_SFF_2_n10), .C2(
        state3FF_inputPar[22]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_6_SFF_2_n11) );
  INV_X1 state3FF_state_gff_6_SFF_2_U2 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_6_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_6_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_6_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[37]), 
        .QN(state3FF_state_gff_6_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_6_SFF_3_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_6_SFF_3_n8), .A(state3FF_state_gff_6_SFF_3_n11), 
        .ZN(state3FF_state_gff_6_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_6_SFF_3_U3 ( .B1(state3FF_state_n9), .B2(
        state3FF_inputPar[52]), .C1(state3FF_state_gff_6_SFF_3_n10), .C2(
        state3FF_inputPar[23]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_6_SFF_3_n11) );
  INV_X1 state3FF_state_gff_6_SFF_3_U2 ( .A(state3FF_state_n9), .ZN(
        state3FF_state_gff_6_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_6_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_6_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[53]), 
        .QN(state3FF_state_gff_6_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_7_SFF_0_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_7_SFF_0_n8), .A(state3FF_state_gff_7_SFF_0_n11), 
        .ZN(state3FF_state_gff_7_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_7_SFF_0_U3 ( .B1(state3FF_state_n11), .B2(
        state3FF_inputPar[5]), .C1(state3FF_state_gff_7_SFF_0_n10), .C2(
        state3FF_inputPar[24]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_7_SFF_0_n11) );
  INV_X1 state3FF_state_gff_7_SFF_0_U2 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_7_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_7_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_7_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[6]), 
        .QN(state3FF_state_gff_7_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_7_SFF_1_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_7_SFF_1_n8), .A(state3FF_state_gff_7_SFF_1_n11), 
        .ZN(state3FF_state_gff_7_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_7_SFF_1_U3 ( .B1(state3FF_state_n11), .B2(
        state3FF_inputPar[21]), .C1(state3FF_state_gff_7_SFF_1_n10), .C2(
        state3FF_inputPar[25]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_7_SFF_1_n11) );
  INV_X1 state3FF_state_gff_7_SFF_1_U2 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_7_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_7_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_7_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[22]), 
        .QN(state3FF_state_gff_7_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_7_SFF_2_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_7_SFF_2_n7), .A(state3FF_state_gff_7_SFF_2_n11), 
        .ZN(state3FF_state_gff_7_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_7_SFF_2_U4 ( .B1(state3FF_state_gff_7_SFF_2_n9), 
        .B2(state3FF_inputPar[37]), .C1(state3FF_state_gff_7_SFF_2_n10), .C2(
        state3FF_inputPar[26]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_7_SFF_2_n11) );
  INV_X1 state3FF_state_gff_7_SFF_2_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_7_SFF_2_n10) );
  INV_X1 state3FF_state_gff_7_SFF_2_U2 ( .A(state3FF_state_gff_7_SFF_2_n10), 
        .ZN(state3FF_state_gff_7_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_7_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_7_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[38]), 
        .QN(state3FF_state_gff_7_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_7_SFF_3_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_7_SFF_3_n7), .A(state3FF_state_gff_7_SFF_3_n11), 
        .ZN(state3FF_state_gff_7_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_7_SFF_3_U4 ( .B1(state3FF_state_gff_7_SFF_3_n9), 
        .B2(state3FF_inputPar[53]), .C1(state3FF_state_gff_7_SFF_3_n10), .C2(
        state3FF_inputPar[27]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_7_SFF_3_n11) );
  INV_X1 state3FF_state_gff_7_SFF_3_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_7_SFF_3_n10) );
  INV_X1 state3FF_state_gff_7_SFF_3_U2 ( .A(state3FF_state_gff_7_SFF_3_n10), 
        .ZN(state3FF_state_gff_7_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_7_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_7_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[54]), 
        .QN(state3FF_state_gff_7_SFF_3_n7) );
  OAI21_X1 state3FF_state_gff_8_SFF_0_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_8_SFF_0_n7), .A(state3FF_state_gff_8_SFF_0_n11), 
        .ZN(state3FF_state_gff_8_SFF_0_n6) );
  OAI221_X1 state3FF_state_gff_8_SFF_0_U4 ( .B1(state3FF_state_gff_8_SFF_0_n9), 
        .B2(state3FF_inputPar[6]), .C1(state3FF_state_gff_8_SFF_0_n10), .C2(
        state3FF_inputPar[28]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_8_SFF_0_n11) );
  INV_X1 state3FF_state_gff_8_SFF_0_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_8_SFF_0_n10) );
  INV_X1 state3FF_state_gff_8_SFF_0_U2 ( .A(state3FF_state_gff_8_SFF_0_n10), 
        .ZN(state3FF_state_gff_8_SFF_0_n9) );
  DFF_X1 state3FF_state_gff_8_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_8_SFF_0_n6), .CK(clk), .Q(state3FF_inputPar[7]), 
        .QN(state3FF_state_gff_8_SFF_0_n7) );
  OAI21_X1 state3FF_state_gff_8_SFF_1_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_8_SFF_1_n7), .A(state3FF_state_gff_8_SFF_1_n11), 
        .ZN(state3FF_state_gff_8_SFF_1_n6) );
  OAI221_X1 state3FF_state_gff_8_SFF_1_U4 ( .B1(state3FF_state_gff_8_SFF_1_n9), 
        .B2(state3FF_inputPar[22]), .C1(state3FF_state_gff_8_SFF_1_n10), .C2(
        state3FF_inputPar[29]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_8_SFF_1_n11) );
  INV_X1 state3FF_state_gff_8_SFF_1_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_8_SFF_1_n10) );
  INV_X1 state3FF_state_gff_8_SFF_1_U2 ( .A(state3FF_state_gff_8_SFF_1_n10), 
        .ZN(state3FF_state_gff_8_SFF_1_n9) );
  DFF_X1 state3FF_state_gff_8_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_8_SFF_1_n6), .CK(clk), .Q(state3FF_inputPar[23]), 
        .QN(state3FF_state_gff_8_SFF_1_n7) );
  OAI21_X1 state3FF_state_gff_8_SFF_2_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_8_SFF_2_n7), .A(state3FF_state_gff_8_SFF_2_n11), 
        .ZN(state3FF_state_gff_8_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_8_SFF_2_U4 ( .B1(state3FF_state_gff_8_SFF_2_n9), 
        .B2(state3FF_inputPar[38]), .C1(state3FF_state_gff_8_SFF_2_n10), .C2(
        state3FF_inputPar[30]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_8_SFF_2_n11) );
  INV_X1 state3FF_state_gff_8_SFF_2_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_8_SFF_2_n10) );
  INV_X1 state3FF_state_gff_8_SFF_2_U2 ( .A(state3FF_state_gff_8_SFF_2_n10), 
        .ZN(state3FF_state_gff_8_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_8_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_8_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[39]), 
        .QN(state3FF_state_gff_8_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_8_SFF_3_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_8_SFF_3_n7), .A(state3FF_state_gff_8_SFF_3_n11), 
        .ZN(state3FF_state_gff_8_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_8_SFF_3_U4 ( .B1(state3FF_state_gff_8_SFF_3_n9), 
        .B2(state3FF_inputPar[54]), .C1(state3FF_state_gff_8_SFF_3_n10), .C2(
        state3FF_inputPar[31]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_8_SFF_3_n11) );
  INV_X1 state3FF_state_gff_8_SFF_3_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_8_SFF_3_n10) );
  INV_X1 state3FF_state_gff_8_SFF_3_U2 ( .A(state3FF_state_gff_8_SFF_3_n10), 
        .ZN(state3FF_state_gff_8_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_8_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_8_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[55]), 
        .QN(state3FF_state_gff_8_SFF_3_n7) );
  OAI21_X1 state3FF_state_gff_9_SFF_0_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_9_SFF_0_n8), .A(state3FF_state_gff_9_SFF_0_n12), 
        .ZN(state3FF_state_gff_9_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_9_SFF_0_U4 ( .B1(state3FF_state_gff_9_SFF_0_n10), .B2(state3FF_inputPar[7]), .C1(state3FF_state_gff_9_SFF_0_n11), .C2(
        state3FF_inputPar[32]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_9_SFF_0_n12) );
  INV_X1 state3FF_state_gff_9_SFF_0_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_9_SFF_0_n11) );
  INV_X1 state3FF_state_gff_9_SFF_0_U2 ( .A(state3FF_state_gff_9_SFF_0_n11), 
        .ZN(state3FF_state_gff_9_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_9_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_9_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[8]), 
        .QN(state3FF_state_gff_9_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_9_SFF_1_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_9_SFF_1_n8), .A(state3FF_state_gff_9_SFF_1_n12), 
        .ZN(state3FF_state_gff_9_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_9_SFF_1_U4 ( .B1(state3FF_state_gff_9_SFF_1_n10), .B2(state3FF_inputPar[23]), .C1(state3FF_state_gff_9_SFF_1_n11), .C2(
        state3FF_inputPar[33]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_9_SFF_1_n12) );
  INV_X1 state3FF_state_gff_9_SFF_1_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_9_SFF_1_n11) );
  INV_X1 state3FF_state_gff_9_SFF_1_U2 ( .A(state3FF_state_gff_9_SFF_1_n11), 
        .ZN(state3FF_state_gff_9_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_9_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_9_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[24]), 
        .QN(state3FF_state_gff_9_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_9_SFF_2_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_9_SFF_2_n8), .A(state3FF_state_gff_9_SFF_2_n12), 
        .ZN(state3FF_state_gff_9_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_9_SFF_2_U4 ( .B1(state3FF_state_gff_9_SFF_2_n10), .B2(state3FF_inputPar[39]), .C1(state3FF_state_gff_9_SFF_2_n11), .C2(
        state3FF_inputPar[34]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_9_SFF_2_n12) );
  INV_X1 state3FF_state_gff_9_SFF_2_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_9_SFF_2_n11) );
  INV_X1 state3FF_state_gff_9_SFF_2_U2 ( .A(state3FF_state_gff_9_SFF_2_n11), 
        .ZN(state3FF_state_gff_9_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_9_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_9_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[40]), 
        .QN(state3FF_state_gff_9_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_9_SFF_3_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_9_SFF_3_n8), .A(state3FF_state_gff_9_SFF_3_n12), 
        .ZN(state3FF_state_gff_9_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_9_SFF_3_U4 ( .B1(state3FF_state_gff_9_SFF_3_n10), .B2(state3FF_inputPar[55]), .C1(state3FF_state_gff_9_SFF_3_n11), .C2(
        state3FF_inputPar[35]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_9_SFF_3_n12) );
  INV_X1 state3FF_state_gff_9_SFF_3_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_9_SFF_3_n11) );
  INV_X1 state3FF_state_gff_9_SFF_3_U2 ( .A(state3FF_state_gff_9_SFF_3_n11), 
        .ZN(state3FF_state_gff_9_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_9_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_9_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[56]), 
        .QN(state3FF_state_gff_9_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_10_SFF_0_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_10_SFF_0_n8), .A(state3FF_state_gff_10_SFF_0_n12), 
        .ZN(state3FF_state_gff_10_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_10_SFF_0_U4 ( .B1(
        state3FF_state_gff_10_SFF_0_n10), .B2(state3FF_inputPar[8]), .C1(
        state3FF_state_gff_10_SFF_0_n11), .C2(state3FF_inputPar[36]), .A(
        state3FF_state_n6), .ZN(state3FF_state_gff_10_SFF_0_n12) );
  INV_X1 state3FF_state_gff_10_SFF_0_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_10_SFF_0_n11) );
  INV_X1 state3FF_state_gff_10_SFF_0_U2 ( .A(state3FF_state_gff_10_SFF_0_n11), 
        .ZN(state3FF_state_gff_10_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_10_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_10_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[9]), 
        .QN(state3FF_state_gff_10_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_10_SFF_1_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_10_SFF_1_n8), .A(state3FF_state_gff_10_SFF_1_n12), 
        .ZN(state3FF_state_gff_10_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_10_SFF_1_U4 ( .B1(
        state3FF_state_gff_10_SFF_1_n10), .B2(state3FF_inputPar[24]), .C1(
        state3FF_state_gff_10_SFF_1_n11), .C2(state3FF_inputPar[37]), .A(
        state3FF_state_n6), .ZN(state3FF_state_gff_10_SFF_1_n12) );
  INV_X1 state3FF_state_gff_10_SFF_1_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_10_SFF_1_n11) );
  INV_X1 state3FF_state_gff_10_SFF_1_U2 ( .A(state3FF_state_gff_10_SFF_1_n11), 
        .ZN(state3FF_state_gff_10_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_10_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_10_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[25]), 
        .QN(state3FF_state_gff_10_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_10_SFF_2_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_10_SFF_2_n8), .A(state3FF_state_gff_10_SFF_2_n12), 
        .ZN(state3FF_state_gff_10_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_10_SFF_2_U4 ( .B1(
        state3FF_state_gff_10_SFF_2_n10), .B2(state3FF_inputPar[40]), .C1(
        state3FF_state_gff_10_SFF_2_n11), .C2(state3FF_inputPar[38]), .A(
        state3FF_state_n6), .ZN(state3FF_state_gff_10_SFF_2_n12) );
  INV_X1 state3FF_state_gff_10_SFF_2_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_10_SFF_2_n11) );
  INV_X1 state3FF_state_gff_10_SFF_2_U2 ( .A(state3FF_state_gff_10_SFF_2_n11), 
        .ZN(state3FF_state_gff_10_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_10_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_10_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[41]), 
        .QN(state3FF_state_gff_10_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_10_SFF_3_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_10_SFF_3_n8), .A(state3FF_state_gff_10_SFF_3_n12), 
        .ZN(state3FF_state_gff_10_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_10_SFF_3_U4 ( .B1(
        state3FF_state_gff_10_SFF_3_n10), .B2(state3FF_inputPar[56]), .C1(
        state3FF_state_gff_10_SFF_3_n11), .C2(state3FF_inputPar[39]), .A(
        state3FF_state_n6), .ZN(state3FF_state_gff_10_SFF_3_n12) );
  INV_X1 state3FF_state_gff_10_SFF_3_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_10_SFF_3_n11) );
  INV_X1 state3FF_state_gff_10_SFF_3_U2 ( .A(state3FF_state_gff_10_SFF_3_n11), 
        .ZN(state3FF_state_gff_10_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_10_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_10_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[57]), 
        .QN(state3FF_state_gff_10_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_11_SFF_0_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_11_SFF_0_n8), .A(state3FF_state_gff_11_SFF_0_n11), 
        .ZN(state3FF_state_gff_11_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_11_SFF_0_U3 ( .B1(state3FF_state_n11), .B2(
        state3FF_inputPar[9]), .C1(state3FF_state_gff_11_SFF_0_n10), .C2(
        state3FF_inputPar[40]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_11_SFF_0_n11) );
  INV_X1 state3FF_state_gff_11_SFF_0_U2 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_11_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_11_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_11_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[10]), 
        .QN(state3FF_state_gff_11_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_11_SFF_1_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_11_SFF_1_n8), .A(state3FF_state_gff_11_SFF_1_n11), 
        .ZN(state3FF_state_gff_11_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_11_SFF_1_U3 ( .B1(state3FF_state_n11), .B2(
        state3FF_inputPar[25]), .C1(state3FF_state_gff_11_SFF_1_n10), .C2(
        state3FF_inputPar[41]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_11_SFF_1_n11) );
  INV_X1 state3FF_state_gff_11_SFF_1_U2 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_11_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_11_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_11_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[26]), 
        .QN(state3FF_state_gff_11_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_11_SFF_2_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_11_SFF_2_n7), .A(state3FF_state_gff_11_SFF_2_n11), 
        .ZN(state3FF_state_gff_11_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_11_SFF_2_U4 ( .B1(
        state3FF_state_gff_11_SFF_2_n9), .B2(state3FF_inputPar[41]), .C1(
        state3FF_state_gff_11_SFF_2_n10), .C2(state3FF_inputPar[42]), .A(
        state3FF_state_n7), .ZN(state3FF_state_gff_11_SFF_2_n11) );
  INV_X1 state3FF_state_gff_11_SFF_2_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_11_SFF_2_n10) );
  INV_X1 state3FF_state_gff_11_SFF_2_U2 ( .A(state3FF_state_gff_11_SFF_2_n10), 
        .ZN(state3FF_state_gff_11_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_11_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_11_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[42]), 
        .QN(state3FF_state_gff_11_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_11_SFF_3_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_11_SFF_3_n7), .A(state3FF_state_gff_11_SFF_3_n11), 
        .ZN(state3FF_state_gff_11_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_11_SFF_3_U4 ( .B1(
        state3FF_state_gff_11_SFF_3_n9), .B2(state3FF_inputPar[57]), .C1(
        state3FF_state_gff_11_SFF_3_n10), .C2(state3FF_inputPar[43]), .A(
        state3FF_state_n7), .ZN(state3FF_state_gff_11_SFF_3_n11) );
  INV_X1 state3FF_state_gff_11_SFF_3_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_11_SFF_3_n10) );
  INV_X1 state3FF_state_gff_11_SFF_3_U2 ( .A(state3FF_state_gff_11_SFF_3_n10), 
        .ZN(state3FF_state_gff_11_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_11_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_11_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[58]), 
        .QN(state3FF_state_gff_11_SFF_3_n7) );
  OAI21_X1 state3FF_state_gff_12_SFF_0_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_12_SFF_0_n7), .A(state3FF_state_gff_12_SFF_0_n11), 
        .ZN(state3FF_state_gff_12_SFF_0_n6) );
  OAI221_X1 state3FF_state_gff_12_SFF_0_U4 ( .B1(
        state3FF_state_gff_12_SFF_0_n9), .B2(state3FF_inputPar[10]), .C1(
        state3FF_state_gff_12_SFF_0_n10), .C2(state3FF_inputPar[44]), .A(
        state3FF_state_n8), .ZN(state3FF_state_gff_12_SFF_0_n11) );
  INV_X1 state3FF_state_gff_12_SFF_0_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_12_SFF_0_n10) );
  INV_X1 state3FF_state_gff_12_SFF_0_U2 ( .A(state3FF_state_gff_12_SFF_0_n10), 
        .ZN(state3FF_state_gff_12_SFF_0_n9) );
  DFF_X1 state3FF_state_gff_12_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_12_SFF_0_n6), .CK(clk), .Q(state3FF_inputPar[11]), 
        .QN(state3FF_state_gff_12_SFF_0_n7) );
  OAI21_X1 state3FF_state_gff_12_SFF_1_U5 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_12_SFF_1_n7), .A(state3FF_state_gff_12_SFF_1_n11), 
        .ZN(state3FF_state_gff_12_SFF_1_n6) );
  OAI221_X1 state3FF_state_gff_12_SFF_1_U4 ( .B1(
        state3FF_state_gff_12_SFF_1_n9), .B2(state3FF_inputPar[26]), .C1(
        state3FF_state_gff_12_SFF_1_n10), .C2(state3FF_inputPar[45]), .A(
        state3FF_state_n8), .ZN(state3FF_state_gff_12_SFF_1_n11) );
  INV_X1 state3FF_state_gff_12_SFF_1_U3 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_12_SFF_1_n10) );
  INV_X1 state3FF_state_gff_12_SFF_1_U2 ( .A(state3FF_state_gff_12_SFF_1_n10), 
        .ZN(state3FF_state_gff_12_SFF_1_n9) );
  DFF_X1 state3FF_state_gff_12_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_12_SFF_1_n6), .CK(clk), .Q(state3FF_inputPar[27]), 
        .QN(state3FF_state_gff_12_SFF_1_n7) );
  OAI21_X1 state3FF_state_gff_12_SFF_2_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_12_SFF_2_n7), .A(state3FF_state_gff_12_SFF_2_n10), 
        .ZN(state3FF_state_gff_12_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_12_SFF_2_U3 ( .B1(state3FF_state_n12), .B2(
        state3FF_inputPar[42]), .C1(state3FF_state_gff_12_SFF_2_n9), .C2(
        state3FF_inputPar[46]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_12_SFF_2_n10) );
  INV_X1 state3FF_state_gff_12_SFF_2_U2 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_12_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_12_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_12_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[43]), 
        .QN(state3FF_state_gff_12_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_12_SFF_3_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_12_SFF_3_n7), .A(state3FF_state_gff_12_SFF_3_n10), 
        .ZN(state3FF_state_gff_12_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_12_SFF_3_U3 ( .B1(state3FF_state_n12), .B2(
        state3FF_inputPar[58]), .C1(state3FF_state_gff_12_SFF_3_n9), .C2(
        state3FF_inputPar[47]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_12_SFF_3_n10) );
  INV_X1 state3FF_state_gff_12_SFF_3_U2 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_12_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_12_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_12_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[59]), 
        .QN(state3FF_state_gff_12_SFF_3_n7) );
  OAI21_X1 state3FF_state_gff_13_SFF_0_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_13_SFF_0_n8), .A(state3FF_state_gff_13_SFF_0_n12), 
        .ZN(state3FF_state_gff_13_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_13_SFF_0_U4 ( .B1(
        state3FF_state_gff_13_SFF_0_n10), .B2(state3FF_inputPar[11]), .C1(
        state3FF_state_gff_13_SFF_0_n11), .C2(state3FF_inputPar[48]), .A(
        state3FF_state_n6), .ZN(state3FF_state_gff_13_SFF_0_n12) );
  INV_X1 state3FF_state_gff_13_SFF_0_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_13_SFF_0_n11) );
  INV_X1 state3FF_state_gff_13_SFF_0_U2 ( .A(state3FF_state_gff_13_SFF_0_n11), 
        .ZN(state3FF_state_gff_13_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_13_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_13_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[12]), 
        .QN(state3FF_state_gff_13_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_13_SFF_1_U5 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_13_SFF_1_n8), .A(state3FF_state_gff_13_SFF_1_n12), 
        .ZN(state3FF_state_gff_13_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_13_SFF_1_U4 ( .B1(
        state3FF_state_gff_13_SFF_1_n10), .B2(state3FF_inputPar[27]), .C1(
        state3FF_state_gff_13_SFF_1_n11), .C2(state3FF_inputPar[49]), .A(
        state3FF_state_n6), .ZN(state3FF_state_gff_13_SFF_1_n12) );
  INV_X1 state3FF_state_gff_13_SFF_1_U3 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_13_SFF_1_n11) );
  INV_X1 state3FF_state_gff_13_SFF_1_U2 ( .A(state3FF_state_gff_13_SFF_1_n11), 
        .ZN(state3FF_state_gff_13_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_13_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_13_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[28]), 
        .QN(state3FF_state_gff_13_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_13_SFF_2_U4 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_13_SFF_2_n8), .A(state3FF_state_gff_13_SFF_2_n11), 
        .ZN(state3FF_state_gff_13_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_13_SFF_2_U3 ( .B1(state3FF_state_n10), .B2(
        state3FF_inputPar[43]), .C1(state3FF_state_gff_13_SFF_2_n10), .C2(
        state3FF_inputPar[50]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_13_SFF_2_n11) );
  INV_X1 state3FF_state_gff_13_SFF_2_U2 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_13_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_13_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_13_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[44]), 
        .QN(state3FF_state_gff_13_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_13_SFF_3_U4 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_13_SFF_3_n8), .A(state3FF_state_gff_13_SFF_3_n11), 
        .ZN(state3FF_state_gff_13_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_13_SFF_3_U3 ( .B1(state3FF_state_n10), .B2(
        state3FF_inputPar[59]), .C1(state3FF_state_gff_13_SFF_3_n10), .C2(
        state3FF_inputPar[51]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_13_SFF_3_n11) );
  INV_X1 state3FF_state_gff_13_SFF_3_U2 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_13_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_13_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_13_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[60]), 
        .QN(state3FF_state_gff_13_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_14_SFF_0_U4 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_14_SFF_0_n8), .A(state3FF_state_gff_14_SFF_0_n11), 
        .ZN(state3FF_state_gff_14_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_14_SFF_0_U3 ( .B1(state3FF_state_n10), .B2(
        state3FF_inputPar[12]), .C1(state3FF_state_gff_14_SFF_0_n10), .C2(
        state3FF_inputPar[52]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_14_SFF_0_n11) );
  INV_X1 state3FF_state_gff_14_SFF_0_U2 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_14_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_14_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_14_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[13]), 
        .QN(state3FF_state_gff_14_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_14_SFF_1_U4 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_14_SFF_1_n8), .A(state3FF_state_gff_14_SFF_1_n11), 
        .ZN(state3FF_state_gff_14_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_14_SFF_1_U3 ( .B1(state3FF_state_n10), .B2(
        state3FF_inputPar[28]), .C1(state3FF_state_gff_14_SFF_1_n10), .C2(
        state3FF_inputPar[53]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_14_SFF_1_n11) );
  INV_X1 state3FF_state_gff_14_SFF_1_U2 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_14_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_14_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_14_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[29]), 
        .QN(state3FF_state_gff_14_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_14_SFF_2_U4 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_14_SFF_2_n8), .A(state3FF_state_gff_14_SFF_2_n11), 
        .ZN(state3FF_state_gff_14_SFF_2_n7) );
  OAI221_X1 state3FF_state_gff_14_SFF_2_U3 ( .B1(state3FF_state_n10), .B2(
        state3FF_inputPar[44]), .C1(state3FF_state_gff_14_SFF_2_n10), .C2(
        state3FF_inputPar[54]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_14_SFF_2_n11) );
  INV_X1 state3FF_state_gff_14_SFF_2_U2 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_14_SFF_2_n10) );
  DFF_X1 state3FF_state_gff_14_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_14_SFF_2_n7), .CK(clk), .Q(state3FF_inputPar[45]), 
        .QN(state3FF_state_gff_14_SFF_2_n8) );
  OAI21_X1 state3FF_state_gff_14_SFF_3_U4 ( .B1(state3FF_state_n6), .B2(
        state3FF_state_gff_14_SFF_3_n8), .A(state3FF_state_gff_14_SFF_3_n11), 
        .ZN(state3FF_state_gff_14_SFF_3_n7) );
  OAI221_X1 state3FF_state_gff_14_SFF_3_U3 ( .B1(state3FF_state_n10), .B2(
        state3FF_inputPar[60]), .C1(state3FF_state_gff_14_SFF_3_n10), .C2(
        state3FF_inputPar[55]), .A(state3FF_state_n6), .ZN(
        state3FF_state_gff_14_SFF_3_n11) );
  INV_X1 state3FF_state_gff_14_SFF_3_U2 ( .A(state3FF_state_n10), .ZN(
        state3FF_state_gff_14_SFF_3_n10) );
  DFF_X1 state3FF_state_gff_14_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_14_SFF_3_n7), .CK(clk), .Q(state3FF_inputPar[61]), 
        .QN(state3FF_state_gff_14_SFF_3_n8) );
  OAI21_X1 state3FF_state_gff_15_SFF_0_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_15_SFF_0_n8), .A(state3FF_state_gff_15_SFF_0_n11), 
        .ZN(state3FF_state_gff_15_SFF_0_n7) );
  OAI221_X1 state3FF_state_gff_15_SFF_0_U3 ( .B1(state3FF_state_n11), .B2(
        state3FF_inputPar[13]), .C1(state3FF_state_gff_15_SFF_0_n10), .C2(
        state3FF_inputPar[56]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_15_SFF_0_n11) );
  INV_X1 state3FF_state_gff_15_SFF_0_U2 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_15_SFF_0_n10) );
  DFF_X1 state3FF_state_gff_15_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_15_SFF_0_n7), .CK(clk), .Q(state3FF_inputPar[14]), 
        .QN(state3FF_state_gff_15_SFF_0_n8) );
  OAI21_X1 state3FF_state_gff_15_SFF_1_U4 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_15_SFF_1_n8), .A(state3FF_state_gff_15_SFF_1_n11), 
        .ZN(state3FF_state_gff_15_SFF_1_n7) );
  OAI221_X1 state3FF_state_gff_15_SFF_1_U3 ( .B1(state3FF_state_n11), .B2(
        state3FF_inputPar[29]), .C1(state3FF_state_gff_15_SFF_1_n10), .C2(
        state3FF_inputPar[57]), .A(state3FF_state_n7), .ZN(
        state3FF_state_gff_15_SFF_1_n11) );
  INV_X1 state3FF_state_gff_15_SFF_1_U2 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_15_SFF_1_n10) );
  DFF_X1 state3FF_state_gff_15_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_15_SFF_1_n7), .CK(clk), .Q(state3FF_inputPar[30]), 
        .QN(state3FF_state_gff_15_SFF_1_n8) );
  OAI21_X1 state3FF_state_gff_15_SFF_2_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_15_SFF_2_n7), .A(state3FF_state_gff_15_SFF_2_n11), 
        .ZN(state3FF_state_gff_15_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_15_SFF_2_U4 ( .B1(
        state3FF_state_gff_15_SFF_2_n9), .B2(state3FF_inputPar[45]), .C1(
        state3FF_state_gff_15_SFF_2_n10), .C2(state3FF_inputPar[58]), .A(
        state3FF_state_n7), .ZN(state3FF_state_gff_15_SFF_2_n11) );
  INV_X1 state3FF_state_gff_15_SFF_2_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_15_SFF_2_n10) );
  INV_X1 state3FF_state_gff_15_SFF_2_U2 ( .A(state3FF_state_gff_15_SFF_2_n10), 
        .ZN(state3FF_state_gff_15_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_15_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_15_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[46]), 
        .QN(state3FF_state_gff_15_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_15_SFF_3_U5 ( .B1(state3FF_state_n7), .B2(
        state3FF_state_gff_15_SFF_3_n7), .A(state3FF_state_gff_15_SFF_3_n11), 
        .ZN(state3FF_state_gff_15_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_15_SFF_3_U4 ( .B1(
        state3FF_state_gff_15_SFF_3_n9), .B2(state3FF_inputPar[61]), .C1(
        state3FF_state_gff_15_SFF_3_n10), .C2(state3FF_inputPar[59]), .A(
        state3FF_state_n7), .ZN(state3FF_state_gff_15_SFF_3_n11) );
  INV_X1 state3FF_state_gff_15_SFF_3_U3 ( .A(state3FF_state_n11), .ZN(
        state3FF_state_gff_15_SFF_3_n10) );
  INV_X1 state3FF_state_gff_15_SFF_3_U2 ( .A(state3FF_state_gff_15_SFF_3_n10), 
        .ZN(state3FF_state_gff_15_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_15_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_15_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[62]), 
        .QN(state3FF_state_gff_15_SFF_3_n7) );
  OAI21_X1 state3FF_state_gff_16_SFF_0_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_16_SFF_0_n7), .A(state3FF_state_gff_16_SFF_0_n10), 
        .ZN(state3FF_state_gff_16_SFF_0_n6) );
  OAI221_X1 state3FF_state_gff_16_SFF_0_U3 ( .B1(state3FF_state_n12), .B2(
        state3FF_inputPar[14]), .C1(state3FF_state_gff_16_SFF_0_n9), .C2(
        state3FF_inputPar[60]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_16_SFF_0_n10) );
  INV_X1 state3FF_state_gff_16_SFF_0_U2 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_16_SFF_0_n9) );
  DFF_X1 state3FF_state_gff_16_SFF_0_Cell_reg ( .D(
        state3FF_state_gff_16_SFF_0_n6), .CK(clk), .Q(state3FF_inputPar[15]), 
        .QN(state3FF_state_gff_16_SFF_0_n7) );
  OAI21_X1 state3FF_state_gff_16_SFF_1_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_16_SFF_1_n7), .A(state3FF_state_gff_16_SFF_1_n10), 
        .ZN(state3FF_state_gff_16_SFF_1_n6) );
  OAI221_X1 state3FF_state_gff_16_SFF_1_U3 ( .B1(state3FF_state_n12), .B2(
        state3FF_inputPar[30]), .C1(state3FF_state_gff_16_SFF_1_n9), .C2(
        state3FF_inputPar[61]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_16_SFF_1_n10) );
  INV_X1 state3FF_state_gff_16_SFF_1_U2 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_16_SFF_1_n9) );
  DFF_X1 state3FF_state_gff_16_SFF_1_Cell_reg ( .D(
        state3FF_state_gff_16_SFF_1_n6), .CK(clk), .Q(state3FF_inputPar[31]), 
        .QN(state3FF_state_gff_16_SFF_1_n7) );
  OAI21_X1 state3FF_state_gff_16_SFF_2_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_16_SFF_2_n7), .A(state3FF_state_gff_16_SFF_2_n10), 
        .ZN(state3FF_state_gff_16_SFF_2_n6) );
  OAI221_X1 state3FF_state_gff_16_SFF_2_U3 ( .B1(state3FF_state_n12), .B2(
        state3FF_inputPar[46]), .C1(state3FF_state_gff_16_SFF_2_n9), .C2(
        state3FF_inputPar[62]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_16_SFF_2_n10) );
  INV_X1 state3FF_state_gff_16_SFF_2_U2 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_16_SFF_2_n9) );
  DFF_X1 state3FF_state_gff_16_SFF_2_Cell_reg ( .D(
        state3FF_state_gff_16_SFF_2_n6), .CK(clk), .Q(state3FF_inputPar[47]), 
        .QN(state3FF_state_gff_16_SFF_2_n7) );
  OAI21_X1 state3FF_state_gff_16_SFF_3_U4 ( .B1(state3FF_state_n8), .B2(
        state3FF_state_gff_16_SFF_3_n7), .A(state3FF_state_gff_16_SFF_3_n10), 
        .ZN(state3FF_state_gff_16_SFF_3_n6) );
  OAI221_X1 state3FF_state_gff_16_SFF_3_U3 ( .B1(state3FF_state_n12), .B2(
        state3FF_inputPar[62]), .C1(state3FF_state_gff_16_SFF_3_n9), .C2(
        state3FF_inputPar[63]), .A(state3FF_state_n8), .ZN(
        state3FF_state_gff_16_SFF_3_n10) );
  INV_X1 state3FF_state_gff_16_SFF_3_U2 ( .A(state3FF_state_n12), .ZN(
        state3FF_state_gff_16_SFF_3_n9) );
  DFF_X1 state3FF_state_gff_16_SFF_3_Cell_reg ( .D(
        state3FF_state_gff_16_SFF_3_n6), .CK(clk), .Q(state3FF_inputPar[63]), 
        .QN(state3FF_state_gff_16_SFF_3_n7) );
  MUX2_X1 key1FF_U10 ( .A(roundkey1[0]), .B(key1[0]), .S(n4), .Z(key1FF_n1) );
  MUX2_X1 key1FF_U9 ( .A(roundkey1[1]), .B(key1[1]), .S(n4), .Z(key1FF_n2) );
  MUX2_X1 key1FF_U8 ( .A(roundkey1[2]), .B(key1[2]), .S(n4), .Z(key1FF_n3) );
  MUX2_X1 key1FF_U7 ( .A(roundkey1[3]), .B(key1[3]), .S(n4), .Z(key1FF_n4) );
  XOR2_X1 key1FF_U6 ( .A(counter[4]), .B(key1FF_outputPar[22]), .Z(
        key1FF_counterAdd[4]) );
  XOR2_X1 key1FF_U5 ( .A(counter[3]), .B(key1FF_outputPar[21]), .Z(
        key1FF_counterAdd[3]) );
  XOR2_X1 key1FF_U4 ( .A(counter[2]), .B(key1FF_outputPar[20]), .Z(
        key1FF_counterAdd[2]) );
  XOR2_X1 key1FF_U3 ( .A(counter[1]), .B(key1FF_outputPar[19]), .Z(
        key1FF_counterAdd[1]) );
  XOR2_X1 key1FF_U2 ( .A(counter[0]), .B(key1FF_outputPar[18]), .Z(
        key1FF_counterAdd[0]) );
  BUF_X2 key1FF_keystate_U9 ( .A(enKey), .Z(key1FF_keystate_n12) );
  BUF_X1 key1FF_keystate_U8 ( .A(selP), .Z(key1FF_keystate_n17) );
  BUF_X2 key1FF_keystate_U7 ( .A(enKey), .Z(key1FF_keystate_n11) );
  BUF_X1 key1FF_keystate_U6 ( .A(selP), .Z(key1FF_keystate_n16) );
  BUF_X2 key1FF_keystate_U5 ( .A(enKey), .Z(key1FF_keystate_n10) );
  BUF_X1 key1FF_keystate_U4 ( .A(selP), .Z(key1FF_keystate_n15) );
  BUF_X2 key1FF_keystate_U3 ( .A(enKey), .Z(key1FF_keystate_n13) );
  BUF_X1 key1FF_keystate_U2 ( .A(selP), .Z(key1FF_keystate_n14) );
  BUF_X1 key1FF_keystate_U1 ( .A(selP), .Z(key1FF_keystate_n18) );
  OAI21_X1 key1FF_keystate_gff_1_SFF_0_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_1_SFF_0_n8), .A(key1FF_keystate_gff_1_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_1_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_1_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_1_SFF_0_n10), .B2(key1FF_n1), .C1(
        key1FF_keystate_gff_1_SFF_0_n11), .C2(key1FF_outputPar[3]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_1_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_1_SFF_0_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_1_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_1_SFF_0_U2 ( .A(key1FF_keystate_gff_1_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_1_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_1_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_1_SFF_0_n7), .CK(clk), .Q(keyRegKS1[1]), .QN(
        key1FF_keystate_gff_1_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_1_SFF_1_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_1_SFF_1_n8), .A(key1FF_keystate_gff_1_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_1_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_1_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_1_SFF_1_n10), .B2(key1FF_n2), .C1(
        key1FF_keystate_gff_1_SFF_1_n11), .C2(key1FF_outputPar[4]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_1_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_1_SFF_1_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_1_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_1_SFF_1_U2 ( .A(key1FF_keystate_gff_1_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_1_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_1_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_1_SFF_1_n7), .CK(clk), .Q(keyRegKS1[2]), .QN(
        key1FF_keystate_gff_1_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_1_SFF_2_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_1_SFF_2_n8), .A(key1FF_keystate_gff_1_SFF_2_n12), 
        .ZN(key1FF_keystate_gff_1_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_1_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_1_SFF_2_n10), .B2(key1FF_n3), .C1(
        key1FF_keystate_gff_1_SFF_2_n11), .C2(key1FF_outputPar[5]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_1_SFF_2_n12) );
  INV_X1 key1FF_keystate_gff_1_SFF_2_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_1_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_1_SFF_2_U2 ( .A(key1FF_keystate_gff_1_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_1_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_1_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_1_SFF_2_n7), .CK(clk), .Q(keyRegKS1[3]), .QN(
        key1FF_keystate_gff_1_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_1_SFF_3_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_1_SFF_3_n8), .A(key1FF_keystate_gff_1_SFF_3_n12), 
        .ZN(key1FF_keystate_gff_1_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_1_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_1_SFF_3_n10), .B2(key1FF_n4), .C1(
        key1FF_keystate_gff_1_SFF_3_n11), .C2(key1FF_outputPar[6]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_1_SFF_3_n12) );
  INV_X1 key1FF_keystate_gff_1_SFF_3_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_1_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_1_SFF_3_U2 ( .A(key1FF_keystate_gff_1_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_1_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_1_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_1_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[3]), 
        .QN(key1FF_keystate_gff_1_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_2_SFF_0_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_2_SFF_0_n8), .A(key1FF_keystate_gff_2_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_2_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_2_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_2_SFF_0_n10), .B2(keyRegKS1[1]), .C1(
        key1FF_keystate_gff_2_SFF_0_n11), .C2(key1FF_outputPar[7]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_2_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_2_SFF_0_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_2_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_2_SFF_0_U2 ( .A(key1FF_keystate_gff_2_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_2_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_2_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_2_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[4]), 
        .QN(key1FF_keystate_gff_2_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_2_SFF_1_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_2_SFF_1_n8), .A(key1FF_keystate_gff_2_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_2_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_2_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_2_SFF_1_n10), .B2(keyRegKS1[2]), .C1(
        key1FF_keystate_gff_2_SFF_1_n11), .C2(key1FF_outputPar[8]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_2_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_2_SFF_1_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_2_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_2_SFF_1_U2 ( .A(key1FF_keystate_gff_2_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_2_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_2_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_2_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[5]), 
        .QN(key1FF_keystate_gff_2_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_2_SFF_2_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_2_SFF_2_n8), .A(key1FF_keystate_gff_2_SFF_2_n12), 
        .ZN(key1FF_keystate_gff_2_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_2_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_2_SFF_2_n10), .B2(keyRegKS1[3]), .C1(
        key1FF_keystate_gff_2_SFF_2_n11), .C2(key1FF_outputPar[9]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_2_SFF_2_n12) );
  INV_X1 key1FF_keystate_gff_2_SFF_2_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_2_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_2_SFF_2_U2 ( .A(key1FF_keystate_gff_2_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_2_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_2_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_2_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[6]), 
        .QN(key1FF_keystate_gff_2_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_2_SFF_3_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_2_SFF_3_n8), .A(key1FF_keystate_gff_2_SFF_3_n12), 
        .ZN(key1FF_keystate_gff_2_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_2_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_2_SFF_3_n10), .B2(key1FF_outputPar[3]), .C1(
        key1FF_keystate_gff_2_SFF_3_n11), .C2(key1FF_outputPar[10]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_2_SFF_3_n12) );
  INV_X1 key1FF_keystate_gff_2_SFF_3_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_2_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_2_SFF_3_U2 ( .A(key1FF_keystate_gff_2_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_2_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_2_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_2_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[7]), 
        .QN(key1FF_keystate_gff_2_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_3_SFF_0_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_3_SFF_0_n8), .A(key1FF_keystate_gff_3_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_3_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_3_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_3_SFF_0_n10), .B2(key1FF_outputPar[4]), .C1(
        key1FF_keystate_gff_3_SFF_0_n11), .C2(key1FF_outputPar[11]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_3_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_3_SFF_0_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_3_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_3_SFF_0_U2 ( .A(key1FF_keystate_gff_3_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_3_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_3_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_3_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[8]), 
        .QN(key1FF_keystate_gff_3_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_3_SFF_1_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_3_SFF_1_n8), .A(key1FF_keystate_gff_3_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_3_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_3_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_3_SFF_1_n10), .B2(key1FF_outputPar[5]), .C1(
        key1FF_keystate_gff_3_SFF_1_n11), .C2(key1FF_outputPar[12]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_3_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_3_SFF_1_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_3_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_3_SFF_1_U2 ( .A(key1FF_keystate_gff_3_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_3_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_3_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_3_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[9]), 
        .QN(key1FF_keystate_gff_3_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_3_SFF_2_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_3_SFF_2_n7), .A(key1FF_keystate_gff_3_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_3_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_3_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_3_SFF_2_n9), .B2(key1FF_outputPar[6]), .C1(
        key1FF_keystate_gff_3_SFF_2_n10), .C2(key1FF_outputPar[13]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_3_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_3_SFF_2_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_3_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_3_SFF_2_U2 ( .A(key1FF_keystate_gff_3_SFF_2_n10), 
        .ZN(key1FF_keystate_gff_3_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_3_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_3_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[10]), 
        .QN(key1FF_keystate_gff_3_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_3_SFF_3_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_3_SFF_3_n7), .A(key1FF_keystate_gff_3_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_3_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_3_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_3_SFF_3_n9), .B2(key1FF_outputPar[7]), .C1(
        key1FF_keystate_gff_3_SFF_3_n10), .C2(key1FF_outputPar[14]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_3_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_3_SFF_3_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_3_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_3_SFF_3_U2 ( .A(key1FF_keystate_gff_3_SFF_3_n10), 
        .ZN(key1FF_keystate_gff_3_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_3_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_3_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[11]), 
        .QN(key1FF_keystate_gff_3_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_4_SFF_0_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_4_SFF_0_n7), .A(key1FF_keystate_gff_4_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_4_SFF_0_n6) );
  OAI221_X1 key1FF_keystate_gff_4_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_4_SFF_0_n9), .B2(key1FF_outputPar[8]), .C1(
        key1FF_keystate_gff_4_SFF_0_n10), .C2(key1FF_outputPar[15]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_4_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_4_SFF_0_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_4_SFF_0_n10) );
  INV_X1 key1FF_keystate_gff_4_SFF_0_U2 ( .A(key1FF_keystate_gff_4_SFF_0_n10), 
        .ZN(key1FF_keystate_gff_4_SFF_0_n9) );
  DFF_X1 key1FF_keystate_gff_4_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_4_SFF_0_n6), .CK(clk), .Q(key1FF_outputPar[12]), 
        .QN(key1FF_keystate_gff_4_SFF_0_n7) );
  OAI21_X1 key1FF_keystate_gff_4_SFF_1_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_4_SFF_1_n7), .A(key1FF_keystate_gff_4_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_4_SFF_1_n6) );
  OAI221_X1 key1FF_keystate_gff_4_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_4_SFF_1_n9), .B2(key1FF_outputPar[9]), .C1(
        key1FF_keystate_gff_4_SFF_1_n10), .C2(key1FF_outputPar[16]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_4_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_4_SFF_1_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_4_SFF_1_n10) );
  INV_X1 key1FF_keystate_gff_4_SFF_1_U2 ( .A(key1FF_keystate_gff_4_SFF_1_n10), 
        .ZN(key1FF_keystate_gff_4_SFF_1_n9) );
  DFF_X1 key1FF_keystate_gff_4_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_4_SFF_1_n6), .CK(clk), .Q(key1FF_outputPar[13]), 
        .QN(key1FF_keystate_gff_4_SFF_1_n7) );
  OAI21_X1 key1FF_keystate_gff_4_SFF_2_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_4_SFF_2_n7), .A(key1FF_keystate_gff_4_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_4_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_4_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_4_SFF_2_n9), .B2(key1FF_outputPar[10]), .C1(
        key1FF_keystate_gff_4_SFF_2_n10), .C2(key1FF_outputPar[17]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_4_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_4_SFF_2_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_4_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_4_SFF_2_U2 ( .A(key1FF_keystate_gff_4_SFF_2_n10), 
        .ZN(key1FF_keystate_gff_4_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_4_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_4_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[14]), 
        .QN(key1FF_keystate_gff_4_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_4_SFF_3_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_4_SFF_3_n7), .A(key1FF_keystate_gff_4_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_4_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_4_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_4_SFF_3_n9), .B2(key1FF_outputPar[11]), .C1(
        key1FF_keystate_gff_4_SFF_3_n10), .C2(key1FF_counterAdd[0]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_4_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_4_SFF_3_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_4_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_4_SFF_3_U2 ( .A(key1FF_keystate_gff_4_SFF_3_n10), 
        .ZN(key1FF_keystate_gff_4_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_4_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_4_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[15]), 
        .QN(key1FF_keystate_gff_4_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_5_SFF_0_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_5_SFF_0_n8), .A(key1FF_keystate_gff_5_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_5_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_5_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_5_SFF_0_n10), .B2(key1FF_outputPar[12]), .C1(
        key1FF_keystate_gff_5_SFF_0_n11), .C2(key1FF_counterAdd[1]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_5_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_5_SFF_0_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_5_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_5_SFF_0_U2 ( .A(key1FF_keystate_gff_5_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_5_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_5_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_5_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[16]), 
        .QN(key1FF_keystate_gff_5_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_5_SFF_1_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_5_SFF_1_n8), .A(key1FF_keystate_gff_5_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_5_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_5_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_5_SFF_1_n10), .B2(key1FF_outputPar[13]), .C1(
        key1FF_keystate_gff_5_SFF_1_n11), .C2(key1FF_counterAdd[2]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_5_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_5_SFF_1_U3 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_5_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_5_SFF_1_U2 ( .A(key1FF_keystate_gff_5_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_5_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_5_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_5_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[17]), 
        .QN(key1FF_keystate_gff_5_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_5_SFF_2_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_5_SFF_2_n8), .A(key1FF_keystate_gff_5_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_5_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_5_SFF_2_U3 ( .B1(key1FF_keystate_n14), .B2(
        key1FF_outputPar[14]), .C1(key1FF_keystate_gff_5_SFF_2_n10), .C2(
        key1FF_counterAdd[3]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_5_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_5_SFF_2_U2 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_5_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_5_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_5_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[18]), 
        .QN(key1FF_keystate_gff_5_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_5_SFF_3_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_5_SFF_3_n8), .A(key1FF_keystate_gff_5_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_5_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_5_SFF_3_U3 ( .B1(key1FF_keystate_n14), .B2(
        key1FF_outputPar[15]), .C1(key1FF_keystate_gff_5_SFF_3_n10), .C2(
        key1FF_counterAdd[4]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_5_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_5_SFF_3_U2 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_5_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_5_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_5_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[19]), 
        .QN(key1FF_keystate_gff_5_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_6_SFF_0_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_6_SFF_0_n8), .A(key1FF_keystate_gff_6_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_6_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_6_SFF_0_U3 ( .B1(key1FF_keystate_n14), .B2(
        key1FF_outputPar[16]), .C1(key1FF_keystate_gff_6_SFF_0_n10), .C2(
        key1FF_outputPar[23]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_6_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_6_SFF_0_U2 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_6_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_6_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_6_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[20]), 
        .QN(key1FF_keystate_gff_6_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_6_SFF_1_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_6_SFF_1_n8), .A(key1FF_keystate_gff_6_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_6_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_6_SFF_1_U3 ( .B1(key1FF_keystate_n14), .B2(
        key1FF_outputPar[17]), .C1(key1FF_keystate_gff_6_SFF_1_n10), .C2(
        key1FF_outputPar[24]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_6_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_6_SFF_1_U2 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_6_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_6_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_6_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[21]), 
        .QN(key1FF_keystate_gff_6_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_6_SFF_2_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_6_SFF_2_n8), .A(key1FF_keystate_gff_6_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_6_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_6_SFF_2_U3 ( .B1(key1FF_keystate_n14), .B2(
        key1FF_outputPar[18]), .C1(key1FF_keystate_gff_6_SFF_2_n10), .C2(
        key1FF_outputPar[25]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_6_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_6_SFF_2_U2 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_6_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_6_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_6_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[22]), 
        .QN(key1FF_keystate_gff_6_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_6_SFF_3_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_6_SFF_3_n8), .A(key1FF_keystate_gff_6_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_6_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_6_SFF_3_U3 ( .B1(key1FF_keystate_n14), .B2(
        key1FF_outputPar[19]), .C1(key1FF_keystate_gff_6_SFF_3_n10), .C2(
        key1FF_outputPar[26]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_6_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_6_SFF_3_U2 ( .A(key1FF_keystate_n14), .ZN(
        key1FF_keystate_gff_6_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_6_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_6_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[23]), 
        .QN(key1FF_keystate_gff_6_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_7_SFF_0_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_7_SFF_0_n8), .A(key1FF_keystate_gff_7_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_7_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_7_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_7_SFF_0_n10), .B2(key1FF_outputPar[20]), .C1(
        key1FF_keystate_gff_7_SFF_0_n11), .C2(key1FF_outputPar[27]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_7_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_7_SFF_0_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_7_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_7_SFF_0_U2 ( .A(key1FF_keystate_gff_7_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_7_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_7_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_7_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[24]), 
        .QN(key1FF_keystate_gff_7_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_7_SFF_1_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_7_SFF_1_n8), .A(key1FF_keystate_gff_7_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_7_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_7_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_7_SFF_1_n10), .B2(key1FF_outputPar[21]), .C1(
        key1FF_keystate_gff_7_SFF_1_n11), .C2(key1FF_outputPar[28]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_7_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_7_SFF_1_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_7_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_7_SFF_1_U2 ( .A(key1FF_keystate_gff_7_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_7_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_7_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_7_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[25]), 
        .QN(key1FF_keystate_gff_7_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_7_SFF_2_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_7_SFF_2_n7), .A(key1FF_keystate_gff_7_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_7_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_7_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_7_SFF_2_n9), .B2(key1FF_outputPar[22]), .C1(
        key1FF_keystate_gff_7_SFF_2_n10), .C2(key1FF_outputPar[29]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_7_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_7_SFF_2_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_7_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_7_SFF_2_U2 ( .A(key1FF_keystate_gff_7_SFF_2_n10), 
        .ZN(key1FF_keystate_gff_7_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_7_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_7_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[26]), 
        .QN(key1FF_keystate_gff_7_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_7_SFF_3_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_7_SFF_3_n7), .A(key1FF_keystate_gff_7_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_7_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_7_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_7_SFF_3_n9), .B2(key1FF_outputPar[23]), .C1(
        key1FF_keystate_gff_7_SFF_3_n10), .C2(key1FF_outputPar[30]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_7_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_7_SFF_3_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_7_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_7_SFF_3_U2 ( .A(key1FF_keystate_gff_7_SFF_3_n10), 
        .ZN(key1FF_keystate_gff_7_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_7_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_7_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[27]), 
        .QN(key1FF_keystate_gff_7_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_8_SFF_0_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_8_SFF_0_n7), .A(key1FF_keystate_gff_8_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_8_SFF_0_n6) );
  OAI221_X1 key1FF_keystate_gff_8_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_8_SFF_0_n9), .B2(key1FF_outputPar[24]), .C1(
        key1FF_keystate_gff_8_SFF_0_n10), .C2(key1FF_outputPar[31]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_8_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_8_SFF_0_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_8_SFF_0_n10) );
  INV_X1 key1FF_keystate_gff_8_SFF_0_U2 ( .A(key1FF_keystate_gff_8_SFF_0_n10), 
        .ZN(key1FF_keystate_gff_8_SFF_0_n9) );
  DFF_X1 key1FF_keystate_gff_8_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_8_SFF_0_n6), .CK(clk), .Q(key1FF_outputPar[28]), 
        .QN(key1FF_keystate_gff_8_SFF_0_n7) );
  OAI21_X1 key1FF_keystate_gff_8_SFF_1_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_8_SFF_1_n7), .A(key1FF_keystate_gff_8_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_8_SFF_1_n6) );
  OAI221_X1 key1FF_keystate_gff_8_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_8_SFF_1_n9), .B2(key1FF_outputPar[25]), .C1(
        key1FF_keystate_gff_8_SFF_1_n10), .C2(key1FF_outputPar[32]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_8_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_8_SFF_1_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_8_SFF_1_n10) );
  INV_X1 key1FF_keystate_gff_8_SFF_1_U2 ( .A(key1FF_keystate_gff_8_SFF_1_n10), 
        .ZN(key1FF_keystate_gff_8_SFF_1_n9) );
  DFF_X1 key1FF_keystate_gff_8_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_8_SFF_1_n6), .CK(clk), .Q(key1FF_outputPar[29]), 
        .QN(key1FF_keystate_gff_8_SFF_1_n7) );
  OAI21_X1 key1FF_keystate_gff_8_SFF_2_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_8_SFF_2_n7), .A(key1FF_keystate_gff_8_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_8_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_8_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_8_SFF_2_n9), .B2(key1FF_outputPar[26]), .C1(
        key1FF_keystate_gff_8_SFF_2_n10), .C2(key1FF_outputPar[33]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_8_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_8_SFF_2_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_8_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_8_SFF_2_U2 ( .A(key1FF_keystate_gff_8_SFF_2_n10), 
        .ZN(key1FF_keystate_gff_8_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_8_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_8_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[30]), 
        .QN(key1FF_keystate_gff_8_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_8_SFF_3_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_8_SFF_3_n7), .A(key1FF_keystate_gff_8_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_8_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_8_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_8_SFF_3_n9), .B2(key1FF_outputPar[27]), .C1(
        key1FF_keystate_gff_8_SFF_3_n10), .C2(key1FF_outputPar[34]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_8_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_8_SFF_3_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_8_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_8_SFF_3_U2 ( .A(key1FF_keystate_gff_8_SFF_3_n10), 
        .ZN(key1FF_keystate_gff_8_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_8_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_8_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[31]), 
        .QN(key1FF_keystate_gff_8_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_9_SFF_0_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_9_SFF_0_n8), .A(key1FF_keystate_gff_9_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_9_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_9_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_9_SFF_0_n10), .B2(key1FF_outputPar[28]), .C1(
        key1FF_keystate_gff_9_SFF_0_n11), .C2(key1FF_outputPar[35]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_9_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_9_SFF_0_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_9_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_9_SFF_0_U2 ( .A(key1FF_keystate_gff_9_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_9_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_9_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_9_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[32]), 
        .QN(key1FF_keystate_gff_9_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_9_SFF_1_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_9_SFF_1_n8), .A(key1FF_keystate_gff_9_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_9_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_9_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_9_SFF_1_n10), .B2(key1FF_outputPar[29]), .C1(
        key1FF_keystate_gff_9_SFF_1_n11), .C2(key1FF_outputPar[36]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_9_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_9_SFF_1_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_9_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_9_SFF_1_U2 ( .A(key1FF_keystate_gff_9_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_9_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_9_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_9_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[33]), 
        .QN(key1FF_keystate_gff_9_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_9_SFF_2_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_9_SFF_2_n8), .A(key1FF_keystate_gff_9_SFF_2_n12), 
        .ZN(key1FF_keystate_gff_9_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_9_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_9_SFF_2_n10), .B2(key1FF_outputPar[30]), .C1(
        key1FF_keystate_gff_9_SFF_2_n11), .C2(key1FF_outputPar[37]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_9_SFF_2_n12) );
  INV_X1 key1FF_keystate_gff_9_SFF_2_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_9_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_9_SFF_2_U2 ( .A(key1FF_keystate_gff_9_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_9_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_9_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_9_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[34]), 
        .QN(key1FF_keystate_gff_9_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_9_SFF_3_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_9_SFF_3_n8), .A(key1FF_keystate_gff_9_SFF_3_n12), 
        .ZN(key1FF_keystate_gff_9_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_9_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_9_SFF_3_n10), .B2(key1FF_outputPar[31]), .C1(
        key1FF_keystate_gff_9_SFF_3_n11), .C2(key1FF_outputPar[38]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_9_SFF_3_n12) );
  INV_X1 key1FF_keystate_gff_9_SFF_3_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_9_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_9_SFF_3_U2 ( .A(key1FF_keystate_gff_9_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_9_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_9_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_9_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[35]), 
        .QN(key1FF_keystate_gff_9_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_10_SFF_0_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_10_SFF_0_n8), .A(key1FF_keystate_gff_10_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_10_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_10_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_10_SFF_0_n10), .B2(key1FF_outputPar[32]), .C1(
        key1FF_keystate_gff_10_SFF_0_n11), .C2(key1FF_outputPar[39]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_10_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_10_SFF_0_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_10_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_10_SFF_0_U2 ( .A(key1FF_keystate_gff_10_SFF_0_n11), .ZN(key1FF_keystate_gff_10_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_10_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_10_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[36]), 
        .QN(key1FF_keystate_gff_10_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_10_SFF_1_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_10_SFF_1_n8), .A(key1FF_keystate_gff_10_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_10_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_10_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_10_SFF_1_n10), .B2(key1FF_outputPar[33]), .C1(
        key1FF_keystate_gff_10_SFF_1_n11), .C2(key1FF_outputPar[40]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_10_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_10_SFF_1_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_10_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_10_SFF_1_U2 ( .A(key1FF_keystate_gff_10_SFF_1_n11), .ZN(key1FF_keystate_gff_10_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_10_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_10_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[37]), 
        .QN(key1FF_keystate_gff_10_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_10_SFF_2_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_10_SFF_2_n8), .A(key1FF_keystate_gff_10_SFF_2_n12), 
        .ZN(key1FF_keystate_gff_10_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_10_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_10_SFF_2_n10), .B2(key1FF_outputPar[34]), .C1(
        key1FF_keystate_gff_10_SFF_2_n11), .C2(key1FF_outputPar[41]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_10_SFF_2_n12) );
  INV_X1 key1FF_keystate_gff_10_SFF_2_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_10_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_10_SFF_2_U2 ( .A(key1FF_keystate_gff_10_SFF_2_n11), .ZN(key1FF_keystate_gff_10_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_10_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_10_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[38]), 
        .QN(key1FF_keystate_gff_10_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_10_SFF_3_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_10_SFF_3_n8), .A(key1FF_keystate_gff_10_SFF_3_n12), 
        .ZN(key1FF_keystate_gff_10_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_10_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_10_SFF_3_n10), .B2(key1FF_outputPar[35]), .C1(
        key1FF_keystate_gff_10_SFF_3_n11), .C2(key1FF_outputPar[42]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_10_SFF_3_n12) );
  INV_X1 key1FF_keystate_gff_10_SFF_3_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_10_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_10_SFF_3_U2 ( .A(key1FF_keystate_gff_10_SFF_3_n11), .ZN(key1FF_keystate_gff_10_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_10_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_10_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[39]), 
        .QN(key1FF_keystate_gff_10_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_11_SFF_0_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_11_SFF_0_n8), .A(key1FF_keystate_gff_11_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_11_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_11_SFF_0_U3 ( .B1(key1FF_keystate_n17), .B2(
        key1FF_outputPar[36]), .C1(key1FF_keystate_gff_11_SFF_0_n10), .C2(
        key1FF_outputPar[43]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_11_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_11_SFF_0_U2 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_11_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_11_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_11_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[40]), 
        .QN(key1FF_keystate_gff_11_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_11_SFF_1_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_11_SFF_1_n8), .A(key1FF_keystate_gff_11_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_11_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_11_SFF_1_U3 ( .B1(key1FF_keystate_n17), .B2(
        key1FF_outputPar[37]), .C1(key1FF_keystate_gff_11_SFF_1_n10), .C2(
        key1FF_outputPar[44]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_11_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_11_SFF_1_U2 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_11_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_11_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_11_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[41]), 
        .QN(key1FF_keystate_gff_11_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_11_SFF_2_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_11_SFF_2_n7), .A(key1FF_keystate_gff_11_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_11_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_11_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_11_SFF_2_n9), .B2(key1FF_outputPar[38]), .C1(
        key1FF_keystate_gff_11_SFF_2_n10), .C2(key1FF_outputPar[45]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_11_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_11_SFF_2_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_11_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_11_SFF_2_U2 ( .A(key1FF_keystate_gff_11_SFF_2_n10), .ZN(key1FF_keystate_gff_11_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_11_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_11_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[42]), 
        .QN(key1FF_keystate_gff_11_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_11_SFF_3_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_11_SFF_3_n7), .A(key1FF_keystate_gff_11_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_11_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_11_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_11_SFF_3_n9), .B2(key1FF_outputPar[39]), .C1(
        key1FF_keystate_gff_11_SFF_3_n10), .C2(key1FF_outputPar[46]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_11_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_11_SFF_3_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_11_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_11_SFF_3_U2 ( .A(key1FF_keystate_gff_11_SFF_3_n10), .ZN(key1FF_keystate_gff_11_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_11_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_11_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[43]), 
        .QN(key1FF_keystate_gff_11_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_12_SFF_0_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_12_SFF_0_n7), .A(key1FF_keystate_gff_12_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_12_SFF_0_n6) );
  OAI221_X1 key1FF_keystate_gff_12_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_12_SFF_0_n9), .B2(key1FF_outputPar[40]), .C1(
        key1FF_keystate_gff_12_SFF_0_n10), .C2(key1FF_outputPar[47]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_12_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_12_SFF_0_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_12_SFF_0_n10) );
  INV_X1 key1FF_keystate_gff_12_SFF_0_U2 ( .A(key1FF_keystate_gff_12_SFF_0_n10), .ZN(key1FF_keystate_gff_12_SFF_0_n9) );
  DFF_X1 key1FF_keystate_gff_12_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_12_SFF_0_n6), .CK(clk), .Q(key1FF_outputPar[44]), 
        .QN(key1FF_keystate_gff_12_SFF_0_n7) );
  OAI21_X1 key1FF_keystate_gff_12_SFF_1_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_12_SFF_1_n7), .A(key1FF_keystate_gff_12_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_12_SFF_1_n6) );
  OAI221_X1 key1FF_keystate_gff_12_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_12_SFF_1_n9), .B2(key1FF_outputPar[41]), .C1(
        key1FF_keystate_gff_12_SFF_1_n10), .C2(key1FF_outputPar[48]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_12_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_12_SFF_1_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_12_SFF_1_n10) );
  INV_X1 key1FF_keystate_gff_12_SFF_1_U2 ( .A(key1FF_keystate_gff_12_SFF_1_n10), .ZN(key1FF_keystate_gff_12_SFF_1_n9) );
  DFF_X1 key1FF_keystate_gff_12_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_12_SFF_1_n6), .CK(clk), .Q(key1FF_outputPar[45]), 
        .QN(key1FF_keystate_gff_12_SFF_1_n7) );
  OAI21_X1 key1FF_keystate_gff_12_SFF_2_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_12_SFF_2_n7), .A(key1FF_keystate_gff_12_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_12_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_12_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_12_SFF_2_n9), .B2(key1FF_outputPar[42]), .C1(
        key1FF_keystate_gff_12_SFF_2_n10), .C2(key1FF_outputPar[49]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_12_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_12_SFF_2_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_12_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_12_SFF_2_U2 ( .A(key1FF_keystate_gff_12_SFF_2_n10), .ZN(key1FF_keystate_gff_12_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_12_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_12_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[46]), 
        .QN(key1FF_keystate_gff_12_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_12_SFF_3_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_12_SFF_3_n7), .A(key1FF_keystate_gff_12_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_12_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_12_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_12_SFF_3_n9), .B2(key1FF_outputPar[43]), .C1(
        key1FF_keystate_gff_12_SFF_3_n10), .C2(key1FF_outputPar[50]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_12_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_12_SFF_3_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_12_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_12_SFF_3_U2 ( .A(key1FF_keystate_gff_12_SFF_3_n10), .ZN(key1FF_keystate_gff_12_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_12_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_12_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[47]), 
        .QN(key1FF_keystate_gff_12_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_13_SFF_0_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_13_SFF_0_n8), .A(key1FF_keystate_gff_13_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_13_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_13_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_13_SFF_0_n10), .B2(key1FF_outputPar[44]), .C1(
        key1FF_keystate_gff_13_SFF_0_n11), .C2(key1FF_outputPar[51]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_13_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_13_SFF_0_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_13_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_13_SFF_0_U2 ( .A(key1FF_keystate_gff_13_SFF_0_n11), .ZN(key1FF_keystate_gff_13_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_13_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_13_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[48]), 
        .QN(key1FF_keystate_gff_13_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_13_SFF_1_U5 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_13_SFF_1_n8), .A(key1FF_keystate_gff_13_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_13_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_13_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_13_SFF_1_n10), .B2(key1FF_outputPar[45]), .C1(
        key1FF_keystate_gff_13_SFF_1_n11), .C2(key1FF_outputPar[52]), .A(
        key1FF_keystate_n10), .ZN(key1FF_keystate_gff_13_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_13_SFF_1_U3 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_13_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_13_SFF_1_U2 ( .A(key1FF_keystate_gff_13_SFF_1_n11), .ZN(key1FF_keystate_gff_13_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_13_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_13_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[49]), 
        .QN(key1FF_keystate_gff_13_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_13_SFF_2_U4 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_13_SFF_2_n8), .A(key1FF_keystate_gff_13_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_13_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_13_SFF_2_U3 ( .B1(key1FF_keystate_n15), .B2(
        key1FF_outputPar[46]), .C1(key1FF_keystate_gff_13_SFF_2_n10), .C2(
        key1FF_outputPar[53]), .A(key1FF_keystate_n10), .ZN(
        key1FF_keystate_gff_13_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_13_SFF_2_U2 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_13_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_13_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_13_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[50]), 
        .QN(key1FF_keystate_gff_13_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_13_SFF_3_U4 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_13_SFF_3_n8), .A(key1FF_keystate_gff_13_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_13_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_13_SFF_3_U3 ( .B1(key1FF_keystate_n15), .B2(
        key1FF_outputPar[47]), .C1(key1FF_keystate_gff_13_SFF_3_n10), .C2(
        key1FF_outputPar[54]), .A(key1FF_keystate_n10), .ZN(
        key1FF_keystate_gff_13_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_13_SFF_3_U2 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_13_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_13_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_13_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[51]), 
        .QN(key1FF_keystate_gff_13_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_14_SFF_0_U4 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_14_SFF_0_n8), .A(key1FF_keystate_gff_14_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_14_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_14_SFF_0_U3 ( .B1(key1FF_keystate_n15), .B2(
        key1FF_outputPar[48]), .C1(key1FF_keystate_gff_14_SFF_0_n10), .C2(
        key1FF_outputPar[55]), .A(key1FF_keystate_n10), .ZN(
        key1FF_keystate_gff_14_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_14_SFF_0_U2 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_14_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_14_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_14_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[52]), 
        .QN(key1FF_keystate_gff_14_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_14_SFF_1_U4 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_14_SFF_1_n8), .A(key1FF_keystate_gff_14_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_14_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_14_SFF_1_U3 ( .B1(key1FF_keystate_n15), .B2(
        key1FF_outputPar[49]), .C1(key1FF_keystate_gff_14_SFF_1_n10), .C2(
        key1FF_outputPar[56]), .A(key1FF_keystate_n10), .ZN(
        key1FF_keystate_gff_14_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_14_SFF_1_U2 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_14_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_14_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_14_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[53]), 
        .QN(key1FF_keystate_gff_14_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_14_SFF_2_U4 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_14_SFF_2_n8), .A(key1FF_keystate_gff_14_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_14_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_14_SFF_2_U3 ( .B1(key1FF_keystate_n15), .B2(
        key1FF_outputPar[50]), .C1(key1FF_keystate_gff_14_SFF_2_n10), .C2(
        key1FF_outputPar[57]), .A(key1FF_keystate_n10), .ZN(
        key1FF_keystate_gff_14_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_14_SFF_2_U2 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_14_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_14_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_14_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[54]), 
        .QN(key1FF_keystate_gff_14_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_14_SFF_3_U4 ( .B1(key1FF_keystate_n10), .B2(
        key1FF_keystate_gff_14_SFF_3_n8), .A(key1FF_keystate_gff_14_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_14_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_14_SFF_3_U3 ( .B1(key1FF_keystate_n15), .B2(
        key1FF_outputPar[51]), .C1(key1FF_keystate_gff_14_SFF_3_n10), .C2(
        key1FF_outputPar[58]), .A(key1FF_keystate_n10), .ZN(
        key1FF_keystate_gff_14_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_14_SFF_3_U2 ( .A(key1FF_keystate_n15), .ZN(
        key1FF_keystate_gff_14_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_14_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_14_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[55]), 
        .QN(key1FF_keystate_gff_14_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_15_SFF_0_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_15_SFF_0_n8), .A(key1FF_keystate_gff_15_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_15_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_15_SFF_0_U3 ( .B1(key1FF_keystate_n17), .B2(
        key1FF_outputPar[52]), .C1(key1FF_keystate_gff_15_SFF_0_n10), .C2(
        key1FF_outputPar[59]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_15_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_15_SFF_0_U2 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_15_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_15_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_15_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[56]), 
        .QN(key1FF_keystate_gff_15_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_15_SFF_1_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_15_SFF_1_n8), .A(key1FF_keystate_gff_15_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_15_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_15_SFF_1_U3 ( .B1(key1FF_keystate_n17), .B2(
        key1FF_outputPar[53]), .C1(key1FF_keystate_gff_15_SFF_1_n10), .C2(
        key1FF_outputPar[60]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_15_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_15_SFF_1_U2 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_15_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_15_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_15_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[57]), 
        .QN(key1FF_keystate_gff_15_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_15_SFF_2_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_15_SFF_2_n7), .A(key1FF_keystate_gff_15_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_15_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_15_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_15_SFF_2_n9), .B2(key1FF_outputPar[54]), .C1(
        key1FF_keystate_gff_15_SFF_2_n10), .C2(key1FF_outputPar[61]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_15_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_15_SFF_2_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_15_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_15_SFF_2_U2 ( .A(key1FF_keystate_gff_15_SFF_2_n10), .ZN(key1FF_keystate_gff_15_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_15_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_15_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[58]), 
        .QN(key1FF_keystate_gff_15_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_15_SFF_3_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_15_SFF_3_n7), .A(key1FF_keystate_gff_15_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_15_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_15_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_15_SFF_3_n9), .B2(key1FF_outputPar[55]), .C1(
        key1FF_keystate_gff_15_SFF_3_n10), .C2(key1FF_outputPar[62]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_15_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_15_SFF_3_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_15_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_15_SFF_3_U2 ( .A(key1FF_keystate_gff_15_SFF_3_n10), .ZN(key1FF_keystate_gff_15_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_15_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_15_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[59]), 
        .QN(key1FF_keystate_gff_15_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_16_SFF_0_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_16_SFF_0_n7), .A(key1FF_keystate_gff_16_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_16_SFF_0_n6) );
  OAI221_X1 key1FF_keystate_gff_16_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_16_SFF_0_n9), .B2(key1FF_outputPar[56]), .C1(
        key1FF_keystate_gff_16_SFF_0_n10), .C2(key1FF_outputPar[63]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_16_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_16_SFF_0_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_16_SFF_0_n10) );
  INV_X1 key1FF_keystate_gff_16_SFF_0_U2 ( .A(key1FF_keystate_gff_16_SFF_0_n10), .ZN(key1FF_keystate_gff_16_SFF_0_n9) );
  DFF_X1 key1FF_keystate_gff_16_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_16_SFF_0_n6), .CK(clk), .Q(key1FF_outputPar[60]), 
        .QN(key1FF_keystate_gff_16_SFF_0_n7) );
  OAI21_X1 key1FF_keystate_gff_16_SFF_1_U5 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_16_SFF_1_n7), .A(key1FF_keystate_gff_16_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_16_SFF_1_n6) );
  OAI221_X1 key1FF_keystate_gff_16_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_16_SFF_1_n9), .B2(key1FF_outputPar[57]), .C1(
        key1FF_keystate_gff_16_SFF_1_n10), .C2(key1FF_outputPar[64]), .A(
        key1FF_keystate_n13), .ZN(key1FF_keystate_gff_16_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_16_SFF_1_U3 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_16_SFF_1_n10) );
  INV_X1 key1FF_keystate_gff_16_SFF_1_U2 ( .A(key1FF_keystate_gff_16_SFF_1_n10), .ZN(key1FF_keystate_gff_16_SFF_1_n9) );
  DFF_X1 key1FF_keystate_gff_16_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_16_SFF_1_n6), .CK(clk), .Q(key1FF_outputPar[61]), 
        .QN(key1FF_keystate_gff_16_SFF_1_n7) );
  OAI21_X1 key1FF_keystate_gff_16_SFF_2_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_16_SFF_2_n7), .A(key1FF_keystate_gff_16_SFF_2_n10), 
        .ZN(key1FF_keystate_gff_16_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_16_SFF_2_U3 ( .B1(key1FF_keystate_n18), .B2(
        key1FF_outputPar[58]), .C1(key1FF_keystate_gff_16_SFF_2_n9), .C2(
        key1FF_outputPar[65]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_16_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_16_SFF_2_U2 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_16_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_16_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_16_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[62]), 
        .QN(key1FF_keystate_gff_16_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_16_SFF_3_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_16_SFF_3_n7), .A(key1FF_keystate_gff_16_SFF_3_n10), 
        .ZN(key1FF_keystate_gff_16_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_16_SFF_3_U3 ( .B1(key1FF_keystate_n18), .B2(
        key1FF_outputPar[59]), .C1(key1FF_keystate_gff_16_SFF_3_n9), .C2(
        key1FF_outputPar[66]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_16_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_16_SFF_3_U2 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_16_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_16_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_16_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[63]), 
        .QN(key1FF_keystate_gff_16_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_17_SFF_0_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_17_SFF_0_n8), .A(key1FF_keystate_gff_17_SFF_0_n12), 
        .ZN(key1FF_keystate_gff_17_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_17_SFF_0_U4 ( .B1(
        key1FF_keystate_gff_17_SFF_0_n10), .B2(key1FF_outputPar[60]), .C1(
        key1FF_keystate_gff_17_SFF_0_n11), .C2(key1FF_outputPar[67]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_17_SFF_0_n12) );
  INV_X1 key1FF_keystate_gff_17_SFF_0_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_17_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_17_SFF_0_U2 ( .A(key1FF_keystate_gff_17_SFF_0_n11), .ZN(key1FF_keystate_gff_17_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_17_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_17_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[64]), 
        .QN(key1FF_keystate_gff_17_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_17_SFF_1_U5 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_17_SFF_1_n8), .A(key1FF_keystate_gff_17_SFF_1_n12), 
        .ZN(key1FF_keystate_gff_17_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_17_SFF_1_U4 ( .B1(
        key1FF_keystate_gff_17_SFF_1_n10), .B2(key1FF_outputPar[61]), .C1(
        key1FF_keystate_gff_17_SFF_1_n11), .C2(key1FF_outputPar[68]), .A(
        key1FF_keystate_n11), .ZN(key1FF_keystate_gff_17_SFF_1_n12) );
  INV_X1 key1FF_keystate_gff_17_SFF_1_U3 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_17_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_17_SFF_1_U2 ( .A(key1FF_keystate_gff_17_SFF_1_n11), .ZN(key1FF_keystate_gff_17_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_17_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_17_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[65]), 
        .QN(key1FF_keystate_gff_17_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_17_SFF_2_U4 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_17_SFF_2_n8), .A(key1FF_keystate_gff_17_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_17_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_17_SFF_2_U3 ( .B1(key1FF_keystate_n16), .B2(
        key1FF_outputPar[62]), .C1(key1FF_keystate_gff_17_SFF_2_n10), .C2(
        key1FF_outputPar[69]), .A(key1FF_keystate_n11), .ZN(
        key1FF_keystate_gff_17_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_17_SFF_2_U2 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_17_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_17_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_17_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[66]), 
        .QN(key1FF_keystate_gff_17_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_17_SFF_3_U4 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_17_SFF_3_n8), .A(key1FF_keystate_gff_17_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_17_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_17_SFF_3_U3 ( .B1(key1FF_keystate_n16), .B2(
        key1FF_outputPar[63]), .C1(key1FF_keystate_gff_17_SFF_3_n10), .C2(
        key1FF_outputPar[70]), .A(key1FF_keystate_n11), .ZN(
        key1FF_keystate_gff_17_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_17_SFF_3_U2 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_17_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_17_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_17_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[67]), 
        .QN(key1FF_keystate_gff_17_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_18_SFF_0_U4 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_18_SFF_0_n8), .A(key1FF_keystate_gff_18_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_18_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_18_SFF_0_U3 ( .B1(key1FF_keystate_n16), .B2(
        key1FF_outputPar[64]), .C1(key1FF_keystate_gff_18_SFF_0_n10), .C2(
        key1FF_outputPar[71]), .A(key1FF_keystate_n11), .ZN(
        key1FF_keystate_gff_18_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_18_SFF_0_U2 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_18_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_18_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_18_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[68]), 
        .QN(key1FF_keystate_gff_18_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_18_SFF_1_U4 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_18_SFF_1_n8), .A(key1FF_keystate_gff_18_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_18_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_18_SFF_1_U3 ( .B1(key1FF_keystate_n16), .B2(
        key1FF_outputPar[65]), .C1(key1FF_keystate_gff_18_SFF_1_n10), .C2(
        key1FF_outputPar[72]), .A(key1FF_keystate_n11), .ZN(
        key1FF_keystate_gff_18_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_18_SFF_1_U2 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_18_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_18_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_18_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[69]), 
        .QN(key1FF_keystate_gff_18_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_18_SFF_2_U4 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_18_SFF_2_n8), .A(key1FF_keystate_gff_18_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_18_SFF_2_n7) );
  OAI221_X1 key1FF_keystate_gff_18_SFF_2_U3 ( .B1(key1FF_keystate_n16), .B2(
        key1FF_outputPar[66]), .C1(key1FF_keystate_gff_18_SFF_2_n10), .C2(
        key1FF_outputPar[73]), .A(key1FF_keystate_n11), .ZN(
        key1FF_keystate_gff_18_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_18_SFF_2_U2 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_18_SFF_2_n10) );
  DFF_X1 key1FF_keystate_gff_18_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_18_SFF_2_n7), .CK(clk), .Q(key1FF_outputPar[70]), 
        .QN(key1FF_keystate_gff_18_SFF_2_n8) );
  OAI21_X1 key1FF_keystate_gff_18_SFF_3_U4 ( .B1(key1FF_keystate_n11), .B2(
        key1FF_keystate_gff_18_SFF_3_n8), .A(key1FF_keystate_gff_18_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_18_SFF_3_n7) );
  OAI221_X1 key1FF_keystate_gff_18_SFF_3_U3 ( .B1(key1FF_keystate_n16), .B2(
        key1FF_outputPar[67]), .C1(key1FF_keystate_gff_18_SFF_3_n10), .C2(
        key1FF_outputPar[74]), .A(key1FF_keystate_n11), .ZN(
        key1FF_keystate_gff_18_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_18_SFF_3_U2 ( .A(key1FF_keystate_n16), .ZN(
        key1FF_keystate_gff_18_SFF_3_n10) );
  DFF_X1 key1FF_keystate_gff_18_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_18_SFF_3_n7), .CK(clk), .Q(key1FF_outputPar[71]), 
        .QN(key1FF_keystate_gff_18_SFF_3_n8) );
  OAI21_X1 key1FF_keystate_gff_19_SFF_0_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_19_SFF_0_n8), .A(key1FF_keystate_gff_19_SFF_0_n11), 
        .ZN(key1FF_keystate_gff_19_SFF_0_n7) );
  OAI221_X1 key1FF_keystate_gff_19_SFF_0_U3 ( .B1(key1FF_keystate_n17), .B2(
        key1FF_outputPar[68]), .C1(key1FF_keystate_gff_19_SFF_0_n10), .C2(
        key1FF_outputPar[75]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_19_SFF_0_n11) );
  INV_X1 key1FF_keystate_gff_19_SFF_0_U2 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_19_SFF_0_n10) );
  DFF_X1 key1FF_keystate_gff_19_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_19_SFF_0_n7), .CK(clk), .Q(key1FF_outputPar[72]), 
        .QN(key1FF_keystate_gff_19_SFF_0_n8) );
  OAI21_X1 key1FF_keystate_gff_19_SFF_1_U4 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_19_SFF_1_n8), .A(key1FF_keystate_gff_19_SFF_1_n11), 
        .ZN(key1FF_keystate_gff_19_SFF_1_n7) );
  OAI221_X1 key1FF_keystate_gff_19_SFF_1_U3 ( .B1(key1FF_keystate_n17), .B2(
        key1FF_outputPar[69]), .C1(key1FF_keystate_gff_19_SFF_1_n10), .C2(
        roundkey1[0]), .A(key1FF_keystate_n12), .ZN(
        key1FF_keystate_gff_19_SFF_1_n11) );
  INV_X1 key1FF_keystate_gff_19_SFF_1_U2 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_19_SFF_1_n10) );
  DFF_X1 key1FF_keystate_gff_19_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_19_SFF_1_n7), .CK(clk), .Q(key1FF_outputPar[73]), 
        .QN(key1FF_keystate_gff_19_SFF_1_n8) );
  OAI21_X1 key1FF_keystate_gff_19_SFF_2_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_19_SFF_2_n7), .A(key1FF_keystate_gff_19_SFF_2_n11), 
        .ZN(key1FF_keystate_gff_19_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_19_SFF_2_U4 ( .B1(
        key1FF_keystate_gff_19_SFF_2_n9), .B2(key1FF_outputPar[70]), .C1(
        key1FF_keystate_gff_19_SFF_2_n10), .C2(roundkey1[1]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_19_SFF_2_n11) );
  INV_X1 key1FF_keystate_gff_19_SFF_2_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_19_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_19_SFF_2_U2 ( .A(key1FF_keystate_gff_19_SFF_2_n10), .ZN(key1FF_keystate_gff_19_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_19_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_19_SFF_2_n6), .CK(clk), .Q(key1FF_outputPar[74]), 
        .QN(key1FF_keystate_gff_19_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_19_SFF_3_U5 ( .B1(key1FF_keystate_n12), .B2(
        key1FF_keystate_gff_19_SFF_3_n7), .A(key1FF_keystate_gff_19_SFF_3_n11), 
        .ZN(key1FF_keystate_gff_19_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_19_SFF_3_U4 ( .B1(
        key1FF_keystate_gff_19_SFF_3_n9), .B2(key1FF_outputPar[71]), .C1(
        key1FF_keystate_gff_19_SFF_3_n10), .C2(roundkey1[2]), .A(
        key1FF_keystate_n12), .ZN(key1FF_keystate_gff_19_SFF_3_n11) );
  INV_X1 key1FF_keystate_gff_19_SFF_3_U3 ( .A(key1FF_keystate_n17), .ZN(
        key1FF_keystate_gff_19_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_19_SFF_3_U2 ( .A(key1FF_keystate_gff_19_SFF_3_n10), .ZN(key1FF_keystate_gff_19_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_19_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_19_SFF_3_n6), .CK(clk), .Q(key1FF_outputPar[75]), 
        .QN(key1FF_keystate_gff_19_SFF_3_n7) );
  OAI21_X1 key1FF_keystate_gff_20_SFF_0_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_20_SFF_0_n7), .A(key1FF_keystate_gff_20_SFF_0_n10), 
        .ZN(key1FF_keystate_gff_20_SFF_0_n6) );
  OAI221_X1 key1FF_keystate_gff_20_SFF_0_U3 ( .B1(key1FF_keystate_n18), .B2(
        key1FF_outputPar[72]), .C1(key1FF_keystate_gff_20_SFF_0_n9), .C2(
        sboxOut1[0]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_20_SFF_0_n10) );
  INV_X1 key1FF_keystate_gff_20_SFF_0_U2 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_20_SFF_0_n9) );
  DFF_X1 key1FF_keystate_gff_20_SFF_0_Cell_reg ( .D(
        key1FF_keystate_gff_20_SFF_0_n6), .CK(clk), .Q(roundkey1[0]), .QN(
        key1FF_keystate_gff_20_SFF_0_n7) );
  OAI21_X1 key1FF_keystate_gff_20_SFF_1_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_20_SFF_1_n7), .A(key1FF_keystate_gff_20_SFF_1_n10), 
        .ZN(key1FF_keystate_gff_20_SFF_1_n6) );
  OAI221_X1 key1FF_keystate_gff_20_SFF_1_U3 ( .B1(key1FF_keystate_n18), .B2(
        key1FF_outputPar[73]), .C1(key1FF_keystate_gff_20_SFF_1_n9), .C2(
        sboxOut1[1]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_20_SFF_1_n10) );
  INV_X1 key1FF_keystate_gff_20_SFF_1_U2 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_20_SFF_1_n9) );
  DFF_X1 key1FF_keystate_gff_20_SFF_1_Cell_reg ( .D(
        key1FF_keystate_gff_20_SFF_1_n6), .CK(clk), .Q(roundkey1[1]), .QN(
        key1FF_keystate_gff_20_SFF_1_n7) );
  OAI21_X1 key1FF_keystate_gff_20_SFF_2_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_20_SFF_2_n7), .A(key1FF_keystate_gff_20_SFF_2_n10), 
        .ZN(key1FF_keystate_gff_20_SFF_2_n6) );
  OAI221_X1 key1FF_keystate_gff_20_SFF_2_U3 ( .B1(key1FF_keystate_n18), .B2(
        key1FF_outputPar[74]), .C1(key1FF_keystate_gff_20_SFF_2_n9), .C2(
        sboxOut1[2]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_20_SFF_2_n10) );
  INV_X1 key1FF_keystate_gff_20_SFF_2_U2 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_20_SFF_2_n9) );
  DFF_X1 key1FF_keystate_gff_20_SFF_2_Cell_reg ( .D(
        key1FF_keystate_gff_20_SFF_2_n6), .CK(clk), .Q(roundkey1[2]), .QN(
        key1FF_keystate_gff_20_SFF_2_n7) );
  OAI21_X1 key1FF_keystate_gff_20_SFF_3_U4 ( .B1(key1FF_keystate_n13), .B2(
        key1FF_keystate_gff_20_SFF_3_n7), .A(key1FF_keystate_gff_20_SFF_3_n10), 
        .ZN(key1FF_keystate_gff_20_SFF_3_n6) );
  OAI221_X1 key1FF_keystate_gff_20_SFF_3_U3 ( .B1(key1FF_keystate_n18), .B2(
        key1FF_outputPar[75]), .C1(key1FF_keystate_gff_20_SFF_3_n9), .C2(
        sboxOut1[3]), .A(key1FF_keystate_n13), .ZN(
        key1FF_keystate_gff_20_SFF_3_n10) );
  INV_X1 key1FF_keystate_gff_20_SFF_3_U2 ( .A(key1FF_keystate_n18), .ZN(
        key1FF_keystate_gff_20_SFF_3_n9) );
  DFF_X1 key1FF_keystate_gff_20_SFF_3_Cell_reg ( .D(
        key1FF_keystate_gff_20_SFF_3_n6), .CK(clk), .Q(roundkey1[3]), .QN(
        key1FF_keystate_gff_20_SFF_3_n7) );
  MUX2_X1 key2FF_U10 ( .A(roundkey2[0]), .B(key2[0]), .S(n4), .Z(key2FF_n1) );
  MUX2_X1 key2FF_U9 ( .A(roundkey2[1]), .B(key2[1]), .S(n4), .Z(key2FF_n2) );
  MUX2_X1 key2FF_U8 ( .A(roundkey2[2]), .B(key2[2]), .S(n4), .Z(key2FF_n3) );
  MUX2_X1 key2FF_U7 ( .A(roundkey2[3]), .B(key2[3]), .S(n4), .Z(key2FF_n4) );
  XOR2_X1 key2FF_U6 ( .A(1'b0), .B(key2FF_outputPar[22]), .Z(
        key2FF_counterAdd[4]) );
  XOR2_X1 key2FF_U5 ( .A(1'b0), .B(key2FF_outputPar[21]), .Z(
        key2FF_counterAdd[3]) );
  XOR2_X1 key2FF_U4 ( .A(1'b0), .B(key2FF_outputPar[20]), .Z(
        key2FF_counterAdd[2]) );
  XOR2_X1 key2FF_U3 ( .A(1'b0), .B(key2FF_outputPar[19]), .Z(
        key2FF_counterAdd[1]) );
  XOR2_X1 key2FF_U2 ( .A(1'b0), .B(key2FF_outputPar[18]), .Z(
        key2FF_counterAdd[0]) );
  BUF_X2 key2FF_keystate_U9 ( .A(enKey), .Z(key2FF_keystate_n12) );
  BUF_X1 key2FF_keystate_U8 ( .A(selP), .Z(key2FF_keystate_n17) );
  BUF_X2 key2FF_keystate_U7 ( .A(enKey), .Z(key2FF_keystate_n11) );
  BUF_X1 key2FF_keystate_U6 ( .A(selP), .Z(key2FF_keystate_n16) );
  BUF_X2 key2FF_keystate_U5 ( .A(enKey), .Z(key2FF_keystate_n10) );
  BUF_X1 key2FF_keystate_U4 ( .A(selP), .Z(key2FF_keystate_n15) );
  BUF_X2 key2FF_keystate_U3 ( .A(enKey), .Z(key2FF_keystate_n13) );
  BUF_X1 key2FF_keystate_U2 ( .A(selP), .Z(key2FF_keystate_n14) );
  BUF_X1 key2FF_keystate_U1 ( .A(selP), .Z(key2FF_keystate_n18) );
  OAI21_X1 key2FF_keystate_gff_1_SFF_0_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_1_SFF_0_n8), .A(key2FF_keystate_gff_1_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_1_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_1_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_1_SFF_0_n10), .B2(key2FF_n1), .C1(
        key2FF_keystate_gff_1_SFF_0_n11), .C2(key2FF_outputPar[3]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_1_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_1_SFF_0_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_1_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_1_SFF_0_U2 ( .A(key2FF_keystate_gff_1_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_1_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_1_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_1_SFF_0_n7), .CK(clk), .Q(keyRegKS2[1]), .QN(
        key2FF_keystate_gff_1_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_1_SFF_1_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_1_SFF_1_n8), .A(key2FF_keystate_gff_1_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_1_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_1_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_1_SFF_1_n10), .B2(key2FF_n2), .C1(
        key2FF_keystate_gff_1_SFF_1_n11), .C2(key2FF_outputPar[4]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_1_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_1_SFF_1_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_1_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_1_SFF_1_U2 ( .A(key2FF_keystate_gff_1_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_1_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_1_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_1_SFF_1_n7), .CK(clk), .Q(keyRegKS2[2]), .QN(
        key2FF_keystate_gff_1_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_1_SFF_2_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_1_SFF_2_n8), .A(key2FF_keystate_gff_1_SFF_2_n12), 
        .ZN(key2FF_keystate_gff_1_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_1_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_1_SFF_2_n10), .B2(key2FF_n3), .C1(
        key2FF_keystate_gff_1_SFF_2_n11), .C2(key2FF_outputPar[5]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_1_SFF_2_n12) );
  INV_X1 key2FF_keystate_gff_1_SFF_2_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_1_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_1_SFF_2_U2 ( .A(key2FF_keystate_gff_1_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_1_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_1_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_1_SFF_2_n7), .CK(clk), .Q(keyRegKS2[3]), .QN(
        key2FF_keystate_gff_1_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_1_SFF_3_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_1_SFF_3_n8), .A(key2FF_keystate_gff_1_SFF_3_n12), 
        .ZN(key2FF_keystate_gff_1_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_1_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_1_SFF_3_n10), .B2(key2FF_n4), .C1(
        key2FF_keystate_gff_1_SFF_3_n11), .C2(key2FF_outputPar[6]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_1_SFF_3_n12) );
  INV_X1 key2FF_keystate_gff_1_SFF_3_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_1_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_1_SFF_3_U2 ( .A(key2FF_keystate_gff_1_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_1_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_1_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_1_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[3]), 
        .QN(key2FF_keystate_gff_1_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_2_SFF_0_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_2_SFF_0_n8), .A(key2FF_keystate_gff_2_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_2_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_2_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_2_SFF_0_n10), .B2(keyRegKS2[1]), .C1(
        key2FF_keystate_gff_2_SFF_0_n11), .C2(key2FF_outputPar[7]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_2_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_2_SFF_0_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_2_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_2_SFF_0_U2 ( .A(key2FF_keystate_gff_2_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_2_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_2_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_2_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[4]), 
        .QN(key2FF_keystate_gff_2_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_2_SFF_1_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_2_SFF_1_n8), .A(key2FF_keystate_gff_2_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_2_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_2_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_2_SFF_1_n10), .B2(keyRegKS2[2]), .C1(
        key2FF_keystate_gff_2_SFF_1_n11), .C2(key2FF_outputPar[8]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_2_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_2_SFF_1_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_2_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_2_SFF_1_U2 ( .A(key2FF_keystate_gff_2_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_2_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_2_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_2_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[5]), 
        .QN(key2FF_keystate_gff_2_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_2_SFF_2_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_2_SFF_2_n8), .A(key2FF_keystate_gff_2_SFF_2_n12), 
        .ZN(key2FF_keystate_gff_2_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_2_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_2_SFF_2_n10), .B2(keyRegKS2[3]), .C1(
        key2FF_keystate_gff_2_SFF_2_n11), .C2(key2FF_outputPar[9]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_2_SFF_2_n12) );
  INV_X1 key2FF_keystate_gff_2_SFF_2_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_2_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_2_SFF_2_U2 ( .A(key2FF_keystate_gff_2_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_2_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_2_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_2_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[6]), 
        .QN(key2FF_keystate_gff_2_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_2_SFF_3_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_2_SFF_3_n8), .A(key2FF_keystate_gff_2_SFF_3_n12), 
        .ZN(key2FF_keystate_gff_2_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_2_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_2_SFF_3_n10), .B2(key2FF_outputPar[3]), .C1(
        key2FF_keystate_gff_2_SFF_3_n11), .C2(key2FF_outputPar[10]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_2_SFF_3_n12) );
  INV_X1 key2FF_keystate_gff_2_SFF_3_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_2_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_2_SFF_3_U2 ( .A(key2FF_keystate_gff_2_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_2_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_2_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_2_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[7]), 
        .QN(key2FF_keystate_gff_2_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_3_SFF_0_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_3_SFF_0_n8), .A(key2FF_keystate_gff_3_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_3_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_3_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_3_SFF_0_n10), .B2(key2FF_outputPar[4]), .C1(
        key2FF_keystate_gff_3_SFF_0_n11), .C2(key2FF_outputPar[11]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_3_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_3_SFF_0_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_3_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_3_SFF_0_U2 ( .A(key2FF_keystate_gff_3_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_3_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_3_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_3_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[8]), 
        .QN(key2FF_keystate_gff_3_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_3_SFF_1_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_3_SFF_1_n8), .A(key2FF_keystate_gff_3_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_3_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_3_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_3_SFF_1_n10), .B2(key2FF_outputPar[5]), .C1(
        key2FF_keystate_gff_3_SFF_1_n11), .C2(key2FF_outputPar[12]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_3_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_3_SFF_1_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_3_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_3_SFF_1_U2 ( .A(key2FF_keystate_gff_3_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_3_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_3_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_3_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[9]), 
        .QN(key2FF_keystate_gff_3_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_3_SFF_2_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_3_SFF_2_n7), .A(key2FF_keystate_gff_3_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_3_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_3_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_3_SFF_2_n9), .B2(key2FF_outputPar[6]), .C1(
        key2FF_keystate_gff_3_SFF_2_n10), .C2(key2FF_outputPar[13]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_3_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_3_SFF_2_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_3_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_3_SFF_2_U2 ( .A(key2FF_keystate_gff_3_SFF_2_n10), 
        .ZN(key2FF_keystate_gff_3_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_3_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_3_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[10]), 
        .QN(key2FF_keystate_gff_3_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_3_SFF_3_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_3_SFF_3_n7), .A(key2FF_keystate_gff_3_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_3_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_3_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_3_SFF_3_n9), .B2(key2FF_outputPar[7]), .C1(
        key2FF_keystate_gff_3_SFF_3_n10), .C2(key2FF_outputPar[14]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_3_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_3_SFF_3_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_3_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_3_SFF_3_U2 ( .A(key2FF_keystate_gff_3_SFF_3_n10), 
        .ZN(key2FF_keystate_gff_3_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_3_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_3_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[11]), 
        .QN(key2FF_keystate_gff_3_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_4_SFF_0_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_4_SFF_0_n7), .A(key2FF_keystate_gff_4_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_4_SFF_0_n6) );
  OAI221_X1 key2FF_keystate_gff_4_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_4_SFF_0_n9), .B2(key2FF_outputPar[8]), .C1(
        key2FF_keystate_gff_4_SFF_0_n10), .C2(key2FF_outputPar[15]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_4_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_4_SFF_0_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_4_SFF_0_n10) );
  INV_X1 key2FF_keystate_gff_4_SFF_0_U2 ( .A(key2FF_keystate_gff_4_SFF_0_n10), 
        .ZN(key2FF_keystate_gff_4_SFF_0_n9) );
  DFF_X1 key2FF_keystate_gff_4_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_4_SFF_0_n6), .CK(clk), .Q(key2FF_outputPar[12]), 
        .QN(key2FF_keystate_gff_4_SFF_0_n7) );
  OAI21_X1 key2FF_keystate_gff_4_SFF_1_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_4_SFF_1_n7), .A(key2FF_keystate_gff_4_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_4_SFF_1_n6) );
  OAI221_X1 key2FF_keystate_gff_4_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_4_SFF_1_n9), .B2(key2FF_outputPar[9]), .C1(
        key2FF_keystate_gff_4_SFF_1_n10), .C2(key2FF_outputPar[16]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_4_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_4_SFF_1_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_4_SFF_1_n10) );
  INV_X1 key2FF_keystate_gff_4_SFF_1_U2 ( .A(key2FF_keystate_gff_4_SFF_1_n10), 
        .ZN(key2FF_keystate_gff_4_SFF_1_n9) );
  DFF_X1 key2FF_keystate_gff_4_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_4_SFF_1_n6), .CK(clk), .Q(key2FF_outputPar[13]), 
        .QN(key2FF_keystate_gff_4_SFF_1_n7) );
  OAI21_X1 key2FF_keystate_gff_4_SFF_2_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_4_SFF_2_n7), .A(key2FF_keystate_gff_4_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_4_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_4_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_4_SFF_2_n9), .B2(key2FF_outputPar[10]), .C1(
        key2FF_keystate_gff_4_SFF_2_n10), .C2(key2FF_outputPar[17]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_4_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_4_SFF_2_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_4_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_4_SFF_2_U2 ( .A(key2FF_keystate_gff_4_SFF_2_n10), 
        .ZN(key2FF_keystate_gff_4_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_4_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_4_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[14]), 
        .QN(key2FF_keystate_gff_4_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_4_SFF_3_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_4_SFF_3_n7), .A(key2FF_keystate_gff_4_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_4_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_4_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_4_SFF_3_n9), .B2(key2FF_outputPar[11]), .C1(
        key2FF_keystate_gff_4_SFF_3_n10), .C2(key2FF_counterAdd[0]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_4_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_4_SFF_3_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_4_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_4_SFF_3_U2 ( .A(key2FF_keystate_gff_4_SFF_3_n10), 
        .ZN(key2FF_keystate_gff_4_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_4_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_4_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[15]), 
        .QN(key2FF_keystate_gff_4_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_5_SFF_0_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_5_SFF_0_n8), .A(key2FF_keystate_gff_5_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_5_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_5_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_5_SFF_0_n10), .B2(key2FF_outputPar[12]), .C1(
        key2FF_keystate_gff_5_SFF_0_n11), .C2(key2FF_counterAdd[1]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_5_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_5_SFF_0_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_5_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_5_SFF_0_U2 ( .A(key2FF_keystate_gff_5_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_5_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_5_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_5_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[16]), 
        .QN(key2FF_keystate_gff_5_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_5_SFF_1_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_5_SFF_1_n8), .A(key2FF_keystate_gff_5_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_5_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_5_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_5_SFF_1_n10), .B2(key2FF_outputPar[13]), .C1(
        key2FF_keystate_gff_5_SFF_1_n11), .C2(key2FF_counterAdd[2]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_5_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_5_SFF_1_U3 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_5_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_5_SFF_1_U2 ( .A(key2FF_keystate_gff_5_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_5_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_5_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_5_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[17]), 
        .QN(key2FF_keystate_gff_5_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_5_SFF_2_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_5_SFF_2_n8), .A(key2FF_keystate_gff_5_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_5_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_5_SFF_2_U3 ( .B1(key2FF_keystate_n14), .B2(
        key2FF_outputPar[14]), .C1(key2FF_keystate_gff_5_SFF_2_n10), .C2(
        key2FF_counterAdd[3]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_5_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_5_SFF_2_U2 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_5_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_5_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_5_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[18]), 
        .QN(key2FF_keystate_gff_5_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_5_SFF_3_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_5_SFF_3_n8), .A(key2FF_keystate_gff_5_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_5_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_5_SFF_3_U3 ( .B1(key2FF_keystate_n14), .B2(
        key2FF_outputPar[15]), .C1(key2FF_keystate_gff_5_SFF_3_n10), .C2(
        key2FF_counterAdd[4]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_5_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_5_SFF_3_U2 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_5_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_5_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_5_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[19]), 
        .QN(key2FF_keystate_gff_5_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_6_SFF_0_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_6_SFF_0_n8), .A(key2FF_keystate_gff_6_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_6_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_6_SFF_0_U3 ( .B1(key2FF_keystate_n14), .B2(
        key2FF_outputPar[16]), .C1(key2FF_keystate_gff_6_SFF_0_n10), .C2(
        key2FF_outputPar[23]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_6_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_6_SFF_0_U2 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_6_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_6_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_6_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[20]), 
        .QN(key2FF_keystate_gff_6_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_6_SFF_1_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_6_SFF_1_n8), .A(key2FF_keystate_gff_6_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_6_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_6_SFF_1_U3 ( .B1(key2FF_keystate_n14), .B2(
        key2FF_outputPar[17]), .C1(key2FF_keystate_gff_6_SFF_1_n10), .C2(
        key2FF_outputPar[24]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_6_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_6_SFF_1_U2 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_6_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_6_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_6_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[21]), 
        .QN(key2FF_keystate_gff_6_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_6_SFF_2_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_6_SFF_2_n8), .A(key2FF_keystate_gff_6_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_6_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_6_SFF_2_U3 ( .B1(key2FF_keystate_n14), .B2(
        key2FF_outputPar[18]), .C1(key2FF_keystate_gff_6_SFF_2_n10), .C2(
        key2FF_outputPar[25]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_6_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_6_SFF_2_U2 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_6_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_6_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_6_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[22]), 
        .QN(key2FF_keystate_gff_6_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_6_SFF_3_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_6_SFF_3_n8), .A(key2FF_keystate_gff_6_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_6_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_6_SFF_3_U3 ( .B1(key2FF_keystate_n14), .B2(
        key2FF_outputPar[19]), .C1(key2FF_keystate_gff_6_SFF_3_n10), .C2(
        key2FF_outputPar[26]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_6_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_6_SFF_3_U2 ( .A(key2FF_keystate_n14), .ZN(
        key2FF_keystate_gff_6_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_6_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_6_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[23]), 
        .QN(key2FF_keystate_gff_6_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_7_SFF_0_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_7_SFF_0_n8), .A(key2FF_keystate_gff_7_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_7_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_7_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_7_SFF_0_n10), .B2(key2FF_outputPar[20]), .C1(
        key2FF_keystate_gff_7_SFF_0_n11), .C2(key2FF_outputPar[27]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_7_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_7_SFF_0_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_7_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_7_SFF_0_U2 ( .A(key2FF_keystate_gff_7_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_7_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_7_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_7_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[24]), 
        .QN(key2FF_keystate_gff_7_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_7_SFF_1_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_7_SFF_1_n8), .A(key2FF_keystate_gff_7_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_7_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_7_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_7_SFF_1_n10), .B2(key2FF_outputPar[21]), .C1(
        key2FF_keystate_gff_7_SFF_1_n11), .C2(key2FF_outputPar[28]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_7_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_7_SFF_1_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_7_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_7_SFF_1_U2 ( .A(key2FF_keystate_gff_7_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_7_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_7_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_7_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[25]), 
        .QN(key2FF_keystate_gff_7_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_7_SFF_2_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_7_SFF_2_n7), .A(key2FF_keystate_gff_7_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_7_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_7_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_7_SFF_2_n9), .B2(key2FF_outputPar[22]), .C1(
        key2FF_keystate_gff_7_SFF_2_n10), .C2(key2FF_outputPar[29]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_7_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_7_SFF_2_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_7_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_7_SFF_2_U2 ( .A(key2FF_keystate_gff_7_SFF_2_n10), 
        .ZN(key2FF_keystate_gff_7_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_7_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_7_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[26]), 
        .QN(key2FF_keystate_gff_7_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_7_SFF_3_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_7_SFF_3_n7), .A(key2FF_keystate_gff_7_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_7_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_7_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_7_SFF_3_n9), .B2(key2FF_outputPar[23]), .C1(
        key2FF_keystate_gff_7_SFF_3_n10), .C2(key2FF_outputPar[30]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_7_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_7_SFF_3_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_7_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_7_SFF_3_U2 ( .A(key2FF_keystate_gff_7_SFF_3_n10), 
        .ZN(key2FF_keystate_gff_7_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_7_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_7_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[27]), 
        .QN(key2FF_keystate_gff_7_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_8_SFF_0_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_8_SFF_0_n7), .A(key2FF_keystate_gff_8_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_8_SFF_0_n6) );
  OAI221_X1 key2FF_keystate_gff_8_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_8_SFF_0_n9), .B2(key2FF_outputPar[24]), .C1(
        key2FF_keystate_gff_8_SFF_0_n10), .C2(key2FF_outputPar[31]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_8_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_8_SFF_0_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_8_SFF_0_n10) );
  INV_X1 key2FF_keystate_gff_8_SFF_0_U2 ( .A(key2FF_keystate_gff_8_SFF_0_n10), 
        .ZN(key2FF_keystate_gff_8_SFF_0_n9) );
  DFF_X1 key2FF_keystate_gff_8_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_8_SFF_0_n6), .CK(clk), .Q(key2FF_outputPar[28]), 
        .QN(key2FF_keystate_gff_8_SFF_0_n7) );
  OAI21_X1 key2FF_keystate_gff_8_SFF_1_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_8_SFF_1_n7), .A(key2FF_keystate_gff_8_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_8_SFF_1_n6) );
  OAI221_X1 key2FF_keystate_gff_8_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_8_SFF_1_n9), .B2(key2FF_outputPar[25]), .C1(
        key2FF_keystate_gff_8_SFF_1_n10), .C2(key2FF_outputPar[32]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_8_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_8_SFF_1_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_8_SFF_1_n10) );
  INV_X1 key2FF_keystate_gff_8_SFF_1_U2 ( .A(key2FF_keystate_gff_8_SFF_1_n10), 
        .ZN(key2FF_keystate_gff_8_SFF_1_n9) );
  DFF_X1 key2FF_keystate_gff_8_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_8_SFF_1_n6), .CK(clk), .Q(key2FF_outputPar[29]), 
        .QN(key2FF_keystate_gff_8_SFF_1_n7) );
  OAI21_X1 key2FF_keystate_gff_8_SFF_2_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_8_SFF_2_n7), .A(key2FF_keystate_gff_8_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_8_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_8_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_8_SFF_2_n9), .B2(key2FF_outputPar[26]), .C1(
        key2FF_keystate_gff_8_SFF_2_n10), .C2(key2FF_outputPar[33]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_8_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_8_SFF_2_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_8_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_8_SFF_2_U2 ( .A(key2FF_keystate_gff_8_SFF_2_n10), 
        .ZN(key2FF_keystate_gff_8_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_8_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_8_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[30]), 
        .QN(key2FF_keystate_gff_8_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_8_SFF_3_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_8_SFF_3_n7), .A(key2FF_keystate_gff_8_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_8_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_8_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_8_SFF_3_n9), .B2(key2FF_outputPar[27]), .C1(
        key2FF_keystate_gff_8_SFF_3_n10), .C2(key2FF_outputPar[34]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_8_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_8_SFF_3_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_8_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_8_SFF_3_U2 ( .A(key2FF_keystate_gff_8_SFF_3_n10), 
        .ZN(key2FF_keystate_gff_8_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_8_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_8_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[31]), 
        .QN(key2FF_keystate_gff_8_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_9_SFF_0_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_9_SFF_0_n8), .A(key2FF_keystate_gff_9_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_9_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_9_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_9_SFF_0_n10), .B2(key2FF_outputPar[28]), .C1(
        key2FF_keystate_gff_9_SFF_0_n11), .C2(key2FF_outputPar[35]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_9_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_9_SFF_0_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_9_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_9_SFF_0_U2 ( .A(key2FF_keystate_gff_9_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_9_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_9_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_9_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[32]), 
        .QN(key2FF_keystate_gff_9_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_9_SFF_1_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_9_SFF_1_n8), .A(key2FF_keystate_gff_9_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_9_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_9_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_9_SFF_1_n10), .B2(key2FF_outputPar[29]), .C1(
        key2FF_keystate_gff_9_SFF_1_n11), .C2(key2FF_outputPar[36]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_9_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_9_SFF_1_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_9_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_9_SFF_1_U2 ( .A(key2FF_keystate_gff_9_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_9_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_9_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_9_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[33]), 
        .QN(key2FF_keystate_gff_9_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_9_SFF_2_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_9_SFF_2_n8), .A(key2FF_keystate_gff_9_SFF_2_n12), 
        .ZN(key2FF_keystate_gff_9_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_9_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_9_SFF_2_n10), .B2(key2FF_outputPar[30]), .C1(
        key2FF_keystate_gff_9_SFF_2_n11), .C2(key2FF_outputPar[37]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_9_SFF_2_n12) );
  INV_X1 key2FF_keystate_gff_9_SFF_2_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_9_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_9_SFF_2_U2 ( .A(key2FF_keystate_gff_9_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_9_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_9_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_9_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[34]), 
        .QN(key2FF_keystate_gff_9_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_9_SFF_3_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_9_SFF_3_n8), .A(key2FF_keystate_gff_9_SFF_3_n12), 
        .ZN(key2FF_keystate_gff_9_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_9_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_9_SFF_3_n10), .B2(key2FF_outputPar[31]), .C1(
        key2FF_keystate_gff_9_SFF_3_n11), .C2(key2FF_outputPar[38]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_9_SFF_3_n12) );
  INV_X1 key2FF_keystate_gff_9_SFF_3_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_9_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_9_SFF_3_U2 ( .A(key2FF_keystate_gff_9_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_9_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_9_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_9_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[35]), 
        .QN(key2FF_keystate_gff_9_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_10_SFF_0_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_10_SFF_0_n8), .A(key2FF_keystate_gff_10_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_10_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_10_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_10_SFF_0_n10), .B2(key2FF_outputPar[32]), .C1(
        key2FF_keystate_gff_10_SFF_0_n11), .C2(key2FF_outputPar[39]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_10_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_10_SFF_0_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_10_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_10_SFF_0_U2 ( .A(key2FF_keystate_gff_10_SFF_0_n11), .ZN(key2FF_keystate_gff_10_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_10_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_10_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[36]), 
        .QN(key2FF_keystate_gff_10_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_10_SFF_1_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_10_SFF_1_n8), .A(key2FF_keystate_gff_10_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_10_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_10_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_10_SFF_1_n10), .B2(key2FF_outputPar[33]), .C1(
        key2FF_keystate_gff_10_SFF_1_n11), .C2(key2FF_outputPar[40]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_10_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_10_SFF_1_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_10_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_10_SFF_1_U2 ( .A(key2FF_keystate_gff_10_SFF_1_n11), .ZN(key2FF_keystate_gff_10_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_10_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_10_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[37]), 
        .QN(key2FF_keystate_gff_10_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_10_SFF_2_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_10_SFF_2_n8), .A(key2FF_keystate_gff_10_SFF_2_n12), 
        .ZN(key2FF_keystate_gff_10_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_10_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_10_SFF_2_n10), .B2(key2FF_outputPar[34]), .C1(
        key2FF_keystate_gff_10_SFF_2_n11), .C2(key2FF_outputPar[41]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_10_SFF_2_n12) );
  INV_X1 key2FF_keystate_gff_10_SFF_2_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_10_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_10_SFF_2_U2 ( .A(key2FF_keystate_gff_10_SFF_2_n11), .ZN(key2FF_keystate_gff_10_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_10_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_10_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[38]), 
        .QN(key2FF_keystate_gff_10_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_10_SFF_3_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_10_SFF_3_n8), .A(key2FF_keystate_gff_10_SFF_3_n12), 
        .ZN(key2FF_keystate_gff_10_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_10_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_10_SFF_3_n10), .B2(key2FF_outputPar[35]), .C1(
        key2FF_keystate_gff_10_SFF_3_n11), .C2(key2FF_outputPar[42]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_10_SFF_3_n12) );
  INV_X1 key2FF_keystate_gff_10_SFF_3_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_10_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_10_SFF_3_U2 ( .A(key2FF_keystate_gff_10_SFF_3_n11), .ZN(key2FF_keystate_gff_10_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_10_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_10_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[39]), 
        .QN(key2FF_keystate_gff_10_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_11_SFF_0_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_11_SFF_0_n8), .A(key2FF_keystate_gff_11_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_11_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_11_SFF_0_U3 ( .B1(key2FF_keystate_n17), .B2(
        key2FF_outputPar[36]), .C1(key2FF_keystate_gff_11_SFF_0_n10), .C2(
        key2FF_outputPar[43]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_11_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_11_SFF_0_U2 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_11_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_11_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_11_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[40]), 
        .QN(key2FF_keystate_gff_11_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_11_SFF_1_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_11_SFF_1_n8), .A(key2FF_keystate_gff_11_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_11_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_11_SFF_1_U3 ( .B1(key2FF_keystate_n17), .B2(
        key2FF_outputPar[37]), .C1(key2FF_keystate_gff_11_SFF_1_n10), .C2(
        key2FF_outputPar[44]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_11_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_11_SFF_1_U2 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_11_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_11_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_11_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[41]), 
        .QN(key2FF_keystate_gff_11_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_11_SFF_2_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_11_SFF_2_n7), .A(key2FF_keystate_gff_11_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_11_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_11_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_11_SFF_2_n9), .B2(key2FF_outputPar[38]), .C1(
        key2FF_keystate_gff_11_SFF_2_n10), .C2(key2FF_outputPar[45]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_11_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_11_SFF_2_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_11_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_11_SFF_2_U2 ( .A(key2FF_keystate_gff_11_SFF_2_n10), .ZN(key2FF_keystate_gff_11_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_11_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_11_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[42]), 
        .QN(key2FF_keystate_gff_11_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_11_SFF_3_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_11_SFF_3_n7), .A(key2FF_keystate_gff_11_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_11_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_11_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_11_SFF_3_n9), .B2(key2FF_outputPar[39]), .C1(
        key2FF_keystate_gff_11_SFF_3_n10), .C2(key2FF_outputPar[46]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_11_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_11_SFF_3_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_11_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_11_SFF_3_U2 ( .A(key2FF_keystate_gff_11_SFF_3_n10), .ZN(key2FF_keystate_gff_11_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_11_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_11_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[43]), 
        .QN(key2FF_keystate_gff_11_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_12_SFF_0_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_12_SFF_0_n7), .A(key2FF_keystate_gff_12_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_12_SFF_0_n6) );
  OAI221_X1 key2FF_keystate_gff_12_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_12_SFF_0_n9), .B2(key2FF_outputPar[40]), .C1(
        key2FF_keystate_gff_12_SFF_0_n10), .C2(key2FF_outputPar[47]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_12_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_12_SFF_0_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_12_SFF_0_n10) );
  INV_X1 key2FF_keystate_gff_12_SFF_0_U2 ( .A(key2FF_keystate_gff_12_SFF_0_n10), .ZN(key2FF_keystate_gff_12_SFF_0_n9) );
  DFF_X1 key2FF_keystate_gff_12_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_12_SFF_0_n6), .CK(clk), .Q(key2FF_outputPar[44]), 
        .QN(key2FF_keystate_gff_12_SFF_0_n7) );
  OAI21_X1 key2FF_keystate_gff_12_SFF_1_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_12_SFF_1_n7), .A(key2FF_keystate_gff_12_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_12_SFF_1_n6) );
  OAI221_X1 key2FF_keystate_gff_12_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_12_SFF_1_n9), .B2(key2FF_outputPar[41]), .C1(
        key2FF_keystate_gff_12_SFF_1_n10), .C2(key2FF_outputPar[48]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_12_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_12_SFF_1_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_12_SFF_1_n10) );
  INV_X1 key2FF_keystate_gff_12_SFF_1_U2 ( .A(key2FF_keystate_gff_12_SFF_1_n10), .ZN(key2FF_keystate_gff_12_SFF_1_n9) );
  DFF_X1 key2FF_keystate_gff_12_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_12_SFF_1_n6), .CK(clk), .Q(key2FF_outputPar[45]), 
        .QN(key2FF_keystate_gff_12_SFF_1_n7) );
  OAI21_X1 key2FF_keystate_gff_12_SFF_2_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_12_SFF_2_n7), .A(key2FF_keystate_gff_12_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_12_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_12_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_12_SFF_2_n9), .B2(key2FF_outputPar[42]), .C1(
        key2FF_keystate_gff_12_SFF_2_n10), .C2(key2FF_outputPar[49]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_12_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_12_SFF_2_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_12_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_12_SFF_2_U2 ( .A(key2FF_keystate_gff_12_SFF_2_n10), .ZN(key2FF_keystate_gff_12_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_12_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_12_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[46]), 
        .QN(key2FF_keystate_gff_12_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_12_SFF_3_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_12_SFF_3_n7), .A(key2FF_keystate_gff_12_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_12_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_12_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_12_SFF_3_n9), .B2(key2FF_outputPar[43]), .C1(
        key2FF_keystate_gff_12_SFF_3_n10), .C2(key2FF_outputPar[50]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_12_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_12_SFF_3_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_12_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_12_SFF_3_U2 ( .A(key2FF_keystate_gff_12_SFF_3_n10), .ZN(key2FF_keystate_gff_12_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_12_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_12_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[47]), 
        .QN(key2FF_keystate_gff_12_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_13_SFF_0_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_13_SFF_0_n8), .A(key2FF_keystate_gff_13_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_13_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_13_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_13_SFF_0_n10), .B2(key2FF_outputPar[44]), .C1(
        key2FF_keystate_gff_13_SFF_0_n11), .C2(key2FF_outputPar[51]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_13_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_13_SFF_0_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_13_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_13_SFF_0_U2 ( .A(key2FF_keystate_gff_13_SFF_0_n11), .ZN(key2FF_keystate_gff_13_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_13_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_13_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[48]), 
        .QN(key2FF_keystate_gff_13_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_13_SFF_1_U5 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_13_SFF_1_n8), .A(key2FF_keystate_gff_13_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_13_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_13_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_13_SFF_1_n10), .B2(key2FF_outputPar[45]), .C1(
        key2FF_keystate_gff_13_SFF_1_n11), .C2(key2FF_outputPar[52]), .A(
        key2FF_keystate_n10), .ZN(key2FF_keystate_gff_13_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_13_SFF_1_U3 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_13_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_13_SFF_1_U2 ( .A(key2FF_keystate_gff_13_SFF_1_n11), .ZN(key2FF_keystate_gff_13_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_13_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_13_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[49]), 
        .QN(key2FF_keystate_gff_13_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_13_SFF_2_U4 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_13_SFF_2_n8), .A(key2FF_keystate_gff_13_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_13_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_13_SFF_2_U3 ( .B1(key2FF_keystate_n15), .B2(
        key2FF_outputPar[46]), .C1(key2FF_keystate_gff_13_SFF_2_n10), .C2(
        key2FF_outputPar[53]), .A(key2FF_keystate_n10), .ZN(
        key2FF_keystate_gff_13_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_13_SFF_2_U2 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_13_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_13_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_13_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[50]), 
        .QN(key2FF_keystate_gff_13_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_13_SFF_3_U4 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_13_SFF_3_n8), .A(key2FF_keystate_gff_13_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_13_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_13_SFF_3_U3 ( .B1(key2FF_keystate_n15), .B2(
        key2FF_outputPar[47]), .C1(key2FF_keystate_gff_13_SFF_3_n10), .C2(
        key2FF_outputPar[54]), .A(key2FF_keystate_n10), .ZN(
        key2FF_keystate_gff_13_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_13_SFF_3_U2 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_13_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_13_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_13_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[51]), 
        .QN(key2FF_keystate_gff_13_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_14_SFF_0_U4 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_14_SFF_0_n8), .A(key2FF_keystate_gff_14_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_14_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_14_SFF_0_U3 ( .B1(key2FF_keystate_n15), .B2(
        key2FF_outputPar[48]), .C1(key2FF_keystate_gff_14_SFF_0_n10), .C2(
        key2FF_outputPar[55]), .A(key2FF_keystate_n10), .ZN(
        key2FF_keystate_gff_14_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_14_SFF_0_U2 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_14_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_14_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_14_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[52]), 
        .QN(key2FF_keystate_gff_14_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_14_SFF_1_U4 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_14_SFF_1_n8), .A(key2FF_keystate_gff_14_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_14_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_14_SFF_1_U3 ( .B1(key2FF_keystate_n15), .B2(
        key2FF_outputPar[49]), .C1(key2FF_keystate_gff_14_SFF_1_n10), .C2(
        key2FF_outputPar[56]), .A(key2FF_keystate_n10), .ZN(
        key2FF_keystate_gff_14_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_14_SFF_1_U2 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_14_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_14_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_14_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[53]), 
        .QN(key2FF_keystate_gff_14_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_14_SFF_2_U4 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_14_SFF_2_n8), .A(key2FF_keystate_gff_14_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_14_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_14_SFF_2_U3 ( .B1(key2FF_keystate_n15), .B2(
        key2FF_outputPar[50]), .C1(key2FF_keystate_gff_14_SFF_2_n10), .C2(
        key2FF_outputPar[57]), .A(key2FF_keystate_n10), .ZN(
        key2FF_keystate_gff_14_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_14_SFF_2_U2 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_14_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_14_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_14_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[54]), 
        .QN(key2FF_keystate_gff_14_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_14_SFF_3_U4 ( .B1(key2FF_keystate_n10), .B2(
        key2FF_keystate_gff_14_SFF_3_n8), .A(key2FF_keystate_gff_14_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_14_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_14_SFF_3_U3 ( .B1(key2FF_keystate_n15), .B2(
        key2FF_outputPar[51]), .C1(key2FF_keystate_gff_14_SFF_3_n10), .C2(
        key2FF_outputPar[58]), .A(key2FF_keystate_n10), .ZN(
        key2FF_keystate_gff_14_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_14_SFF_3_U2 ( .A(key2FF_keystate_n15), .ZN(
        key2FF_keystate_gff_14_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_14_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_14_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[55]), 
        .QN(key2FF_keystate_gff_14_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_15_SFF_0_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_15_SFF_0_n8), .A(key2FF_keystate_gff_15_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_15_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_15_SFF_0_U3 ( .B1(key2FF_keystate_n17), .B2(
        key2FF_outputPar[52]), .C1(key2FF_keystate_gff_15_SFF_0_n10), .C2(
        key2FF_outputPar[59]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_15_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_15_SFF_0_U2 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_15_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_15_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_15_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[56]), 
        .QN(key2FF_keystate_gff_15_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_15_SFF_1_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_15_SFF_1_n8), .A(key2FF_keystate_gff_15_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_15_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_15_SFF_1_U3 ( .B1(key2FF_keystate_n17), .B2(
        key2FF_outputPar[53]), .C1(key2FF_keystate_gff_15_SFF_1_n10), .C2(
        key2FF_outputPar[60]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_15_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_15_SFF_1_U2 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_15_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_15_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_15_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[57]), 
        .QN(key2FF_keystate_gff_15_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_15_SFF_2_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_15_SFF_2_n7), .A(key2FF_keystate_gff_15_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_15_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_15_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_15_SFF_2_n9), .B2(key2FF_outputPar[54]), .C1(
        key2FF_keystate_gff_15_SFF_2_n10), .C2(key2FF_outputPar[61]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_15_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_15_SFF_2_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_15_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_15_SFF_2_U2 ( .A(key2FF_keystate_gff_15_SFF_2_n10), .ZN(key2FF_keystate_gff_15_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_15_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_15_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[58]), 
        .QN(key2FF_keystate_gff_15_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_15_SFF_3_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_15_SFF_3_n7), .A(key2FF_keystate_gff_15_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_15_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_15_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_15_SFF_3_n9), .B2(key2FF_outputPar[55]), .C1(
        key2FF_keystate_gff_15_SFF_3_n10), .C2(key2FF_outputPar[62]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_15_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_15_SFF_3_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_15_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_15_SFF_3_U2 ( .A(key2FF_keystate_gff_15_SFF_3_n10), .ZN(key2FF_keystate_gff_15_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_15_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_15_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[59]), 
        .QN(key2FF_keystate_gff_15_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_16_SFF_0_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_16_SFF_0_n7), .A(key2FF_keystate_gff_16_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_16_SFF_0_n6) );
  OAI221_X1 key2FF_keystate_gff_16_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_16_SFF_0_n9), .B2(key2FF_outputPar[56]), .C1(
        key2FF_keystate_gff_16_SFF_0_n10), .C2(key2FF_outputPar[63]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_16_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_16_SFF_0_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_16_SFF_0_n10) );
  INV_X1 key2FF_keystate_gff_16_SFF_0_U2 ( .A(key2FF_keystate_gff_16_SFF_0_n10), .ZN(key2FF_keystate_gff_16_SFF_0_n9) );
  DFF_X1 key2FF_keystate_gff_16_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_16_SFF_0_n6), .CK(clk), .Q(key2FF_outputPar[60]), 
        .QN(key2FF_keystate_gff_16_SFF_0_n7) );
  OAI21_X1 key2FF_keystate_gff_16_SFF_1_U5 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_16_SFF_1_n7), .A(key2FF_keystate_gff_16_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_16_SFF_1_n6) );
  OAI221_X1 key2FF_keystate_gff_16_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_16_SFF_1_n9), .B2(key2FF_outputPar[57]), .C1(
        key2FF_keystate_gff_16_SFF_1_n10), .C2(key2FF_outputPar[64]), .A(
        key2FF_keystate_n13), .ZN(key2FF_keystate_gff_16_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_16_SFF_1_U3 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_16_SFF_1_n10) );
  INV_X1 key2FF_keystate_gff_16_SFF_1_U2 ( .A(key2FF_keystate_gff_16_SFF_1_n10), .ZN(key2FF_keystate_gff_16_SFF_1_n9) );
  DFF_X1 key2FF_keystate_gff_16_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_16_SFF_1_n6), .CK(clk), .Q(key2FF_outputPar[61]), 
        .QN(key2FF_keystate_gff_16_SFF_1_n7) );
  OAI21_X1 key2FF_keystate_gff_16_SFF_2_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_16_SFF_2_n7), .A(key2FF_keystate_gff_16_SFF_2_n10), 
        .ZN(key2FF_keystate_gff_16_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_16_SFF_2_U3 ( .B1(key2FF_keystate_n18), .B2(
        key2FF_outputPar[58]), .C1(key2FF_keystate_gff_16_SFF_2_n9), .C2(
        key2FF_outputPar[65]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_16_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_16_SFF_2_U2 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_16_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_16_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_16_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[62]), 
        .QN(key2FF_keystate_gff_16_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_16_SFF_3_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_16_SFF_3_n7), .A(key2FF_keystate_gff_16_SFF_3_n10), 
        .ZN(key2FF_keystate_gff_16_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_16_SFF_3_U3 ( .B1(key2FF_keystate_n18), .B2(
        key2FF_outputPar[59]), .C1(key2FF_keystate_gff_16_SFF_3_n9), .C2(
        key2FF_outputPar[66]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_16_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_16_SFF_3_U2 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_16_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_16_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_16_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[63]), 
        .QN(key2FF_keystate_gff_16_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_17_SFF_0_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_17_SFF_0_n8), .A(key2FF_keystate_gff_17_SFF_0_n12), 
        .ZN(key2FF_keystate_gff_17_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_17_SFF_0_U4 ( .B1(
        key2FF_keystate_gff_17_SFF_0_n10), .B2(key2FF_outputPar[60]), .C1(
        key2FF_keystate_gff_17_SFF_0_n11), .C2(key2FF_outputPar[67]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_17_SFF_0_n12) );
  INV_X1 key2FF_keystate_gff_17_SFF_0_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_17_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_17_SFF_0_U2 ( .A(key2FF_keystate_gff_17_SFF_0_n11), .ZN(key2FF_keystate_gff_17_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_17_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_17_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[64]), 
        .QN(key2FF_keystate_gff_17_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_17_SFF_1_U5 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_17_SFF_1_n8), .A(key2FF_keystate_gff_17_SFF_1_n12), 
        .ZN(key2FF_keystate_gff_17_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_17_SFF_1_U4 ( .B1(
        key2FF_keystate_gff_17_SFF_1_n10), .B2(key2FF_outputPar[61]), .C1(
        key2FF_keystate_gff_17_SFF_1_n11), .C2(key2FF_outputPar[68]), .A(
        key2FF_keystate_n11), .ZN(key2FF_keystate_gff_17_SFF_1_n12) );
  INV_X1 key2FF_keystate_gff_17_SFF_1_U3 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_17_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_17_SFF_1_U2 ( .A(key2FF_keystate_gff_17_SFF_1_n11), .ZN(key2FF_keystate_gff_17_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_17_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_17_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[65]), 
        .QN(key2FF_keystate_gff_17_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_17_SFF_2_U4 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_17_SFF_2_n8), .A(key2FF_keystate_gff_17_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_17_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_17_SFF_2_U3 ( .B1(key2FF_keystate_n16), .B2(
        key2FF_outputPar[62]), .C1(key2FF_keystate_gff_17_SFF_2_n10), .C2(
        key2FF_outputPar[69]), .A(key2FF_keystate_n11), .ZN(
        key2FF_keystate_gff_17_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_17_SFF_2_U2 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_17_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_17_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_17_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[66]), 
        .QN(key2FF_keystate_gff_17_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_17_SFF_3_U4 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_17_SFF_3_n8), .A(key2FF_keystate_gff_17_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_17_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_17_SFF_3_U3 ( .B1(key2FF_keystate_n16), .B2(
        key2FF_outputPar[63]), .C1(key2FF_keystate_gff_17_SFF_3_n10), .C2(
        key2FF_outputPar[70]), .A(key2FF_keystate_n11), .ZN(
        key2FF_keystate_gff_17_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_17_SFF_3_U2 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_17_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_17_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_17_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[67]), 
        .QN(key2FF_keystate_gff_17_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_18_SFF_0_U4 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_18_SFF_0_n8), .A(key2FF_keystate_gff_18_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_18_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_18_SFF_0_U3 ( .B1(key2FF_keystate_n16), .B2(
        key2FF_outputPar[64]), .C1(key2FF_keystate_gff_18_SFF_0_n10), .C2(
        key2FF_outputPar[71]), .A(key2FF_keystate_n11), .ZN(
        key2FF_keystate_gff_18_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_18_SFF_0_U2 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_18_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_18_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_18_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[68]), 
        .QN(key2FF_keystate_gff_18_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_18_SFF_1_U4 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_18_SFF_1_n8), .A(key2FF_keystate_gff_18_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_18_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_18_SFF_1_U3 ( .B1(key2FF_keystate_n16), .B2(
        key2FF_outputPar[65]), .C1(key2FF_keystate_gff_18_SFF_1_n10), .C2(
        key2FF_outputPar[72]), .A(key2FF_keystate_n11), .ZN(
        key2FF_keystate_gff_18_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_18_SFF_1_U2 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_18_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_18_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_18_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[69]), 
        .QN(key2FF_keystate_gff_18_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_18_SFF_2_U4 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_18_SFF_2_n8), .A(key2FF_keystate_gff_18_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_18_SFF_2_n7) );
  OAI221_X1 key2FF_keystate_gff_18_SFF_2_U3 ( .B1(key2FF_keystate_n16), .B2(
        key2FF_outputPar[66]), .C1(key2FF_keystate_gff_18_SFF_2_n10), .C2(
        key2FF_outputPar[73]), .A(key2FF_keystate_n11), .ZN(
        key2FF_keystate_gff_18_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_18_SFF_2_U2 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_18_SFF_2_n10) );
  DFF_X1 key2FF_keystate_gff_18_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_18_SFF_2_n7), .CK(clk), .Q(key2FF_outputPar[70]), 
        .QN(key2FF_keystate_gff_18_SFF_2_n8) );
  OAI21_X1 key2FF_keystate_gff_18_SFF_3_U4 ( .B1(key2FF_keystate_n11), .B2(
        key2FF_keystate_gff_18_SFF_3_n8), .A(key2FF_keystate_gff_18_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_18_SFF_3_n7) );
  OAI221_X1 key2FF_keystate_gff_18_SFF_3_U3 ( .B1(key2FF_keystate_n16), .B2(
        key2FF_outputPar[67]), .C1(key2FF_keystate_gff_18_SFF_3_n10), .C2(
        key2FF_outputPar[74]), .A(key2FF_keystate_n11), .ZN(
        key2FF_keystate_gff_18_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_18_SFF_3_U2 ( .A(key2FF_keystate_n16), .ZN(
        key2FF_keystate_gff_18_SFF_3_n10) );
  DFF_X1 key2FF_keystate_gff_18_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_18_SFF_3_n7), .CK(clk), .Q(key2FF_outputPar[71]), 
        .QN(key2FF_keystate_gff_18_SFF_3_n8) );
  OAI21_X1 key2FF_keystate_gff_19_SFF_0_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_19_SFF_0_n8), .A(key2FF_keystate_gff_19_SFF_0_n11), 
        .ZN(key2FF_keystate_gff_19_SFF_0_n7) );
  OAI221_X1 key2FF_keystate_gff_19_SFF_0_U3 ( .B1(key2FF_keystate_n17), .B2(
        key2FF_outputPar[68]), .C1(key2FF_keystate_gff_19_SFF_0_n10), .C2(
        key2FF_outputPar[75]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_19_SFF_0_n11) );
  INV_X1 key2FF_keystate_gff_19_SFF_0_U2 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_19_SFF_0_n10) );
  DFF_X1 key2FF_keystate_gff_19_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_19_SFF_0_n7), .CK(clk), .Q(key2FF_outputPar[72]), 
        .QN(key2FF_keystate_gff_19_SFF_0_n8) );
  OAI21_X1 key2FF_keystate_gff_19_SFF_1_U4 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_19_SFF_1_n8), .A(key2FF_keystate_gff_19_SFF_1_n11), 
        .ZN(key2FF_keystate_gff_19_SFF_1_n7) );
  OAI221_X1 key2FF_keystate_gff_19_SFF_1_U3 ( .B1(key2FF_keystate_n17), .B2(
        key2FF_outputPar[69]), .C1(key2FF_keystate_gff_19_SFF_1_n10), .C2(
        roundkey2[0]), .A(key2FF_keystate_n12), .ZN(
        key2FF_keystate_gff_19_SFF_1_n11) );
  INV_X1 key2FF_keystate_gff_19_SFF_1_U2 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_19_SFF_1_n10) );
  DFF_X1 key2FF_keystate_gff_19_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_19_SFF_1_n7), .CK(clk), .Q(key2FF_outputPar[73]), 
        .QN(key2FF_keystate_gff_19_SFF_1_n8) );
  OAI21_X1 key2FF_keystate_gff_19_SFF_2_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_19_SFF_2_n7), .A(key2FF_keystate_gff_19_SFF_2_n11), 
        .ZN(key2FF_keystate_gff_19_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_19_SFF_2_U4 ( .B1(
        key2FF_keystate_gff_19_SFF_2_n9), .B2(key2FF_outputPar[70]), .C1(
        key2FF_keystate_gff_19_SFF_2_n10), .C2(roundkey2[1]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_19_SFF_2_n11) );
  INV_X1 key2FF_keystate_gff_19_SFF_2_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_19_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_19_SFF_2_U2 ( .A(key2FF_keystate_gff_19_SFF_2_n10), .ZN(key2FF_keystate_gff_19_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_19_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_19_SFF_2_n6), .CK(clk), .Q(key2FF_outputPar[74]), 
        .QN(key2FF_keystate_gff_19_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_19_SFF_3_U5 ( .B1(key2FF_keystate_n12), .B2(
        key2FF_keystate_gff_19_SFF_3_n7), .A(key2FF_keystate_gff_19_SFF_3_n11), 
        .ZN(key2FF_keystate_gff_19_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_19_SFF_3_U4 ( .B1(
        key2FF_keystate_gff_19_SFF_3_n9), .B2(key2FF_outputPar[71]), .C1(
        key2FF_keystate_gff_19_SFF_3_n10), .C2(roundkey2[2]), .A(
        key2FF_keystate_n12), .ZN(key2FF_keystate_gff_19_SFF_3_n11) );
  INV_X1 key2FF_keystate_gff_19_SFF_3_U3 ( .A(key2FF_keystate_n17), .ZN(
        key2FF_keystate_gff_19_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_19_SFF_3_U2 ( .A(key2FF_keystate_gff_19_SFF_3_n10), .ZN(key2FF_keystate_gff_19_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_19_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_19_SFF_3_n6), .CK(clk), .Q(key2FF_outputPar[75]), 
        .QN(key2FF_keystate_gff_19_SFF_3_n7) );
  OAI21_X1 key2FF_keystate_gff_20_SFF_0_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_20_SFF_0_n7), .A(key2FF_keystate_gff_20_SFF_0_n10), 
        .ZN(key2FF_keystate_gff_20_SFF_0_n6) );
  OAI221_X1 key2FF_keystate_gff_20_SFF_0_U3 ( .B1(key2FF_keystate_n18), .B2(
        key2FF_outputPar[72]), .C1(key2FF_keystate_gff_20_SFF_0_n9), .C2(
        sboxOut2[0]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_20_SFF_0_n10) );
  INV_X1 key2FF_keystate_gff_20_SFF_0_U2 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_20_SFF_0_n9) );
  DFF_X1 key2FF_keystate_gff_20_SFF_0_Cell_reg ( .D(
        key2FF_keystate_gff_20_SFF_0_n6), .CK(clk), .Q(roundkey2[0]), .QN(
        key2FF_keystate_gff_20_SFF_0_n7) );
  OAI21_X1 key2FF_keystate_gff_20_SFF_1_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_20_SFF_1_n7), .A(key2FF_keystate_gff_20_SFF_1_n10), 
        .ZN(key2FF_keystate_gff_20_SFF_1_n6) );
  OAI221_X1 key2FF_keystate_gff_20_SFF_1_U3 ( .B1(key2FF_keystate_n18), .B2(
        key2FF_outputPar[73]), .C1(key2FF_keystate_gff_20_SFF_1_n9), .C2(
        sboxOut2[1]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_20_SFF_1_n10) );
  INV_X1 key2FF_keystate_gff_20_SFF_1_U2 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_20_SFF_1_n9) );
  DFF_X1 key2FF_keystate_gff_20_SFF_1_Cell_reg ( .D(
        key2FF_keystate_gff_20_SFF_1_n6), .CK(clk), .Q(roundkey2[1]), .QN(
        key2FF_keystate_gff_20_SFF_1_n7) );
  OAI21_X1 key2FF_keystate_gff_20_SFF_2_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_20_SFF_2_n7), .A(key2FF_keystate_gff_20_SFF_2_n10), 
        .ZN(key2FF_keystate_gff_20_SFF_2_n6) );
  OAI221_X1 key2FF_keystate_gff_20_SFF_2_U3 ( .B1(key2FF_keystate_n18), .B2(
        key2FF_outputPar[74]), .C1(key2FF_keystate_gff_20_SFF_2_n9), .C2(
        sboxOut2[2]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_20_SFF_2_n10) );
  INV_X1 key2FF_keystate_gff_20_SFF_2_U2 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_20_SFF_2_n9) );
  DFF_X1 key2FF_keystate_gff_20_SFF_2_Cell_reg ( .D(
        key2FF_keystate_gff_20_SFF_2_n6), .CK(clk), .Q(roundkey2[2]), .QN(
        key2FF_keystate_gff_20_SFF_2_n7) );
  OAI21_X1 key2FF_keystate_gff_20_SFF_3_U4 ( .B1(key2FF_keystate_n13), .B2(
        key2FF_keystate_gff_20_SFF_3_n7), .A(key2FF_keystate_gff_20_SFF_3_n10), 
        .ZN(key2FF_keystate_gff_20_SFF_3_n6) );
  OAI221_X1 key2FF_keystate_gff_20_SFF_3_U3 ( .B1(key2FF_keystate_n18), .B2(
        key2FF_outputPar[75]), .C1(key2FF_keystate_gff_20_SFF_3_n9), .C2(
        sboxOut2[3]), .A(key2FF_keystate_n13), .ZN(
        key2FF_keystate_gff_20_SFF_3_n10) );
  INV_X1 key2FF_keystate_gff_20_SFF_3_U2 ( .A(key2FF_keystate_n18), .ZN(
        key2FF_keystate_gff_20_SFF_3_n9) );
  DFF_X1 key2FF_keystate_gff_20_SFF_3_Cell_reg ( .D(
        key2FF_keystate_gff_20_SFF_3_n6), .CK(clk), .Q(roundkey2[3]), .QN(
        key2FF_keystate_gff_20_SFF_3_n7) );
  MUX2_X1 key3FF_U10 ( .A(roundkey3[0]), .B(key3[0]), .S(n4), .Z(key3FF_n1) );
  MUX2_X1 key3FF_U9 ( .A(roundkey3[1]), .B(key3[1]), .S(n4), .Z(key3FF_n2) );
  MUX2_X1 key3FF_U8 ( .A(roundkey3[2]), .B(key3[2]), .S(n4), .Z(key3FF_n3) );
  MUX2_X1 key3FF_U7 ( .A(roundkey3[3]), .B(key3[3]), .S(n4), .Z(key3FF_n4) );
  XOR2_X1 key3FF_U6 ( .A(1'b0), .B(key3FF_outputPar[22]), .Z(
        key3FF_counterAdd[4]) );
  XOR2_X1 key3FF_U5 ( .A(1'b0), .B(key3FF_outputPar[21]), .Z(
        key3FF_counterAdd[3]) );
  XOR2_X1 key3FF_U4 ( .A(1'b0), .B(key3FF_outputPar[20]), .Z(
        key3FF_counterAdd[2]) );
  XOR2_X1 key3FF_U3 ( .A(1'b0), .B(key3FF_outputPar[19]), .Z(
        key3FF_counterAdd[1]) );
  XOR2_X1 key3FF_U2 ( .A(1'b0), .B(key3FF_outputPar[18]), .Z(
        key3FF_counterAdd[0]) );
  BUF_X2 key3FF_keystate_U9 ( .A(enKey), .Z(key3FF_keystate_n10) );
  BUF_X1 key3FF_keystate_U8 ( .A(selP), .Z(key3FF_keystate_n15) );
  BUF_X2 key3FF_keystate_U7 ( .A(enKey), .Z(key3FF_keystate_n11) );
  BUF_X1 key3FF_keystate_U6 ( .A(selP), .Z(key3FF_keystate_n16) );
  BUF_X2 key3FF_keystate_U5 ( .A(enKey), .Z(key3FF_keystate_n12) );
  BUF_X1 key3FF_keystate_U4 ( .A(selP), .Z(key3FF_keystate_n14) );
  BUF_X2 key3FF_keystate_U3 ( .A(enKey), .Z(key3FF_keystate_n13) );
  BUF_X1 key3FF_keystate_U2 ( .A(selP), .Z(key3FF_keystate_n18) );
  BUF_X1 key3FF_keystate_U1 ( .A(selP), .Z(key3FF_keystate_n17) );
  OAI21_X1 key3FF_keystate_gff_1_SFF_0_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_1_SFF_0_n8), .A(key3FF_keystate_gff_1_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_1_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_1_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_1_SFF_0_n10), .B2(key3FF_n1), .C1(
        key3FF_keystate_gff_1_SFF_0_n11), .C2(key3FF_outputPar[3]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_1_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_1_SFF_0_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_1_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_1_SFF_0_U2 ( .A(key3FF_keystate_gff_1_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_1_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_1_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_1_SFF_0_n7), .CK(clk), .Q(keyRegKS3[1]), .QN(
        key3FF_keystate_gff_1_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_1_SFF_1_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_1_SFF_1_n8), .A(key3FF_keystate_gff_1_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_1_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_1_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_1_SFF_1_n10), .B2(key3FF_n2), .C1(
        key3FF_keystate_gff_1_SFF_1_n11), .C2(key3FF_outputPar[4]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_1_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_1_SFF_1_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_1_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_1_SFF_1_U2 ( .A(key3FF_keystate_gff_1_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_1_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_1_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_1_SFF_1_n7), .CK(clk), .Q(keyRegKS3[2]), .QN(
        key3FF_keystate_gff_1_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_1_SFF_2_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_1_SFF_2_n8), .A(key3FF_keystate_gff_1_SFF_2_n12), 
        .ZN(key3FF_keystate_gff_1_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_1_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_1_SFF_2_n10), .B2(key3FF_n3), .C1(
        key3FF_keystate_gff_1_SFF_2_n11), .C2(key3FF_outputPar[5]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_1_SFF_2_n12) );
  INV_X1 key3FF_keystate_gff_1_SFF_2_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_1_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_1_SFF_2_U2 ( .A(key3FF_keystate_gff_1_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_1_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_1_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_1_SFF_2_n7), .CK(clk), .Q(keyRegKS3[3]), .QN(
        key3FF_keystate_gff_1_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_1_SFF_3_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_1_SFF_3_n8), .A(key3FF_keystate_gff_1_SFF_3_n12), 
        .ZN(key3FF_keystate_gff_1_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_1_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_1_SFF_3_n10), .B2(key3FF_n4), .C1(
        key3FF_keystate_gff_1_SFF_3_n11), .C2(key3FF_outputPar[6]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_1_SFF_3_n12) );
  INV_X1 key3FF_keystate_gff_1_SFF_3_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_1_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_1_SFF_3_U2 ( .A(key3FF_keystate_gff_1_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_1_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_1_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_1_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[3]), 
        .QN(key3FF_keystate_gff_1_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_2_SFF_0_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_2_SFF_0_n8), .A(key3FF_keystate_gff_2_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_2_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_2_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_2_SFF_0_n10), .B2(keyRegKS3[1]), .C1(
        key3FF_keystate_gff_2_SFF_0_n11), .C2(key3FF_outputPar[7]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_2_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_2_SFF_0_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_2_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_2_SFF_0_U2 ( .A(key3FF_keystate_gff_2_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_2_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_2_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_2_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[4]), 
        .QN(key3FF_keystate_gff_2_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_2_SFF_1_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_2_SFF_1_n8), .A(key3FF_keystate_gff_2_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_2_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_2_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_2_SFF_1_n10), .B2(keyRegKS3[2]), .C1(
        key3FF_keystate_gff_2_SFF_1_n11), .C2(key3FF_outputPar[8]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_2_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_2_SFF_1_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_2_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_2_SFF_1_U2 ( .A(key3FF_keystate_gff_2_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_2_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_2_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_2_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[5]), 
        .QN(key3FF_keystate_gff_2_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_2_SFF_2_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_2_SFF_2_n8), .A(key3FF_keystate_gff_2_SFF_2_n12), 
        .ZN(key3FF_keystate_gff_2_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_2_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_2_SFF_2_n10), .B2(keyRegKS3[3]), .C1(
        key3FF_keystate_gff_2_SFF_2_n11), .C2(key3FF_outputPar[9]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_2_SFF_2_n12) );
  INV_X1 key3FF_keystate_gff_2_SFF_2_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_2_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_2_SFF_2_U2 ( .A(key3FF_keystate_gff_2_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_2_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_2_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_2_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[6]), 
        .QN(key3FF_keystate_gff_2_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_2_SFF_3_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_2_SFF_3_n8), .A(key3FF_keystate_gff_2_SFF_3_n12), 
        .ZN(key3FF_keystate_gff_2_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_2_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_2_SFF_3_n10), .B2(key3FF_outputPar[3]), .C1(
        key3FF_keystate_gff_2_SFF_3_n11), .C2(key3FF_outputPar[10]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_2_SFF_3_n12) );
  INV_X1 key3FF_keystate_gff_2_SFF_3_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_2_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_2_SFF_3_U2 ( .A(key3FF_keystate_gff_2_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_2_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_2_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_2_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[7]), 
        .QN(key3FF_keystate_gff_2_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_3_SFF_0_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_3_SFF_0_n8), .A(key3FF_keystate_gff_3_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_3_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_3_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_3_SFF_0_n10), .B2(key3FF_outputPar[4]), .C1(
        key3FF_keystate_gff_3_SFF_0_n11), .C2(key3FF_outputPar[11]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_3_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_3_SFF_0_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_3_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_3_SFF_0_U2 ( .A(key3FF_keystate_gff_3_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_3_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_3_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_3_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[8]), 
        .QN(key3FF_keystate_gff_3_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_3_SFF_1_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_3_SFF_1_n8), .A(key3FF_keystate_gff_3_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_3_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_3_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_3_SFF_1_n10), .B2(key3FF_outputPar[5]), .C1(
        key3FF_keystate_gff_3_SFF_1_n11), .C2(key3FF_outputPar[12]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_3_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_3_SFF_1_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_3_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_3_SFF_1_U2 ( .A(key3FF_keystate_gff_3_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_3_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_3_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_3_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[9]), 
        .QN(key3FF_keystate_gff_3_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_3_SFF_2_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_3_SFF_2_n7), .A(key3FF_keystate_gff_3_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_3_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_3_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_3_SFF_2_n9), .B2(key3FF_outputPar[6]), .C1(
        key3FF_keystate_gff_3_SFF_2_n10), .C2(key3FF_outputPar[13]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_3_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_3_SFF_2_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_3_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_3_SFF_2_U2 ( .A(key3FF_keystate_gff_3_SFF_2_n10), 
        .ZN(key3FF_keystate_gff_3_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_3_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_3_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[10]), 
        .QN(key3FF_keystate_gff_3_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_3_SFF_3_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_3_SFF_3_n7), .A(key3FF_keystate_gff_3_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_3_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_3_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_3_SFF_3_n9), .B2(key3FF_outputPar[7]), .C1(
        key3FF_keystate_gff_3_SFF_3_n10), .C2(key3FF_outputPar[14]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_3_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_3_SFF_3_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_3_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_3_SFF_3_U2 ( .A(key3FF_keystate_gff_3_SFF_3_n10), 
        .ZN(key3FF_keystate_gff_3_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_3_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_3_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[11]), 
        .QN(key3FF_keystate_gff_3_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_4_SFF_0_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_4_SFF_0_n7), .A(key3FF_keystate_gff_4_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_4_SFF_0_n6) );
  OAI221_X1 key3FF_keystate_gff_4_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_4_SFF_0_n9), .B2(key3FF_outputPar[8]), .C1(
        key3FF_keystate_gff_4_SFF_0_n10), .C2(key3FF_outputPar[15]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_4_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_4_SFF_0_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_4_SFF_0_n10) );
  INV_X1 key3FF_keystate_gff_4_SFF_0_U2 ( .A(key3FF_keystate_gff_4_SFF_0_n10), 
        .ZN(key3FF_keystate_gff_4_SFF_0_n9) );
  DFF_X1 key3FF_keystate_gff_4_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_4_SFF_0_n6), .CK(clk), .Q(key3FF_outputPar[12]), 
        .QN(key3FF_keystate_gff_4_SFF_0_n7) );
  OAI21_X1 key3FF_keystate_gff_4_SFF_1_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_4_SFF_1_n7), .A(key3FF_keystate_gff_4_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_4_SFF_1_n6) );
  OAI221_X1 key3FF_keystate_gff_4_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_4_SFF_1_n9), .B2(key3FF_outputPar[9]), .C1(
        key3FF_keystate_gff_4_SFF_1_n10), .C2(key3FF_outputPar[16]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_4_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_4_SFF_1_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_4_SFF_1_n10) );
  INV_X1 key3FF_keystate_gff_4_SFF_1_U2 ( .A(key3FF_keystate_gff_4_SFF_1_n10), 
        .ZN(key3FF_keystate_gff_4_SFF_1_n9) );
  DFF_X1 key3FF_keystate_gff_4_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_4_SFF_1_n6), .CK(clk), .Q(key3FF_outputPar[13]), 
        .QN(key3FF_keystate_gff_4_SFF_1_n7) );
  OAI21_X1 key3FF_keystate_gff_4_SFF_2_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_4_SFF_2_n7), .A(key3FF_keystate_gff_4_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_4_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_4_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_4_SFF_2_n9), .B2(key3FF_outputPar[10]), .C1(
        key3FF_keystate_gff_4_SFF_2_n10), .C2(key3FF_outputPar[17]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_4_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_4_SFF_2_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_4_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_4_SFF_2_U2 ( .A(key3FF_keystate_gff_4_SFF_2_n10), 
        .ZN(key3FF_keystate_gff_4_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_4_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_4_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[14]), 
        .QN(key3FF_keystate_gff_4_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_4_SFF_3_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_4_SFF_3_n7), .A(key3FF_keystate_gff_4_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_4_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_4_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_4_SFF_3_n9), .B2(key3FF_outputPar[11]), .C1(
        key3FF_keystate_gff_4_SFF_3_n10), .C2(key3FF_counterAdd[0]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_4_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_4_SFF_3_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_4_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_4_SFF_3_U2 ( .A(key3FF_keystate_gff_4_SFF_3_n10), 
        .ZN(key3FF_keystate_gff_4_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_4_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_4_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[15]), 
        .QN(key3FF_keystate_gff_4_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_5_SFF_0_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_5_SFF_0_n8), .A(key3FF_keystate_gff_5_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_5_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_5_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_5_SFF_0_n10), .B2(key3FF_outputPar[12]), .C1(
        key3FF_keystate_gff_5_SFF_0_n11), .C2(key3FF_counterAdd[1]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_5_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_5_SFF_0_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_5_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_5_SFF_0_U2 ( .A(key3FF_keystate_gff_5_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_5_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_5_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_5_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[16]), 
        .QN(key3FF_keystate_gff_5_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_5_SFF_1_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_5_SFF_1_n8), .A(key3FF_keystate_gff_5_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_5_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_5_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_5_SFF_1_n10), .B2(key3FF_outputPar[13]), .C1(
        key3FF_keystate_gff_5_SFF_1_n11), .C2(key3FF_counterAdd[2]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_5_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_5_SFF_1_U3 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_5_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_5_SFF_1_U2 ( .A(key3FF_keystate_gff_5_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_5_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_5_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_5_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[17]), 
        .QN(key3FF_keystate_gff_5_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_5_SFF_2_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_5_SFF_2_n8), .A(key3FF_keystate_gff_5_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_5_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_5_SFF_2_U3 ( .B1(key3FF_keystate_n14), .B2(
        key3FF_outputPar[14]), .C1(key3FF_keystate_gff_5_SFF_2_n10), .C2(
        key3FF_counterAdd[3]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_5_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_5_SFF_2_U2 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_5_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_5_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_5_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[18]), 
        .QN(key3FF_keystate_gff_5_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_5_SFF_3_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_5_SFF_3_n8), .A(key3FF_keystate_gff_5_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_5_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_5_SFF_3_U3 ( .B1(key3FF_keystate_n14), .B2(
        key3FF_outputPar[15]), .C1(key3FF_keystate_gff_5_SFF_3_n10), .C2(
        key3FF_counterAdd[4]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_5_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_5_SFF_3_U2 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_5_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_5_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_5_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[19]), 
        .QN(key3FF_keystate_gff_5_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_6_SFF_0_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_6_SFF_0_n8), .A(key3FF_keystate_gff_6_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_6_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_6_SFF_0_U3 ( .B1(key3FF_keystate_n14), .B2(
        key3FF_outputPar[16]), .C1(key3FF_keystate_gff_6_SFF_0_n10), .C2(
        key3FF_outputPar[23]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_6_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_6_SFF_0_U2 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_6_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_6_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_6_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[20]), 
        .QN(key3FF_keystate_gff_6_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_6_SFF_1_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_6_SFF_1_n8), .A(key3FF_keystate_gff_6_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_6_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_6_SFF_1_U3 ( .B1(key3FF_keystate_n14), .B2(
        key3FF_outputPar[17]), .C1(key3FF_keystate_gff_6_SFF_1_n10), .C2(
        key3FF_outputPar[24]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_6_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_6_SFF_1_U2 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_6_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_6_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_6_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[21]), 
        .QN(key3FF_keystate_gff_6_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_6_SFF_2_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_6_SFF_2_n8), .A(key3FF_keystate_gff_6_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_6_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_6_SFF_2_U3 ( .B1(key3FF_keystate_n14), .B2(
        key3FF_outputPar[18]), .C1(key3FF_keystate_gff_6_SFF_2_n10), .C2(
        key3FF_outputPar[25]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_6_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_6_SFF_2_U2 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_6_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_6_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_6_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[22]), 
        .QN(key3FF_keystate_gff_6_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_6_SFF_3_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_6_SFF_3_n8), .A(key3FF_keystate_gff_6_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_6_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_6_SFF_3_U3 ( .B1(key3FF_keystate_n14), .B2(
        key3FF_outputPar[19]), .C1(key3FF_keystate_gff_6_SFF_3_n10), .C2(
        key3FF_outputPar[26]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_6_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_6_SFF_3_U2 ( .A(key3FF_keystate_n14), .ZN(
        key3FF_keystate_gff_6_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_6_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_6_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[23]), 
        .QN(key3FF_keystate_gff_6_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_7_SFF_0_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_7_SFF_0_n8), .A(key3FF_keystate_gff_7_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_7_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_7_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_7_SFF_0_n10), .B2(key3FF_outputPar[20]), .C1(
        key3FF_keystate_gff_7_SFF_0_n11), .C2(key3FF_outputPar[27]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_7_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_7_SFF_0_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_7_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_7_SFF_0_U2 ( .A(key3FF_keystate_gff_7_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_7_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_7_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_7_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[24]), 
        .QN(key3FF_keystate_gff_7_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_7_SFF_1_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_7_SFF_1_n8), .A(key3FF_keystate_gff_7_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_7_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_7_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_7_SFF_1_n10), .B2(key3FF_outputPar[21]), .C1(
        key3FF_keystate_gff_7_SFF_1_n11), .C2(key3FF_outputPar[28]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_7_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_7_SFF_1_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_7_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_7_SFF_1_U2 ( .A(key3FF_keystate_gff_7_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_7_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_7_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_7_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[25]), 
        .QN(key3FF_keystate_gff_7_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_7_SFF_2_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_7_SFF_2_n7), .A(key3FF_keystate_gff_7_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_7_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_7_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_7_SFF_2_n9), .B2(key3FF_outputPar[22]), .C1(
        key3FF_keystate_gff_7_SFF_2_n10), .C2(key3FF_outputPar[29]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_7_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_7_SFF_2_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_7_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_7_SFF_2_U2 ( .A(key3FF_keystate_gff_7_SFF_2_n10), 
        .ZN(key3FF_keystate_gff_7_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_7_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_7_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[26]), 
        .QN(key3FF_keystate_gff_7_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_7_SFF_3_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_7_SFF_3_n7), .A(key3FF_keystate_gff_7_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_7_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_7_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_7_SFF_3_n9), .B2(key3FF_outputPar[23]), .C1(
        key3FF_keystate_gff_7_SFF_3_n10), .C2(key3FF_outputPar[30]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_7_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_7_SFF_3_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_7_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_7_SFF_3_U2 ( .A(key3FF_keystate_gff_7_SFF_3_n10), 
        .ZN(key3FF_keystate_gff_7_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_7_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_7_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[27]), 
        .QN(key3FF_keystate_gff_7_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_8_SFF_0_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_8_SFF_0_n7), .A(key3FF_keystate_gff_8_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_8_SFF_0_n6) );
  OAI221_X1 key3FF_keystate_gff_8_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_8_SFF_0_n9), .B2(key3FF_outputPar[24]), .C1(
        key3FF_keystate_gff_8_SFF_0_n10), .C2(key3FF_outputPar[31]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_8_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_8_SFF_0_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_8_SFF_0_n10) );
  INV_X1 key3FF_keystate_gff_8_SFF_0_U2 ( .A(key3FF_keystate_gff_8_SFF_0_n10), 
        .ZN(key3FF_keystate_gff_8_SFF_0_n9) );
  DFF_X1 key3FF_keystate_gff_8_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_8_SFF_0_n6), .CK(clk), .Q(key3FF_outputPar[28]), 
        .QN(key3FF_keystate_gff_8_SFF_0_n7) );
  OAI21_X1 key3FF_keystate_gff_8_SFF_1_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_8_SFF_1_n7), .A(key3FF_keystate_gff_8_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_8_SFF_1_n6) );
  OAI221_X1 key3FF_keystate_gff_8_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_8_SFF_1_n9), .B2(key3FF_outputPar[25]), .C1(
        key3FF_keystate_gff_8_SFF_1_n10), .C2(key3FF_outputPar[32]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_8_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_8_SFF_1_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_8_SFF_1_n10) );
  INV_X1 key3FF_keystate_gff_8_SFF_1_U2 ( .A(key3FF_keystate_gff_8_SFF_1_n10), 
        .ZN(key3FF_keystate_gff_8_SFF_1_n9) );
  DFF_X1 key3FF_keystate_gff_8_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_8_SFF_1_n6), .CK(clk), .Q(key3FF_outputPar[29]), 
        .QN(key3FF_keystate_gff_8_SFF_1_n7) );
  OAI21_X1 key3FF_keystate_gff_8_SFF_2_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_8_SFF_2_n7), .A(key3FF_keystate_gff_8_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_8_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_8_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_8_SFF_2_n9), .B2(key3FF_outputPar[26]), .C1(
        key3FF_keystate_gff_8_SFF_2_n10), .C2(key3FF_outputPar[33]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_8_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_8_SFF_2_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_8_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_8_SFF_2_U2 ( .A(key3FF_keystate_gff_8_SFF_2_n10), 
        .ZN(key3FF_keystate_gff_8_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_8_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_8_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[30]), 
        .QN(key3FF_keystate_gff_8_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_8_SFF_3_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_8_SFF_3_n7), .A(key3FF_keystate_gff_8_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_8_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_8_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_8_SFF_3_n9), .B2(key3FF_outputPar[27]), .C1(
        key3FF_keystate_gff_8_SFF_3_n10), .C2(key3FF_outputPar[34]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_8_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_8_SFF_3_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_8_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_8_SFF_3_U2 ( .A(key3FF_keystate_gff_8_SFF_3_n10), 
        .ZN(key3FF_keystate_gff_8_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_8_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_8_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[31]), 
        .QN(key3FF_keystate_gff_8_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_9_SFF_0_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_9_SFF_0_n8), .A(key3FF_keystate_gff_9_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_9_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_9_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_9_SFF_0_n10), .B2(key3FF_outputPar[28]), .C1(
        key3FF_keystate_gff_9_SFF_0_n11), .C2(key3FF_outputPar[35]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_9_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_9_SFF_0_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_9_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_9_SFF_0_U2 ( .A(key3FF_keystate_gff_9_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_9_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_9_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_9_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[32]), 
        .QN(key3FF_keystate_gff_9_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_9_SFF_1_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_9_SFF_1_n8), .A(key3FF_keystate_gff_9_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_9_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_9_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_9_SFF_1_n10), .B2(key3FF_outputPar[29]), .C1(
        key3FF_keystate_gff_9_SFF_1_n11), .C2(key3FF_outputPar[36]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_9_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_9_SFF_1_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_9_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_9_SFF_1_U2 ( .A(key3FF_keystate_gff_9_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_9_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_9_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_9_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[33]), 
        .QN(key3FF_keystate_gff_9_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_9_SFF_2_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_9_SFF_2_n8), .A(key3FF_keystate_gff_9_SFF_2_n12), 
        .ZN(key3FF_keystate_gff_9_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_9_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_9_SFF_2_n10), .B2(key3FF_outputPar[30]), .C1(
        key3FF_keystate_gff_9_SFF_2_n11), .C2(key3FF_outputPar[37]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_9_SFF_2_n12) );
  INV_X1 key3FF_keystate_gff_9_SFF_2_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_9_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_9_SFF_2_U2 ( .A(key3FF_keystate_gff_9_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_9_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_9_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_9_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[34]), 
        .QN(key3FF_keystate_gff_9_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_9_SFF_3_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_9_SFF_3_n8), .A(key3FF_keystate_gff_9_SFF_3_n12), 
        .ZN(key3FF_keystate_gff_9_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_9_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_9_SFF_3_n10), .B2(key3FF_outputPar[31]), .C1(
        key3FF_keystate_gff_9_SFF_3_n11), .C2(key3FF_outputPar[38]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_9_SFF_3_n12) );
  INV_X1 key3FF_keystate_gff_9_SFF_3_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_9_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_9_SFF_3_U2 ( .A(key3FF_keystate_gff_9_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_9_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_9_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_9_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[35]), 
        .QN(key3FF_keystate_gff_9_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_10_SFF_0_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_10_SFF_0_n8), .A(key3FF_keystate_gff_10_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_10_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_10_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_10_SFF_0_n10), .B2(key3FF_outputPar[32]), .C1(
        key3FF_keystate_gff_10_SFF_0_n11), .C2(key3FF_outputPar[39]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_10_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_10_SFF_0_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_10_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_10_SFF_0_U2 ( .A(key3FF_keystate_gff_10_SFF_0_n11), .ZN(key3FF_keystate_gff_10_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_10_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_10_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[36]), 
        .QN(key3FF_keystate_gff_10_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_10_SFF_1_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_10_SFF_1_n8), .A(key3FF_keystate_gff_10_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_10_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_10_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_10_SFF_1_n10), .B2(key3FF_outputPar[33]), .C1(
        key3FF_keystate_gff_10_SFF_1_n11), .C2(key3FF_outputPar[40]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_10_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_10_SFF_1_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_10_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_10_SFF_1_U2 ( .A(key3FF_keystate_gff_10_SFF_1_n11), .ZN(key3FF_keystate_gff_10_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_10_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_10_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[37]), 
        .QN(key3FF_keystate_gff_10_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_10_SFF_2_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_10_SFF_2_n8), .A(key3FF_keystate_gff_10_SFF_2_n12), 
        .ZN(key3FF_keystate_gff_10_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_10_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_10_SFF_2_n10), .B2(key3FF_outputPar[34]), .C1(
        key3FF_keystate_gff_10_SFF_2_n11), .C2(key3FF_outputPar[41]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_10_SFF_2_n12) );
  INV_X1 key3FF_keystate_gff_10_SFF_2_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_10_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_10_SFF_2_U2 ( .A(key3FF_keystate_gff_10_SFF_2_n11), .ZN(key3FF_keystate_gff_10_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_10_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_10_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[38]), 
        .QN(key3FF_keystate_gff_10_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_10_SFF_3_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_10_SFF_3_n8), .A(key3FF_keystate_gff_10_SFF_3_n12), 
        .ZN(key3FF_keystate_gff_10_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_10_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_10_SFF_3_n10), .B2(key3FF_outputPar[35]), .C1(
        key3FF_keystate_gff_10_SFF_3_n11), .C2(key3FF_outputPar[42]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_10_SFF_3_n12) );
  INV_X1 key3FF_keystate_gff_10_SFF_3_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_10_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_10_SFF_3_U2 ( .A(key3FF_keystate_gff_10_SFF_3_n11), .ZN(key3FF_keystate_gff_10_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_10_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_10_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[39]), 
        .QN(key3FF_keystate_gff_10_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_11_SFF_0_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_11_SFF_0_n8), .A(key3FF_keystate_gff_11_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_11_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_11_SFF_0_U3 ( .B1(key3FF_keystate_n17), .B2(
        key3FF_outputPar[36]), .C1(key3FF_keystate_gff_11_SFF_0_n10), .C2(
        key3FF_outputPar[43]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_11_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_11_SFF_0_U2 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_11_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_11_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_11_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[40]), 
        .QN(key3FF_keystate_gff_11_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_11_SFF_1_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_11_SFF_1_n8), .A(key3FF_keystate_gff_11_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_11_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_11_SFF_1_U3 ( .B1(key3FF_keystate_n17), .B2(
        key3FF_outputPar[37]), .C1(key3FF_keystate_gff_11_SFF_1_n10), .C2(
        key3FF_outputPar[44]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_11_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_11_SFF_1_U2 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_11_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_11_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_11_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[41]), 
        .QN(key3FF_keystate_gff_11_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_11_SFF_2_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_11_SFF_2_n7), .A(key3FF_keystate_gff_11_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_11_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_11_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_11_SFF_2_n9), .B2(key3FF_outputPar[38]), .C1(
        key3FF_keystate_gff_11_SFF_2_n10), .C2(key3FF_outputPar[45]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_11_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_11_SFF_2_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_11_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_11_SFF_2_U2 ( .A(key3FF_keystate_gff_11_SFF_2_n10), .ZN(key3FF_keystate_gff_11_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_11_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_11_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[42]), 
        .QN(key3FF_keystate_gff_11_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_11_SFF_3_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_11_SFF_3_n7), .A(key3FF_keystate_gff_11_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_11_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_11_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_11_SFF_3_n9), .B2(key3FF_outputPar[39]), .C1(
        key3FF_keystate_gff_11_SFF_3_n10), .C2(key3FF_outputPar[46]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_11_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_11_SFF_3_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_11_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_11_SFF_3_U2 ( .A(key3FF_keystate_gff_11_SFF_3_n10), .ZN(key3FF_keystate_gff_11_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_11_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_11_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[43]), 
        .QN(key3FF_keystate_gff_11_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_12_SFF_0_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_12_SFF_0_n7), .A(key3FF_keystate_gff_12_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_12_SFF_0_n6) );
  OAI221_X1 key3FF_keystate_gff_12_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_12_SFF_0_n9), .B2(key3FF_outputPar[40]), .C1(
        key3FF_keystate_gff_12_SFF_0_n10), .C2(key3FF_outputPar[47]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_12_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_12_SFF_0_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_12_SFF_0_n10) );
  INV_X1 key3FF_keystate_gff_12_SFF_0_U2 ( .A(key3FF_keystate_gff_12_SFF_0_n10), .ZN(key3FF_keystate_gff_12_SFF_0_n9) );
  DFF_X1 key3FF_keystate_gff_12_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_12_SFF_0_n6), .CK(clk), .Q(key3FF_outputPar[44]), 
        .QN(key3FF_keystate_gff_12_SFF_0_n7) );
  OAI21_X1 key3FF_keystate_gff_12_SFF_1_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_12_SFF_1_n7), .A(key3FF_keystate_gff_12_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_12_SFF_1_n6) );
  OAI221_X1 key3FF_keystate_gff_12_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_12_SFF_1_n9), .B2(key3FF_outputPar[41]), .C1(
        key3FF_keystate_gff_12_SFF_1_n10), .C2(key3FF_outputPar[48]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_12_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_12_SFF_1_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_12_SFF_1_n10) );
  INV_X1 key3FF_keystate_gff_12_SFF_1_U2 ( .A(key3FF_keystate_gff_12_SFF_1_n10), .ZN(key3FF_keystate_gff_12_SFF_1_n9) );
  DFF_X1 key3FF_keystate_gff_12_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_12_SFF_1_n6), .CK(clk), .Q(key3FF_outputPar[45]), 
        .QN(key3FF_keystate_gff_12_SFF_1_n7) );
  OAI21_X1 key3FF_keystate_gff_12_SFF_2_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_12_SFF_2_n7), .A(key3FF_keystate_gff_12_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_12_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_12_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_12_SFF_2_n9), .B2(key3FF_outputPar[42]), .C1(
        key3FF_keystate_gff_12_SFF_2_n10), .C2(key3FF_outputPar[49]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_12_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_12_SFF_2_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_12_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_12_SFF_2_U2 ( .A(key3FF_keystate_gff_12_SFF_2_n10), .ZN(key3FF_keystate_gff_12_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_12_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_12_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[46]), 
        .QN(key3FF_keystate_gff_12_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_12_SFF_3_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_12_SFF_3_n7), .A(key3FF_keystate_gff_12_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_12_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_12_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_12_SFF_3_n9), .B2(key3FF_outputPar[43]), .C1(
        key3FF_keystate_gff_12_SFF_3_n10), .C2(key3FF_outputPar[50]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_12_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_12_SFF_3_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_12_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_12_SFF_3_U2 ( .A(key3FF_keystate_gff_12_SFF_3_n10), .ZN(key3FF_keystate_gff_12_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_12_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_12_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[47]), 
        .QN(key3FF_keystate_gff_12_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_13_SFF_0_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_13_SFF_0_n8), .A(key3FF_keystate_gff_13_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_13_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_13_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_13_SFF_0_n10), .B2(key3FF_outputPar[44]), .C1(
        key3FF_keystate_gff_13_SFF_0_n11), .C2(key3FF_outputPar[51]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_13_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_13_SFF_0_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_13_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_13_SFF_0_U2 ( .A(key3FF_keystate_gff_13_SFF_0_n11), .ZN(key3FF_keystate_gff_13_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_13_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_13_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[48]), 
        .QN(key3FF_keystate_gff_13_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_13_SFF_1_U5 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_13_SFF_1_n8), .A(key3FF_keystate_gff_13_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_13_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_13_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_13_SFF_1_n10), .B2(key3FF_outputPar[45]), .C1(
        key3FF_keystate_gff_13_SFF_1_n11), .C2(key3FF_outputPar[52]), .A(
        key3FF_keystate_n10), .ZN(key3FF_keystate_gff_13_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_13_SFF_1_U3 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_13_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_13_SFF_1_U2 ( .A(key3FF_keystate_gff_13_SFF_1_n11), .ZN(key3FF_keystate_gff_13_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_13_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_13_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[49]), 
        .QN(key3FF_keystate_gff_13_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_13_SFF_2_U4 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_13_SFF_2_n8), .A(key3FF_keystate_gff_13_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_13_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_13_SFF_2_U3 ( .B1(key3FF_keystate_n15), .B2(
        key3FF_outputPar[46]), .C1(key3FF_keystate_gff_13_SFF_2_n10), .C2(
        key3FF_outputPar[53]), .A(key3FF_keystate_n10), .ZN(
        key3FF_keystate_gff_13_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_13_SFF_2_U2 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_13_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_13_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_13_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[50]), 
        .QN(key3FF_keystate_gff_13_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_13_SFF_3_U4 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_13_SFF_3_n8), .A(key3FF_keystate_gff_13_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_13_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_13_SFF_3_U3 ( .B1(key3FF_keystate_n15), .B2(
        key3FF_outputPar[47]), .C1(key3FF_keystate_gff_13_SFF_3_n10), .C2(
        key3FF_outputPar[54]), .A(key3FF_keystate_n10), .ZN(
        key3FF_keystate_gff_13_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_13_SFF_3_U2 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_13_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_13_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_13_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[51]), 
        .QN(key3FF_keystate_gff_13_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_14_SFF_0_U4 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_14_SFF_0_n8), .A(key3FF_keystate_gff_14_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_14_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_14_SFF_0_U3 ( .B1(key3FF_keystate_n15), .B2(
        key3FF_outputPar[48]), .C1(key3FF_keystate_gff_14_SFF_0_n10), .C2(
        key3FF_outputPar[55]), .A(key3FF_keystate_n10), .ZN(
        key3FF_keystate_gff_14_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_14_SFF_0_U2 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_14_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_14_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_14_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[52]), 
        .QN(key3FF_keystate_gff_14_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_14_SFF_1_U4 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_14_SFF_1_n8), .A(key3FF_keystate_gff_14_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_14_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_14_SFF_1_U3 ( .B1(key3FF_keystate_n15), .B2(
        key3FF_outputPar[49]), .C1(key3FF_keystate_gff_14_SFF_1_n10), .C2(
        key3FF_outputPar[56]), .A(key3FF_keystate_n10), .ZN(
        key3FF_keystate_gff_14_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_14_SFF_1_U2 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_14_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_14_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_14_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[53]), 
        .QN(key3FF_keystate_gff_14_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_14_SFF_2_U4 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_14_SFF_2_n8), .A(key3FF_keystate_gff_14_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_14_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_14_SFF_2_U3 ( .B1(key3FF_keystate_n15), .B2(
        key3FF_outputPar[50]), .C1(key3FF_keystate_gff_14_SFF_2_n10), .C2(
        key3FF_outputPar[57]), .A(key3FF_keystate_n10), .ZN(
        key3FF_keystate_gff_14_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_14_SFF_2_U2 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_14_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_14_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_14_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[54]), 
        .QN(key3FF_keystate_gff_14_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_14_SFF_3_U4 ( .B1(key3FF_keystate_n10), .B2(
        key3FF_keystate_gff_14_SFF_3_n8), .A(key3FF_keystate_gff_14_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_14_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_14_SFF_3_U3 ( .B1(key3FF_keystate_n15), .B2(
        key3FF_outputPar[51]), .C1(key3FF_keystate_gff_14_SFF_3_n10), .C2(
        key3FF_outputPar[58]), .A(key3FF_keystate_n10), .ZN(
        key3FF_keystate_gff_14_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_14_SFF_3_U2 ( .A(key3FF_keystate_n15), .ZN(
        key3FF_keystate_gff_14_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_14_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_14_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[55]), 
        .QN(key3FF_keystate_gff_14_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_15_SFF_0_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_15_SFF_0_n8), .A(key3FF_keystate_gff_15_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_15_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_15_SFF_0_U3 ( .B1(key3FF_keystate_n17), .B2(
        key3FF_outputPar[52]), .C1(key3FF_keystate_gff_15_SFF_0_n10), .C2(
        key3FF_outputPar[59]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_15_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_15_SFF_0_U2 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_15_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_15_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_15_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[56]), 
        .QN(key3FF_keystate_gff_15_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_15_SFF_1_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_15_SFF_1_n8), .A(key3FF_keystate_gff_15_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_15_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_15_SFF_1_U3 ( .B1(key3FF_keystate_n17), .B2(
        key3FF_outputPar[53]), .C1(key3FF_keystate_gff_15_SFF_1_n10), .C2(
        key3FF_outputPar[60]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_15_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_15_SFF_1_U2 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_15_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_15_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_15_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[57]), 
        .QN(key3FF_keystate_gff_15_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_15_SFF_2_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_15_SFF_2_n7), .A(key3FF_keystate_gff_15_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_15_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_15_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_15_SFF_2_n9), .B2(key3FF_outputPar[54]), .C1(
        key3FF_keystate_gff_15_SFF_2_n10), .C2(key3FF_outputPar[61]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_15_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_15_SFF_2_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_15_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_15_SFF_2_U2 ( .A(key3FF_keystate_gff_15_SFF_2_n10), .ZN(key3FF_keystate_gff_15_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_15_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_15_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[58]), 
        .QN(key3FF_keystate_gff_15_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_15_SFF_3_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_15_SFF_3_n7), .A(key3FF_keystate_gff_15_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_15_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_15_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_15_SFF_3_n9), .B2(key3FF_outputPar[55]), .C1(
        key3FF_keystate_gff_15_SFF_3_n10), .C2(key3FF_outputPar[62]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_15_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_15_SFF_3_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_15_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_15_SFF_3_U2 ( .A(key3FF_keystate_gff_15_SFF_3_n10), .ZN(key3FF_keystate_gff_15_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_15_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_15_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[59]), 
        .QN(key3FF_keystate_gff_15_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_16_SFF_0_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_16_SFF_0_n7), .A(key3FF_keystate_gff_16_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_16_SFF_0_n6) );
  OAI221_X1 key3FF_keystate_gff_16_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_16_SFF_0_n9), .B2(key3FF_outputPar[56]), .C1(
        key3FF_keystate_gff_16_SFF_0_n10), .C2(key3FF_outputPar[63]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_16_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_16_SFF_0_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_16_SFF_0_n10) );
  INV_X1 key3FF_keystate_gff_16_SFF_0_U2 ( .A(key3FF_keystate_gff_16_SFF_0_n10), .ZN(key3FF_keystate_gff_16_SFF_0_n9) );
  DFF_X1 key3FF_keystate_gff_16_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_16_SFF_0_n6), .CK(clk), .Q(key3FF_outputPar[60]), 
        .QN(key3FF_keystate_gff_16_SFF_0_n7) );
  OAI21_X1 key3FF_keystate_gff_16_SFF_1_U5 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_16_SFF_1_n7), .A(key3FF_keystate_gff_16_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_16_SFF_1_n6) );
  OAI221_X1 key3FF_keystate_gff_16_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_16_SFF_1_n9), .B2(key3FF_outputPar[57]), .C1(
        key3FF_keystate_gff_16_SFF_1_n10), .C2(key3FF_outputPar[64]), .A(
        key3FF_keystate_n13), .ZN(key3FF_keystate_gff_16_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_16_SFF_1_U3 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_16_SFF_1_n10) );
  INV_X1 key3FF_keystate_gff_16_SFF_1_U2 ( .A(key3FF_keystate_gff_16_SFF_1_n10), .ZN(key3FF_keystate_gff_16_SFF_1_n9) );
  DFF_X1 key3FF_keystate_gff_16_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_16_SFF_1_n6), .CK(clk), .Q(key3FF_outputPar[61]), 
        .QN(key3FF_keystate_gff_16_SFF_1_n7) );
  OAI21_X1 key3FF_keystate_gff_16_SFF_2_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_16_SFF_2_n7), .A(key3FF_keystate_gff_16_SFF_2_n10), 
        .ZN(key3FF_keystate_gff_16_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_16_SFF_2_U3 ( .B1(key3FF_keystate_n18), .B2(
        key3FF_outputPar[58]), .C1(key3FF_keystate_gff_16_SFF_2_n9), .C2(
        key3FF_outputPar[65]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_16_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_16_SFF_2_U2 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_16_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_16_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_16_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[62]), 
        .QN(key3FF_keystate_gff_16_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_16_SFF_3_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_16_SFF_3_n7), .A(key3FF_keystate_gff_16_SFF_3_n10), 
        .ZN(key3FF_keystate_gff_16_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_16_SFF_3_U3 ( .B1(key3FF_keystate_n18), .B2(
        key3FF_outputPar[59]), .C1(key3FF_keystate_gff_16_SFF_3_n9), .C2(
        key3FF_outputPar[66]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_16_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_16_SFF_3_U2 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_16_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_16_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_16_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[63]), 
        .QN(key3FF_keystate_gff_16_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_17_SFF_0_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_17_SFF_0_n8), .A(key3FF_keystate_gff_17_SFF_0_n12), 
        .ZN(key3FF_keystate_gff_17_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_17_SFF_0_U4 ( .B1(
        key3FF_keystate_gff_17_SFF_0_n10), .B2(key3FF_outputPar[60]), .C1(
        key3FF_keystate_gff_17_SFF_0_n11), .C2(key3FF_outputPar[67]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_17_SFF_0_n12) );
  INV_X1 key3FF_keystate_gff_17_SFF_0_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_17_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_17_SFF_0_U2 ( .A(key3FF_keystate_gff_17_SFF_0_n11), .ZN(key3FF_keystate_gff_17_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_17_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_17_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[64]), 
        .QN(key3FF_keystate_gff_17_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_17_SFF_1_U5 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_17_SFF_1_n8), .A(key3FF_keystate_gff_17_SFF_1_n12), 
        .ZN(key3FF_keystate_gff_17_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_17_SFF_1_U4 ( .B1(
        key3FF_keystate_gff_17_SFF_1_n10), .B2(key3FF_outputPar[61]), .C1(
        key3FF_keystate_gff_17_SFF_1_n11), .C2(key3FF_outputPar[68]), .A(
        key3FF_keystate_n11), .ZN(key3FF_keystate_gff_17_SFF_1_n12) );
  INV_X1 key3FF_keystate_gff_17_SFF_1_U3 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_17_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_17_SFF_1_U2 ( .A(key3FF_keystate_gff_17_SFF_1_n11), .ZN(key3FF_keystate_gff_17_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_17_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_17_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[65]), 
        .QN(key3FF_keystate_gff_17_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_17_SFF_2_U4 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_17_SFF_2_n8), .A(key3FF_keystate_gff_17_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_17_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_17_SFF_2_U3 ( .B1(key3FF_keystate_n16), .B2(
        key3FF_outputPar[62]), .C1(key3FF_keystate_gff_17_SFF_2_n10), .C2(
        key3FF_outputPar[69]), .A(key3FF_keystate_n11), .ZN(
        key3FF_keystate_gff_17_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_17_SFF_2_U2 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_17_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_17_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_17_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[66]), 
        .QN(key3FF_keystate_gff_17_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_17_SFF_3_U4 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_17_SFF_3_n8), .A(key3FF_keystate_gff_17_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_17_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_17_SFF_3_U3 ( .B1(key3FF_keystate_n16), .B2(
        key3FF_outputPar[63]), .C1(key3FF_keystate_gff_17_SFF_3_n10), .C2(
        key3FF_outputPar[70]), .A(key3FF_keystate_n11), .ZN(
        key3FF_keystate_gff_17_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_17_SFF_3_U2 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_17_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_17_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_17_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[67]), 
        .QN(key3FF_keystate_gff_17_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_18_SFF_0_U4 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_18_SFF_0_n8), .A(key3FF_keystate_gff_18_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_18_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_18_SFF_0_U3 ( .B1(key3FF_keystate_n16), .B2(
        key3FF_outputPar[64]), .C1(key3FF_keystate_gff_18_SFF_0_n10), .C2(
        key3FF_outputPar[71]), .A(key3FF_keystate_n11), .ZN(
        key3FF_keystate_gff_18_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_18_SFF_0_U2 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_18_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_18_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_18_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[68]), 
        .QN(key3FF_keystate_gff_18_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_18_SFF_1_U4 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_18_SFF_1_n8), .A(key3FF_keystate_gff_18_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_18_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_18_SFF_1_U3 ( .B1(key3FF_keystate_n16), .B2(
        key3FF_outputPar[65]), .C1(key3FF_keystate_gff_18_SFF_1_n10), .C2(
        key3FF_outputPar[72]), .A(key3FF_keystate_n11), .ZN(
        key3FF_keystate_gff_18_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_18_SFF_1_U2 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_18_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_18_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_18_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[69]), 
        .QN(key3FF_keystate_gff_18_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_18_SFF_2_U4 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_18_SFF_2_n8), .A(key3FF_keystate_gff_18_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_18_SFF_2_n7) );
  OAI221_X1 key3FF_keystate_gff_18_SFF_2_U3 ( .B1(key3FF_keystate_n16), .B2(
        key3FF_outputPar[66]), .C1(key3FF_keystate_gff_18_SFF_2_n10), .C2(
        key3FF_outputPar[73]), .A(key3FF_keystate_n11), .ZN(
        key3FF_keystate_gff_18_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_18_SFF_2_U2 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_18_SFF_2_n10) );
  DFF_X1 key3FF_keystate_gff_18_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_18_SFF_2_n7), .CK(clk), .Q(key3FF_outputPar[70]), 
        .QN(key3FF_keystate_gff_18_SFF_2_n8) );
  OAI21_X1 key3FF_keystate_gff_18_SFF_3_U4 ( .B1(key3FF_keystate_n11), .B2(
        key3FF_keystate_gff_18_SFF_3_n8), .A(key3FF_keystate_gff_18_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_18_SFF_3_n7) );
  OAI221_X1 key3FF_keystate_gff_18_SFF_3_U3 ( .B1(key3FF_keystate_n16), .B2(
        key3FF_outputPar[67]), .C1(key3FF_keystate_gff_18_SFF_3_n10), .C2(
        key3FF_outputPar[74]), .A(key3FF_keystate_n11), .ZN(
        key3FF_keystate_gff_18_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_18_SFF_3_U2 ( .A(key3FF_keystate_n16), .ZN(
        key3FF_keystate_gff_18_SFF_3_n10) );
  DFF_X1 key3FF_keystate_gff_18_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_18_SFF_3_n7), .CK(clk), .Q(key3FF_outputPar[71]), 
        .QN(key3FF_keystate_gff_18_SFF_3_n8) );
  OAI21_X1 key3FF_keystate_gff_19_SFF_0_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_19_SFF_0_n8), .A(key3FF_keystate_gff_19_SFF_0_n11), 
        .ZN(key3FF_keystate_gff_19_SFF_0_n7) );
  OAI221_X1 key3FF_keystate_gff_19_SFF_0_U3 ( .B1(key3FF_keystate_n17), .B2(
        key3FF_outputPar[68]), .C1(key3FF_keystate_gff_19_SFF_0_n10), .C2(
        key3FF_outputPar[75]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_19_SFF_0_n11) );
  INV_X1 key3FF_keystate_gff_19_SFF_0_U2 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_19_SFF_0_n10) );
  DFF_X1 key3FF_keystate_gff_19_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_19_SFF_0_n7), .CK(clk), .Q(key3FF_outputPar[72]), 
        .QN(key3FF_keystate_gff_19_SFF_0_n8) );
  OAI21_X1 key3FF_keystate_gff_19_SFF_1_U4 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_19_SFF_1_n8), .A(key3FF_keystate_gff_19_SFF_1_n11), 
        .ZN(key3FF_keystate_gff_19_SFF_1_n7) );
  OAI221_X1 key3FF_keystate_gff_19_SFF_1_U3 ( .B1(key3FF_keystate_n17), .B2(
        key3FF_outputPar[69]), .C1(key3FF_keystate_gff_19_SFF_1_n10), .C2(
        roundkey3[0]), .A(key3FF_keystate_n12), .ZN(
        key3FF_keystate_gff_19_SFF_1_n11) );
  INV_X1 key3FF_keystate_gff_19_SFF_1_U2 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_19_SFF_1_n10) );
  DFF_X1 key3FF_keystate_gff_19_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_19_SFF_1_n7), .CK(clk), .Q(key3FF_outputPar[73]), 
        .QN(key3FF_keystate_gff_19_SFF_1_n8) );
  OAI21_X1 key3FF_keystate_gff_19_SFF_2_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_19_SFF_2_n7), .A(key3FF_keystate_gff_19_SFF_2_n11), 
        .ZN(key3FF_keystate_gff_19_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_19_SFF_2_U4 ( .B1(
        key3FF_keystate_gff_19_SFF_2_n9), .B2(key3FF_outputPar[70]), .C1(
        key3FF_keystate_gff_19_SFF_2_n10), .C2(roundkey3[1]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_19_SFF_2_n11) );
  INV_X1 key3FF_keystate_gff_19_SFF_2_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_19_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_19_SFF_2_U2 ( .A(key3FF_keystate_gff_19_SFF_2_n10), .ZN(key3FF_keystate_gff_19_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_19_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_19_SFF_2_n6), .CK(clk), .Q(key3FF_outputPar[74]), 
        .QN(key3FF_keystate_gff_19_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_19_SFF_3_U5 ( .B1(key3FF_keystate_n12), .B2(
        key3FF_keystate_gff_19_SFF_3_n7), .A(key3FF_keystate_gff_19_SFF_3_n11), 
        .ZN(key3FF_keystate_gff_19_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_19_SFF_3_U4 ( .B1(
        key3FF_keystate_gff_19_SFF_3_n9), .B2(key3FF_outputPar[71]), .C1(
        key3FF_keystate_gff_19_SFF_3_n10), .C2(roundkey3[2]), .A(
        key3FF_keystate_n12), .ZN(key3FF_keystate_gff_19_SFF_3_n11) );
  INV_X1 key3FF_keystate_gff_19_SFF_3_U3 ( .A(key3FF_keystate_n17), .ZN(
        key3FF_keystate_gff_19_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_19_SFF_3_U2 ( .A(key3FF_keystate_gff_19_SFF_3_n10), .ZN(key3FF_keystate_gff_19_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_19_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_19_SFF_3_n6), .CK(clk), .Q(key3FF_outputPar[75]), 
        .QN(key3FF_keystate_gff_19_SFF_3_n7) );
  OAI21_X1 key3FF_keystate_gff_20_SFF_0_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_20_SFF_0_n7), .A(key3FF_keystate_gff_20_SFF_0_n10), 
        .ZN(key3FF_keystate_gff_20_SFF_0_n6) );
  OAI221_X1 key3FF_keystate_gff_20_SFF_0_U3 ( .B1(key3FF_keystate_n18), .B2(
        key3FF_outputPar[72]), .C1(key3FF_keystate_gff_20_SFF_0_n9), .C2(
        sboxOut3[0]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_20_SFF_0_n10) );
  INV_X1 key3FF_keystate_gff_20_SFF_0_U2 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_20_SFF_0_n9) );
  DFF_X1 key3FF_keystate_gff_20_SFF_0_Cell_reg ( .D(
        key3FF_keystate_gff_20_SFF_0_n6), .CK(clk), .Q(roundkey3[0]), .QN(
        key3FF_keystate_gff_20_SFF_0_n7) );
  OAI21_X1 key3FF_keystate_gff_20_SFF_1_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_20_SFF_1_n7), .A(key3FF_keystate_gff_20_SFF_1_n10), 
        .ZN(key3FF_keystate_gff_20_SFF_1_n6) );
  OAI221_X1 key3FF_keystate_gff_20_SFF_1_U3 ( .B1(key3FF_keystate_n18), .B2(
        key3FF_outputPar[73]), .C1(key3FF_keystate_gff_20_SFF_1_n9), .C2(
        sboxOut3[1]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_20_SFF_1_n10) );
  INV_X1 key3FF_keystate_gff_20_SFF_1_U2 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_20_SFF_1_n9) );
  DFF_X1 key3FF_keystate_gff_20_SFF_1_Cell_reg ( .D(
        key3FF_keystate_gff_20_SFF_1_n6), .CK(clk), .Q(roundkey3[1]), .QN(
        key3FF_keystate_gff_20_SFF_1_n7) );
  OAI21_X1 key3FF_keystate_gff_20_SFF_2_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_20_SFF_2_n7), .A(key3FF_keystate_gff_20_SFF_2_n10), 
        .ZN(key3FF_keystate_gff_20_SFF_2_n6) );
  OAI221_X1 key3FF_keystate_gff_20_SFF_2_U3 ( .B1(key3FF_keystate_n18), .B2(
        key3FF_outputPar[74]), .C1(key3FF_keystate_gff_20_SFF_2_n9), .C2(
        sboxOut3[2]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_20_SFF_2_n10) );
  INV_X1 key3FF_keystate_gff_20_SFF_2_U2 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_20_SFF_2_n9) );
  DFF_X1 key3FF_keystate_gff_20_SFF_2_Cell_reg ( .D(
        key3FF_keystate_gff_20_SFF_2_n6), .CK(clk), .Q(roundkey3[2]), .QN(
        key3FF_keystate_gff_20_SFF_2_n7) );
  OAI21_X1 key3FF_keystate_gff_20_SFF_3_U4 ( .B1(key3FF_keystate_n13), .B2(
        key3FF_keystate_gff_20_SFF_3_n7), .A(key3FF_keystate_gff_20_SFF_3_n10), 
        .ZN(key3FF_keystate_gff_20_SFF_3_n6) );
  OAI221_X1 key3FF_keystate_gff_20_SFF_3_U3 ( .B1(key3FF_keystate_n18), .B2(
        key3FF_outputPar[75]), .C1(key3FF_keystate_gff_20_SFF_3_n9), .C2(
        sboxOut3[3]), .A(key3FF_keystate_n13), .ZN(
        key3FF_keystate_gff_20_SFF_3_n10) );
  INV_X1 key3FF_keystate_gff_20_SFF_3_U2 ( .A(key3FF_keystate_n18), .ZN(
        key3FF_keystate_gff_20_SFF_3_n9) );
  DFF_X1 key3FF_keystate_gff_20_SFF_3_Cell_reg ( .D(
        key3FF_keystate_gff_20_SFF_3_n6), .CK(clk), .Q(roundkey3[3]), .QN(
        key3FF_keystate_gff_20_SFF_3_n7) );
  MUX2_X1 mux1_U4 ( .A(roundkey1[3]), .B(AddKeyOut1[0]), .S(selSbox), .Z(
        dataOut1[0]) );
  MUX2_X1 mux1_U3 ( .A(keyRegKS1[1]), .B(AddKeyOut1[1]), .S(selSbox), .Z(
        dataOut1[1]) );
  MUX2_X1 mux1_U2 ( .A(keyRegKS1[2]), .B(AddKeyOut1[2]), .S(selSbox), .Z(
        dataOut1[2]) );
  MUX2_X1 mux1_U1 ( .A(keyRegKS1[3]), .B(AddKeyOut1[3]), .S(selSbox), .Z(
        dataOut1[3]) );
  MUX2_X1 mux2_U4 ( .A(roundkey2[3]), .B(AddKeyOut2[0]), .S(selSbox), .Z(
        dataOut2[0]) );
  MUX2_X1 mux2_U3 ( .A(keyRegKS2[1]), .B(AddKeyOut2[1]), .S(selSbox), .Z(
        dataOut2[1]) );
  MUX2_X1 mux2_U2 ( .A(keyRegKS2[2]), .B(AddKeyOut2[2]), .S(selSbox), .Z(
        dataOut2[2]) );
  MUX2_X1 mux2_U1 ( .A(keyRegKS2[3]), .B(AddKeyOut2[3]), .S(selSbox), .Z(
        dataOut2[3]) );
  MUX2_X1 mux3_U4 ( .A(roundkey3[3]), .B(AddKeyOut3[0]), .S(selSbox), .Z(
        dataOut3[0]) );
  MUX2_X1 mux3_U3 ( .A(keyRegKS3[1]), .B(AddKeyOut3[1]), .S(selSbox), .Z(
        dataOut3[1]) );
  MUX2_X1 mux3_U2 ( .A(keyRegKS3[2]), .B(AddKeyOut3[2]), .S(selSbox), .Z(
        dataOut3[2]) );
  MUX2_X1 mux3_U1 ( .A(keyRegKS3[3]), .B(AddKeyOut3[3]), .S(selSbox), .Z(
        dataOut3[3]) );
  DFF_X1 sbox_Rq1_reg_3_ ( .D(sbox_q1[3]), .CK(clk), .Q(sbox_Rq1[3]), .QN() );
  DFF_X1 sbox_Rq1_reg_2_ ( .D(sbox_q1[2]), .CK(clk), .Q(sbox_Rq1[2]), .QN() );
  DFF_X1 sbox_Rq1_reg_1_ ( .D(sbox_q1[1]), .CK(clk), .Q(sbox_Rq1[1]), .QN() );
  DFF_X1 sbox_Rq1_reg_0_ ( .D(sbox_q1[0]), .CK(clk), .Q(sbox_Rq1[0]), .QN() );
  DFF_X1 sbox_Rq2_reg_3_ ( .D(sbox_q2[3]), .CK(clk), .Q(sbox_Rq2[3]), .QN() );
  DFF_X1 sbox_Rq2_reg_2_ ( .D(sbox_q2[2]), .CK(clk), .Q(sbox_Rq2[2]), .QN() );
  DFF_X1 sbox_Rq2_reg_1_ ( .D(sbox_q2[1]), .CK(clk), .Q(sbox_Rq2[1]), .QN() );
  DFF_X1 sbox_Rq2_reg_0_ ( .D(sbox_q2[0]), .CK(clk), .Q(sbox_Rq2[0]), .QN() );
  DFF_X1 sbox_Rq3_reg_3_ ( .D(sbox_q3[3]), .CK(clk), .Q(sbox_Rq3[3]), .QN() );
  DFF_X1 sbox_Rq3_reg_2_ ( .D(sbox_q3[2]), .CK(clk), .Q(sbox_Rq3[2]), .QN() );
  DFF_X1 sbox_Rq3_reg_1_ ( .D(sbox_q3[1]), .CK(clk), .Q(sbox_Rq3[1]), .QN() );
  DFF_X1 sbox_Rq3_reg_0_ ( .D(sbox_q3[0]), .CK(clk), .Q(sbox_Rq3[0]), .QN() );
  DFF_X1 sbox_F_in3_reg_reg_0_ ( .D(dataOut3[0]), .CK(clk), .Q(
        sbox_F_in3_reg[0]), .QN() );
  DFF_X1 sbox_F_in3_reg_reg_1_ ( .D(dataOut3[3]), .CK(clk), .Q(
        sbox_F_in3_reg[1]), .QN() );
  DFF_X1 sbox_F_in3_reg_reg_2_ ( .D(dataOut3[1]), .CK(clk), .Q(
        sbox_F_in3_reg[2]), .QN() );
  DFF_X1 sbox_F_in3_reg_reg_3_ ( .D(sbox_F_in3_3_), .CK(clk), .Q(
        sbox_F_in3_reg[3]), .QN() );
  DFF_X1 sbox_F_in2_reg_reg_0_ ( .D(dataOut2[0]), .CK(clk), .Q(
        sbox_F_in2_reg[0]), .QN() );
  DFF_X1 sbox_F_in2_reg_reg_1_ ( .D(dataOut2[3]), .CK(clk), .Q(
        sbox_F_in2_reg[1]), .QN() );
  DFF_X1 sbox_F_in2_reg_reg_2_ ( .D(dataOut2[1]), .CK(clk), .Q(
        sbox_F_in2_reg[2]), .QN() );
  DFF_X1 sbox_F_in2_reg_reg_3_ ( .D(sbox_F_in2_3_), .CK(clk), .Q(
        sbox_F_in2_reg[3]), .QN() );
  DFF_X1 sbox_F_in1_reg_reg_0_ ( .D(dataOut1[0]), .CK(clk), .Q(
        sbox_F_in1_reg[0]), .QN() );
  DFF_X1 sbox_F_in1_reg_reg_1_ ( .D(dataOut1[3]), .CK(clk), .Q(
        sbox_F_in1_reg[1]), .QN() );
  DFF_X1 sbox_F_in1_reg_reg_2_ ( .D(dataOut1[1]), .CK(clk), .Q(
        sbox_F_in1_reg[2]), .QN() );
  DFF_X1 sbox_F_in1_reg_reg_3_ ( .D(sbox_F_in1_3_), .CK(clk), .Q(
        sbox_F_in1_reg[3]), .QN() );
  XOR2_X1 sbox_InputAffine_U3 ( .A(dataOut3[1]), .B(dataOut3[2]), .Z(
        sbox_F_in3_3_) );
  XOR2_X1 sbox_InputAffine_U2 ( .A(dataOut2[1]), .B(dataOut2[2]), .Z(
        sbox_F_in2_3_) );
  XNOR2_X1 sbox_InputAffine_U1 ( .A(dataOut1[1]), .B(dataOut1[2]), .ZN(
        sbox_F_in1_3_) );
  XNOR2_X1 sbox_F_U18 ( .A(sbox_F_n4), .B(r[3]), .ZN(sbox_q3[3]) );
  XNOR2_X1 sbox_F_U17 ( .A(r[2]), .B(sbox_F_q3[3]), .ZN(sbox_F_n4) );
  XNOR2_X1 sbox_F_U16 ( .A(sbox_F_n3), .B(r[1]), .ZN(sbox_q3[2]) );
  XNOR2_X1 sbox_F_U15 ( .A(r[0]), .B(sbox_F_q3[2]), .ZN(sbox_F_n3) );
  XNOR2_X1 sbox_F_U14 ( .A(sbox_F_n2), .B(r[7]), .ZN(sbox_q3[1]) );
  XNOR2_X1 sbox_F_U13 ( .A(r[6]), .B(sbox_F_q3[1]), .ZN(sbox_F_n2) );
  XNOR2_X1 sbox_F_U12 ( .A(sbox_F_n1), .B(r[5]), .ZN(sbox_q3[0]) );
  XNOR2_X1 sbox_F_U11 ( .A(r[4]), .B(sbox_F_q3[0]), .ZN(sbox_F_n1) );
  XOR2_X1 sbox_F_U10 ( .A(r[3]), .B(sbox_F_q2[3]), .Z(sbox_q2[3]) );
  XOR2_X1 sbox_F_U9 ( .A(r[1]), .B(sbox_F_q2[2]), .Z(sbox_q2[2]) );
  XOR2_X1 sbox_F_U8 ( .A(r[7]), .B(sbox_F_q2[1]), .Z(sbox_q2[1]) );
  XOR2_X1 sbox_F_U7 ( .A(r[5]), .B(sbox_F_q2[0]), .Z(sbox_q2[0]) );
  XOR2_X1 sbox_F_U6 ( .A(r[2]), .B(sbox_F_q1[3]), .Z(sbox_q1[3]) );
  XOR2_X1 sbox_F_U5 ( .A(r[0]), .B(sbox_F_q1[2]), .Z(sbox_q1[2]) );
  XOR2_X1 sbox_F_U4 ( .A(r[6]), .B(sbox_F_q1[1]), .Z(sbox_q1[1]) );
  XOR2_X1 sbox_F_U3 ( .A(r[4]), .B(sbox_F_q1[0]), .Z(sbox_q1[0]) );
  DFF_X1 sbox_F_CF_Reg_reg_0_ ( .D(sbox_F_CF_Out[0]), .CK(clk), .Q(
        sbox_F_CF_Reg[0]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_1_ ( .D(sbox_F_CF_Out[1]), .CK(clk), .Q(
        sbox_F_CF_Reg[1]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_2_ ( .D(sbox_F_CF_Out[2]), .CK(clk), .Q(
        sbox_F_CF_Reg[2]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_3_ ( .D(sbox_F_CF_Out[3]), .CK(clk), .Q(
        sbox_F_CF_Reg[3]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_4_ ( .D(sbox_F_CF_Out[4]), .CK(clk), .Q(
        sbox_F_CF_Reg[4]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_5_ ( .D(sbox_F_CF_Out[5]), .CK(clk), .Q(
        sbox_F_CF_Reg[5]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_6_ ( .D(sbox_F_CF_Out[6]), .CK(clk), .Q(
        sbox_F_CF_Reg[6]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_7_ ( .D(sbox_F_CF_Out[7]), .CK(clk), .Q(
        sbox_F_CF_Reg[7]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_8_ ( .D(sbox_F_CF_Out[8]), .CK(clk), .Q(
        sbox_F_CF_Reg[8]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_9_ ( .D(sbox_F_CF_Out[9]), .CK(clk), .Q(
        sbox_F_CF_Reg[9]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_10_ ( .D(sbox_F_CF_Out[10]), .CK(clk), .Q(
        sbox_F_CF_Reg[10]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_11_ ( .D(sbox_F_CF_Out[11]), .CK(clk), .Q(
        sbox_F_CF_Reg[11]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_12_ ( .D(sbox_F_CF_Out[12]), .CK(clk), .Q(
        sbox_F_CF_Reg[12]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_13_ ( .D(sbox_F_CF_Out[13]), .CK(clk), .Q(
        sbox_F_CF_Reg[13]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_14_ ( .D(sbox_F_CF_Out[14]), .CK(clk), .Q(
        sbox_F_CF_Reg[14]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_15_ ( .D(sbox_F_CF_Out[15]), .CK(clk), .Q(
        sbox_F_CF_Reg[15]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_16_ ( .D(sbox_F_CF_Out[16]), .CK(clk), .Q(
        sbox_F_CF_Reg[16]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_17_ ( .D(sbox_F_CF_Out[17]), .CK(clk), .Q(
        sbox_F_CF_Reg[17]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_18_ ( .D(sbox_F_CF_Out[18]), .CK(clk), .Q(
        sbox_F_CF_Reg[18]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_19_ ( .D(sbox_F_CF_Out[19]), .CK(clk), .Q(
        sbox_F_CF_Reg[19]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_20_ ( .D(sbox_F_CF_Out[20]), .CK(clk), .Q(
        sbox_F_CF_Reg[20]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_21_ ( .D(sbox_F_CF_Out[21]), .CK(clk), .Q(
        sbox_F_CF_Reg[21]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_22_ ( .D(sbox_F_CF_Out[22]), .CK(clk), .Q(
        sbox_F_CF_Reg[22]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_23_ ( .D(sbox_F_CF_Out[23]), .CK(clk), .Q(
        sbox_F_CF_Reg[23]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_24_ ( .D(sbox_F_CF_Out[24]), .CK(clk), .Q(
        sbox_F_CF_Reg[24]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_25_ ( .D(sbox_F_CF_Out[25]), .CK(clk), .Q(
        sbox_F_CF_Reg[25]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_26_ ( .D(sbox_F_CF_Out[26]), .CK(clk), .Q(
        sbox_F_CF_Reg[26]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_27_ ( .D(sbox_F_CF_Out[27]), .CK(clk), .Q(
        sbox_F_CF_Reg[27]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_28_ ( .D(sbox_F_CF_Out[28]), .CK(clk), .Q(
        sbox_F_CF_Reg[28]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_29_ ( .D(sbox_F_CF_Out[29]), .CK(clk), .Q(
        sbox_F_CF_Reg[29]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_30_ ( .D(sbox_F_CF_Out[30]), .CK(clk), .Q(
        sbox_F_CF_Reg[30]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_31_ ( .D(sbox_F_CF_Out[31]), .CK(clk), .Q(
        sbox_F_CF_Reg[31]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_32_ ( .D(sbox_F_CF_Out[32]), .CK(clk), .Q(
        sbox_F_CF_Reg[32]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_33_ ( .D(sbox_F_CF_Out[33]), .CK(clk), .Q(
        sbox_F_CF_Reg[33]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_34_ ( .D(sbox_F_CF_Out[34]), .CK(clk), .Q(
        sbox_F_CF_Reg[34]), .QN() );
  DFF_X1 sbox_F_CF_Reg_reg_35_ ( .D(sbox_F_CF_Out[35]), .CK(clk), .Q(
        sbox_F_CF_Reg[35]), .QN() );
  AND2_X1 sbox_F_Inst_0__CF_Inst_U1 ( .A1(sbox_F_in1_reg[1]), .A2(
        sbox_F_in1_reg[3]), .ZN(sbox_F_CF_Out[0]) );
  XNOR2_X1 sbox_F_Inst_1__CF_Inst_U2 ( .A(sbox_F_Inst_1__CF_Inst_n1), .B(
        sbox_F_in2_reg[2]), .ZN(sbox_F_CF_Out[1]) );
  NAND2_X1 sbox_F_Inst_1__CF_Inst_U1 ( .A1(sbox_F_in2_reg[1]), .A2(
        sbox_F_in1_reg[3]), .ZN(sbox_F_Inst_1__CF_Inst_n1) );
  OR2_X1 sbox_F_Inst_2__CF_Inst_U1 ( .A1(sbox_F_in1_reg[3]), .A2(
        sbox_F_in3_reg[1]), .ZN(sbox_F_CF_Out[2]) );
  XNOR2_X1 sbox_F_Inst_3__CF_Inst_U2 ( .A(sbox_F_Inst_3__CF_Inst_n1), .B(
        sbox_F_in1_reg[2]), .ZN(sbox_F_CF_Out[3]) );
  NAND2_X1 sbox_F_Inst_3__CF_Inst_U1 ( .A1(sbox_F_in1_reg[1]), .A2(
        sbox_F_in2_reg[3]), .ZN(sbox_F_Inst_3__CF_Inst_n1) );
  NOR2_X1 sbox_F_Inst_4__CF_Inst_U2 ( .A1(sbox_F_in2_reg[3]), .A2(
        sbox_F_Inst_4__CF_Inst_n2), .ZN(sbox_F_CF_Out[4]) );
  INV_X1 sbox_F_Inst_4__CF_Inst_U1 ( .A(sbox_F_in2_reg[1]), .ZN(
        sbox_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 sbox_F_Inst_5__CF_Inst_U2 ( .A1(sbox_F_in3_reg[1]), .A2(
        sbox_F_Inst_5__CF_Inst_n2), .ZN(sbox_F_CF_Out[5]) );
  INV_X1 sbox_F_Inst_5__CF_Inst_U1 ( .A(sbox_F_in2_reg[3]), .ZN(
        sbox_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 sbox_F_Inst_6__CF_Inst_U2 ( .A1(sbox_F_in1_reg[1]), .A2(
        sbox_F_Inst_6__CF_Inst_n2), .ZN(sbox_F_CF_Out[6]) );
  INV_X1 sbox_F_Inst_6__CF_Inst_U1 ( .A(sbox_F_in3_reg[3]), .ZN(
        sbox_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 sbox_F_Inst_7__CF_Inst_U2 ( .A1(sbox_F_in3_reg[3]), .A2(
        sbox_F_Inst_7__CF_Inst_n2), .ZN(sbox_F_CF_Out[7]) );
  INV_X1 sbox_F_Inst_7__CF_Inst_U1 ( .A(sbox_F_in2_reg[1]), .ZN(
        sbox_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 sbox_F_Inst_8__CF_Inst_U3 ( .A(sbox_F_in3_reg[2]), .B(
        sbox_F_Inst_8__CF_Inst_n2), .ZN(sbox_F_CF_Out[8]) );
  NAND2_X1 sbox_F_Inst_8__CF_Inst_U2 ( .A1(sbox_F_in3_reg[1]), .A2(
        sbox_F_Inst_8__CF_Inst_n1), .ZN(sbox_F_Inst_8__CF_Inst_n2) );
  INV_X1 sbox_F_Inst_8__CF_Inst_U1 ( .A(sbox_F_in3_reg[3]), .ZN(
        sbox_F_Inst_8__CF_Inst_n1) );
  NOR2_X1 sbox_F_Inst_9__CF_Inst_U2 ( .A1(sbox_F_in1_reg[1]), .A2(
        sbox_F_Inst_9__CF_Inst_n2), .ZN(sbox_F_CF_Out[9]) );
  INV_X1 sbox_F_Inst_9__CF_Inst_U1 ( .A(sbox_F_in1_reg[3]), .ZN(
        sbox_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 sbox_F_Inst_10__CF_Inst_U3 ( .A(sbox_F_in2_reg[2]), .B(
        sbox_F_Inst_10__CF_Inst_n2), .ZN(sbox_F_CF_Out[10]) );
  NAND2_X1 sbox_F_Inst_10__CF_Inst_U2 ( .A1(sbox_F_in1_reg[3]), .A2(
        sbox_F_Inst_10__CF_Inst_n1), .ZN(sbox_F_Inst_10__CF_Inst_n2) );
  INV_X1 sbox_F_Inst_10__CF_Inst_U1 ( .A(sbox_F_in2_reg[1]), .ZN(
        sbox_F_Inst_10__CF_Inst_n1) );
  NOR2_X1 sbox_F_Inst_11__CF_Inst_U2 ( .A1(sbox_F_in1_reg[3]), .A2(
        sbox_F_Inst_11__CF_Inst_n2), .ZN(sbox_F_CF_Out[11]) );
  INV_X1 sbox_F_Inst_11__CF_Inst_U1 ( .A(sbox_F_in3_reg[1]), .ZN(
        sbox_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 sbox_F_Inst_12__CF_Inst_U3 ( .A(sbox_F_in1_reg[2]), .B(
        sbox_F_Inst_12__CF_Inst_n2), .ZN(sbox_F_CF_Out[12]) );
  NAND2_X1 sbox_F_Inst_12__CF_Inst_U2 ( .A1(sbox_F_in2_reg[3]), .A2(
        sbox_F_Inst_12__CF_Inst_n1), .ZN(sbox_F_Inst_12__CF_Inst_n2) );
  INV_X1 sbox_F_Inst_12__CF_Inst_U1 ( .A(sbox_F_in1_reg[1]), .ZN(
        sbox_F_Inst_12__CF_Inst_n1) );
  NOR2_X1 sbox_F_Inst_13__CF_Inst_U2 ( .A1(sbox_F_in2_reg[3]), .A2(
        sbox_F_Inst_13__CF_Inst_n2), .ZN(sbox_F_CF_Out[13]) );
  INV_X1 sbox_F_Inst_13__CF_Inst_U1 ( .A(sbox_F_in2_reg[1]), .ZN(
        sbox_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 sbox_F_Inst_14__CF_Inst_U2 ( .A1(sbox_F_in3_reg[1]), .A2(
        sbox_F_Inst_14__CF_Inst_n2), .ZN(sbox_F_CF_Out[14]) );
  INV_X1 sbox_F_Inst_14__CF_Inst_U1 ( .A(sbox_F_in2_reg[3]), .ZN(
        sbox_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 sbox_F_Inst_15__CF_Inst_U2 ( .A1(sbox_F_in1_reg[1]), .A2(
        sbox_F_Inst_15__CF_Inst_n2), .ZN(sbox_F_CF_Out[15]) );
  INV_X1 sbox_F_Inst_15__CF_Inst_U1 ( .A(sbox_F_in3_reg[3]), .ZN(
        sbox_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 sbox_F_Inst_16__CF_Inst_U2 ( .A1(sbox_F_in3_reg[3]), .A2(
        sbox_F_Inst_16__CF_Inst_n2), .ZN(sbox_F_CF_Out[16]) );
  INV_X1 sbox_F_Inst_16__CF_Inst_U1 ( .A(sbox_F_in2_reg[1]), .ZN(
        sbox_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 sbox_F_Inst_17__CF_Inst_U2 ( .A(sbox_F_Inst_17__CF_Inst_n2), .B(
        sbox_F_in3_reg[2]), .ZN(sbox_F_CF_Out[17]) );
  NOR2_X1 sbox_F_Inst_17__CF_Inst_U1 ( .A1(sbox_F_in3_reg[1]), .A2(
        sbox_F_in3_reg[3]), .ZN(sbox_F_Inst_17__CF_Inst_n2) );
  AOI211_X1 sbox_F_Inst_18__CF_Inst_U2 ( .C1(sbox_F_in1_reg[1]), .C2(
        sbox_F_in1_reg[2]), .A(sbox_F_in1_reg[3]), .B(
        sbox_F_Inst_18__CF_Inst_n1), .ZN(sbox_F_CF_Out[18]) );
  NOR2_X1 sbox_F_Inst_18__CF_Inst_U1 ( .A1(sbox_F_in1_reg[1]), .A2(
        sbox_F_in1_reg[2]), .ZN(sbox_F_Inst_18__CF_Inst_n1) );
  AOI21_X1 sbox_F_Inst_19__CF_Inst_U3 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_Inst_19__CF_Inst_n2), .A(sbox_F_Inst_19__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[19]) );
  OAI21_X1 sbox_F_Inst_19__CF_Inst_U2 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_Inst_19__CF_Inst_n2), .A(sbox_F_in1_reg[3]), .ZN(
        sbox_F_Inst_19__CF_Inst_n1) );
  INV_X1 sbox_F_Inst_19__CF_Inst_U1 ( .A(sbox_F_in2_reg[2]), .ZN(
        sbox_F_Inst_19__CF_Inst_n2) );
  OAI21_X1 sbox_F_Inst_20__CF_Inst_U3 ( .B1(sbox_F_Inst_20__CF_Inst_n2), .B2(
        sbox_F_in3_reg[1]), .A(sbox_F_Inst_20__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[20]) );
  NAND2_X1 sbox_F_Inst_20__CF_Inst_U2 ( .A1(sbox_F_Inst_20__CF_Inst_n2), .A2(
        sbox_F_in3_reg[2]), .ZN(sbox_F_Inst_20__CF_Inst_n1) );
  INV_X1 sbox_F_Inst_20__CF_Inst_U1 ( .A(sbox_F_in1_reg[3]), .ZN(
        sbox_F_Inst_20__CF_Inst_n2) );
  MUX2_X1 sbox_F_Inst_21__CF_Inst_U1 ( .A(sbox_F_in1_reg[1]), .B(
        sbox_F_in1_reg[2]), .S(sbox_F_in2_reg[3]), .Z(sbox_F_CF_Out[21]) );
  AOI21_X1 sbox_F_Inst_22__CF_Inst_U2 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_in2_reg[2]), .A(sbox_F_Inst_22__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[22]) );
  OAI21_X1 sbox_F_Inst_22__CF_Inst_U1 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_in2_reg[2]), .A(sbox_F_in2_reg[3]), .ZN(
        sbox_F_Inst_22__CF_Inst_n1) );
  AOI211_X1 sbox_F_Inst_23__CF_Inst_U2 ( .C1(sbox_F_in3_reg[1]), .C2(
        sbox_F_in3_reg[2]), .A(sbox_F_in2_reg[3]), .B(
        sbox_F_Inst_23__CF_Inst_n1), .ZN(sbox_F_CF_Out[23]) );
  NOR2_X1 sbox_F_Inst_23__CF_Inst_U1 ( .A1(sbox_F_in3_reg[1]), .A2(
        sbox_F_in3_reg[2]), .ZN(sbox_F_Inst_23__CF_Inst_n1) );
  AOI211_X1 sbox_F_Inst_24__CF_Inst_U2 ( .C1(sbox_F_in1_reg[1]), .C2(
        sbox_F_in1_reg[2]), .A(sbox_F_in3_reg[3]), .B(
        sbox_F_Inst_24__CF_Inst_n1), .ZN(sbox_F_CF_Out[24]) );
  NOR2_X1 sbox_F_Inst_24__CF_Inst_U1 ( .A1(sbox_F_in1_reg[1]), .A2(
        sbox_F_in1_reg[2]), .ZN(sbox_F_Inst_24__CF_Inst_n1) );
  MUX2_X1 sbox_F_Inst_25__CF_Inst_U1 ( .A(sbox_F_in2_reg[1]), .B(
        sbox_F_in2_reg[2]), .S(sbox_F_in3_reg[3]), .Z(sbox_F_CF_Out[25]) );
  AOI21_X1 sbox_F_Inst_26__CF_Inst_U2 ( .B1(sbox_F_in3_reg[1]), .B2(
        sbox_F_in3_reg[2]), .A(sbox_F_Inst_26__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[26]) );
  OAI21_X1 sbox_F_Inst_26__CF_Inst_U1 ( .B1(sbox_F_in3_reg[1]), .B2(
        sbox_F_in3_reg[2]), .A(sbox_F_in3_reg[3]), .ZN(
        sbox_F_Inst_26__CF_Inst_n1) );
  XNOR2_X1 sbox_F_Inst_27__CF_Inst_U3 ( .A(sbox_F_in1_reg[0]), .B(
        sbox_F_Inst_27__CF_Inst_n3), .ZN(sbox_F_CF_Out[27]) );
  OAI21_X1 sbox_F_Inst_27__CF_Inst_U2 ( .B1(sbox_F_in1_reg[1]), .B2(
        sbox_F_in1_reg[2]), .A(sbox_F_Inst_27__CF_Inst_n2), .ZN(
        sbox_F_Inst_27__CF_Inst_n3) );
  AOI21_X1 sbox_F_Inst_27__CF_Inst_U1 ( .B1(sbox_F_in1_reg[1]), .B2(
        sbox_F_in1_reg[2]), .A(sbox_F_in1_reg[3]), .ZN(
        sbox_F_Inst_27__CF_Inst_n2) );
  AOI21_X1 sbox_F_Inst_28__CF_Inst_U3 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_Inst_28__CF_Inst_n2), .A(sbox_F_Inst_28__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[28]) );
  OAI21_X1 sbox_F_Inst_28__CF_Inst_U2 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_Inst_28__CF_Inst_n2), .A(sbox_F_in1_reg[3]), .ZN(
        sbox_F_Inst_28__CF_Inst_n1) );
  INV_X1 sbox_F_Inst_28__CF_Inst_U1 ( .A(sbox_F_in2_reg[2]), .ZN(
        sbox_F_Inst_28__CF_Inst_n2) );
  OAI21_X1 sbox_F_Inst_29__CF_Inst_U3 ( .B1(sbox_F_Inst_29__CF_Inst_n2), .B2(
        sbox_F_in3_reg[1]), .A(sbox_F_Inst_29__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[29]) );
  NAND2_X1 sbox_F_Inst_29__CF_Inst_U2 ( .A1(sbox_F_Inst_29__CF_Inst_n2), .A2(
        sbox_F_in3_reg[2]), .ZN(sbox_F_Inst_29__CF_Inst_n1) );
  INV_X1 sbox_F_Inst_29__CF_Inst_U1 ( .A(sbox_F_in1_reg[3]), .ZN(
        sbox_F_Inst_29__CF_Inst_n2) );
  XNOR2_X1 sbox_F_Inst_30__CF_Inst_U3 ( .A(sbox_F_in2_reg[0]), .B(
        sbox_F_Inst_30__CF_Inst_n2), .ZN(sbox_F_CF_Out[30]) );
  AOI22_X1 sbox_F_Inst_30__CF_Inst_U2 ( .A1(sbox_F_in2_reg[3]), .A2(
        sbox_F_in1_reg[2]), .B1(sbox_F_in1_reg[1]), .B2(
        sbox_F_Inst_30__CF_Inst_n1), .ZN(sbox_F_Inst_30__CF_Inst_n2) );
  INV_X1 sbox_F_Inst_30__CF_Inst_U1 ( .A(sbox_F_in2_reg[3]), .ZN(
        sbox_F_Inst_30__CF_Inst_n1) );
  AOI21_X1 sbox_F_Inst_31__CF_Inst_U2 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_in2_reg[2]), .A(sbox_F_Inst_31__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[31]) );
  OAI21_X1 sbox_F_Inst_31__CF_Inst_U1 ( .B1(sbox_F_in2_reg[1]), .B2(
        sbox_F_in2_reg[2]), .A(sbox_F_in2_reg[3]), .ZN(
        sbox_F_Inst_31__CF_Inst_n1) );
  AOI211_X1 sbox_F_Inst_32__CF_Inst_U2 ( .C1(sbox_F_in3_reg[1]), .C2(
        sbox_F_in3_reg[2]), .A(sbox_F_in2_reg[3]), .B(
        sbox_F_Inst_32__CF_Inst_n1), .ZN(sbox_F_CF_Out[32]) );
  NOR2_X1 sbox_F_Inst_32__CF_Inst_U1 ( .A1(sbox_F_in3_reg[1]), .A2(
        sbox_F_in3_reg[2]), .ZN(sbox_F_Inst_32__CF_Inst_n1) );
  XNOR2_X1 sbox_F_Inst_33__CF_Inst_U4 ( .A(sbox_F_in3_reg[0]), .B(
        sbox_F_Inst_33__CF_Inst_n5), .ZN(sbox_F_CF_Out[33]) );
  AOI221_X1 sbox_F_Inst_33__CF_Inst_U3 ( .B1(sbox_F_in1_reg[1]), .B2(
        sbox_F_Inst_33__CF_Inst_n4), .C1(sbox_F_Inst_33__CF_Inst_n3), .C2(
        sbox_F_in1_reg[2]), .A(sbox_F_in3_reg[3]), .ZN(
        sbox_F_Inst_33__CF_Inst_n5) );
  INV_X1 sbox_F_Inst_33__CF_Inst_U2 ( .A(sbox_F_in1_reg[1]), .ZN(
        sbox_F_Inst_33__CF_Inst_n3) );
  INV_X1 sbox_F_Inst_33__CF_Inst_U1 ( .A(sbox_F_in1_reg[2]), .ZN(
        sbox_F_Inst_33__CF_Inst_n4) );
  MUX2_X1 sbox_F_Inst_34__CF_Inst_U1 ( .A(sbox_F_in2_reg[1]), .B(
        sbox_F_in2_reg[2]), .S(sbox_F_in3_reg[3]), .Z(sbox_F_CF_Out[34]) );
  AOI21_X1 sbox_F_Inst_35__CF_Inst_U3 ( .B1(sbox_F_in3_reg[1]), .B2(
        sbox_F_Inst_35__CF_Inst_n2), .A(sbox_F_Inst_35__CF_Inst_n1), .ZN(
        sbox_F_CF_Out[35]) );
  OAI21_X1 sbox_F_Inst_35__CF_Inst_U2 ( .B1(sbox_F_in3_reg[1]), .B2(
        sbox_F_Inst_35__CF_Inst_n2), .A(sbox_F_in3_reg[3]), .ZN(
        sbox_F_Inst_35__CF_Inst_n1) );
  INV_X1 sbox_F_Inst_35__CF_Inst_U1 ( .A(sbox_F_in3_reg[2]), .ZN(
        sbox_F_Inst_35__CF_Inst_n2) );
  XNOR2_X1 sbox_F_InstXOR_0__Compression1_U2 ( .A(
        sbox_F_InstXOR_0__Compression1_n3), .B(sbox_F_CF_Reg[2]), .ZN(
        sbox_F_q1[0]) );
  XNOR2_X1 sbox_F_InstXOR_0__Compression1_U1 ( .A(sbox_F_CF_Reg[0]), .B(
        sbox_F_CF_Reg[1]), .ZN(sbox_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 sbox_F_InstXOR_0__Compression2_U2 ( .A(
        sbox_F_InstXOR_0__Compression2_n3), .B(sbox_F_CF_Reg[5]), .ZN(
        sbox_F_q2[0]) );
  XNOR2_X1 sbox_F_InstXOR_0__Compression2_U1 ( .A(sbox_F_CF_Reg[3]), .B(
        sbox_F_CF_Reg[4]), .ZN(sbox_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 sbox_F_InstXOR_0__Compression3_U2 ( .A(
        sbox_F_InstXOR_0__Compression3_n3), .B(sbox_F_CF_Reg[8]), .ZN(
        sbox_F_q3[0]) );
  XNOR2_X1 sbox_F_InstXOR_0__Compression3_U1 ( .A(sbox_F_CF_Reg[6]), .B(
        sbox_F_CF_Reg[7]), .ZN(sbox_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 sbox_F_InstXOR_1__Compression1_U2 ( .A(
        sbox_F_InstXOR_1__Compression1_n3), .B(sbox_F_CF_Reg[11]), .ZN(
        sbox_F_q1[1]) );
  XNOR2_X1 sbox_F_InstXOR_1__Compression1_U1 ( .A(sbox_F_CF_Reg[9]), .B(
        sbox_F_CF_Reg[10]), .ZN(sbox_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 sbox_F_InstXOR_1__Compression2_U2 ( .A(
        sbox_F_InstXOR_1__Compression2_n3), .B(sbox_F_CF_Reg[14]), .ZN(
        sbox_F_q2[1]) );
  XNOR2_X1 sbox_F_InstXOR_1__Compression2_U1 ( .A(sbox_F_CF_Reg[12]), .B(
        sbox_F_CF_Reg[13]), .ZN(sbox_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 sbox_F_InstXOR_1__Compression3_U2 ( .A(
        sbox_F_InstXOR_1__Compression3_n3), .B(sbox_F_CF_Reg[17]), .ZN(
        sbox_F_q3[1]) );
  XNOR2_X1 sbox_F_InstXOR_1__Compression3_U1 ( .A(sbox_F_CF_Reg[15]), .B(
        sbox_F_CF_Reg[16]), .ZN(sbox_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 sbox_F_InstXOR_2__Compression1_U2 ( .A(
        sbox_F_InstXOR_2__Compression1_n3), .B(sbox_F_CF_Reg[20]), .ZN(
        sbox_F_q1[2]) );
  XNOR2_X1 sbox_F_InstXOR_2__Compression1_U1 ( .A(sbox_F_CF_Reg[18]), .B(
        sbox_F_CF_Reg[19]), .ZN(sbox_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 sbox_F_InstXOR_2__Compression2_U2 ( .A(
        sbox_F_InstXOR_2__Compression2_n3), .B(sbox_F_CF_Reg[23]), .ZN(
        sbox_F_q2[2]) );
  XNOR2_X1 sbox_F_InstXOR_2__Compression2_U1 ( .A(sbox_F_CF_Reg[21]), .B(
        sbox_F_CF_Reg[22]), .ZN(sbox_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 sbox_F_InstXOR_2__Compression3_U2 ( .A(
        sbox_F_InstXOR_2__Compression3_n3), .B(sbox_F_CF_Reg[26]), .ZN(
        sbox_F_q3[2]) );
  XNOR2_X1 sbox_F_InstXOR_2__Compression3_U1 ( .A(sbox_F_CF_Reg[24]), .B(
        sbox_F_CF_Reg[25]), .ZN(sbox_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 sbox_F_InstXOR_3__Compression1_U2 ( .A(
        sbox_F_InstXOR_3__Compression1_n3), .B(sbox_F_CF_Reg[29]), .ZN(
        sbox_F_q1[3]) );
  XNOR2_X1 sbox_F_InstXOR_3__Compression1_U1 ( .A(sbox_F_CF_Reg[27]), .B(
        sbox_F_CF_Reg[28]), .ZN(sbox_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 sbox_F_InstXOR_3__Compression2_U2 ( .A(
        sbox_F_InstXOR_3__Compression2_n3), .B(sbox_F_CF_Reg[32]), .ZN(
        sbox_F_q2[3]) );
  XNOR2_X1 sbox_F_InstXOR_3__Compression2_U1 ( .A(sbox_F_CF_Reg[30]), .B(
        sbox_F_CF_Reg[31]), .ZN(sbox_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 sbox_F_InstXOR_3__Compression3_U2 ( .A(
        sbox_F_InstXOR_3__Compression3_n3), .B(sbox_F_CF_Reg[35]), .ZN(
        sbox_F_q3[3]) );
  XNOR2_X1 sbox_F_InstXOR_3__Compression3_U1 ( .A(sbox_F_CF_Reg[33]), .B(
        sbox_F_CF_Reg[34]), .ZN(sbox_F_InstXOR_3__Compression3_n3) );
  XOR2_X1 sbox_G_U5 ( .A(sbox_Rq2[3]), .B(sbox_Rq2[0]), .Z(sbox_G_N2) );
  XOR2_X1 sbox_G_U4 ( .A(sbox_Rq3[3]), .B(sbox_Rq3[0]), .Z(sbox_G_N3) );
  XNOR2_X1 sbox_G_U3 ( .A(sbox_Rq1[3]), .B(sbox_Rq1[0]), .ZN(sbox_G_n1) );
  DFF_X1 sbox_G_out1_reg_0_ ( .D(sbox_G_n1), .CK(clk), .Q(sboxOut1[0]), .QN()
         );
  DFF_X1 sbox_G_CF_Reg_reg_0_ ( .D(sbox_G_CF_Out[0]), .CK(clk), .Q(
        sbox_G_CF_Reg[0]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_1_ ( .D(sbox_G_CF_Out[1]), .CK(clk), .Q(
        sbox_G_CF_Reg[1]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_2_ ( .D(sbox_G_CF_Out[2]), .CK(clk), .Q(
        sbox_G_CF_Reg[2]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_3_ ( .D(sbox_G_CF_Out[3]), .CK(clk), .Q(
        sbox_G_CF_Reg[3]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_4_ ( .D(sbox_G_CF_Out[4]), .CK(clk), .Q(
        sbox_G_CF_Reg[4]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_5_ ( .D(sbox_G_CF_Out[5]), .CK(clk), .Q(
        sbox_G_CF_Reg[5]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_6_ ( .D(sbox_G_CF_Out[6]), .CK(clk), .Q(
        sbox_G_CF_Reg[6]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_7_ ( .D(sbox_G_CF_Out[7]), .CK(clk), .Q(
        sbox_G_CF_Reg[7]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_8_ ( .D(sbox_G_CF_Out[8]), .CK(clk), .Q(
        sbox_G_CF_Reg[8]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_9_ ( .D(sbox_G_CF_Out[9]), .CK(clk), .Q(
        sbox_G_CF_Reg[9]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_10_ ( .D(sbox_G_CF_Out[10]), .CK(clk), .Q(
        sbox_G_CF_Reg[10]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_11_ ( .D(sbox_G_CF_Out[11]), .CK(clk), .Q(
        sbox_G_CF_Reg[11]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_12_ ( .D(sbox_G_CF_Out[12]), .CK(clk), .Q(
        sbox_G_CF_Reg[12]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_13_ ( .D(sbox_G_CF_Out[13]), .CK(clk), .Q(
        sbox_G_CF_Reg[13]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_14_ ( .D(sbox_G_CF_Out[14]), .CK(clk), .Q(
        sbox_G_CF_Reg[14]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_15_ ( .D(sbox_G_CF_Out[15]), .CK(clk), .Q(
        sbox_G_CF_Reg[15]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_16_ ( .D(sbox_G_CF_Out[16]), .CK(clk), .Q(
        sbox_G_CF_Reg[16]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_17_ ( .D(sbox_G_CF_Out[17]), .CK(clk), .Q(
        sbox_G_CF_Reg[17]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_18_ ( .D(sbox_G_CF_Out[18]), .CK(clk), .Q(
        sbox_G_CF_Reg[18]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_19_ ( .D(sbox_G_CF_Out[19]), .CK(clk), .Q(
        sbox_G_CF_Reg[19]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_20_ ( .D(sbox_G_CF_Out[20]), .CK(clk), .Q(
        sbox_G_CF_Reg[20]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_21_ ( .D(sbox_G_CF_Out[21]), .CK(clk), .Q(
        sbox_G_CF_Reg[21]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_22_ ( .D(sbox_G_CF_Out[22]), .CK(clk), .Q(
        sbox_G_CF_Reg[22]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_23_ ( .D(sbox_G_CF_Out[23]), .CK(clk), .Q(
        sbox_G_CF_Reg[23]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_24_ ( .D(sbox_G_CF_Out[24]), .CK(clk), .Q(
        sbox_G_CF_Reg[24]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_25_ ( .D(sbox_G_CF_Out[25]), .CK(clk), .Q(
        sbox_G_CF_Reg[25]), .QN() );
  DFF_X1 sbox_G_CF_Reg_reg_26_ ( .D(sbox_G_CF_Out[26]), .CK(clk), .Q(
        sbox_G_CF_Reg[26]), .QN() );
  DFF_X1 sbox_G_out3_reg_0_ ( .D(sbox_G_N3), .CK(clk), .Q(sboxOut3[0]), .QN()
         );
  DFF_X1 sbox_G_out2_reg_0_ ( .D(sbox_G_N2), .CK(clk), .Q(sboxOut2[0]), .QN()
         );
  AND2_X1 sbox_G_Inst_0__CF_Inst_U1 ( .A1(sbox_Rq1[2]), .A2(sbox_Rq1[3]), .ZN(
        sbox_G_CF_Out[0]) );
  NOR2_X1 sbox_G_Inst_1__CF_Inst_U2 ( .A1(sbox_Rq1[3]), .A2(
        sbox_G_Inst_1__CF_Inst_n2), .ZN(sbox_G_CF_Out[1]) );
  INV_X1 sbox_G_Inst_1__CF_Inst_U1 ( .A(sbox_Rq2[2]), .ZN(
        sbox_G_Inst_1__CF_Inst_n2) );
  XNOR2_X1 sbox_G_Inst_2__CF_Inst_U3 ( .A(sbox_Rq1[1]), .B(
        sbox_G_Inst_2__CF_Inst_n2), .ZN(sbox_G_CF_Out[2]) );
  NAND2_X1 sbox_G_Inst_2__CF_Inst_U2 ( .A1(sbox_Rq3[2]), .A2(
        sbox_G_Inst_2__CF_Inst_n1), .ZN(sbox_G_Inst_2__CF_Inst_n2) );
  INV_X1 sbox_G_Inst_2__CF_Inst_U1 ( .A(sbox_Rq1[3]), .ZN(
        sbox_G_Inst_2__CF_Inst_n1) );
  NOR2_X1 sbox_G_Inst_3__CF_Inst_U2 ( .A1(sbox_Rq2[3]), .A2(
        sbox_G_Inst_3__CF_Inst_n2), .ZN(sbox_G_CF_Out[3]) );
  INV_X1 sbox_G_Inst_3__CF_Inst_U1 ( .A(sbox_Rq1[2]), .ZN(
        sbox_G_Inst_3__CF_Inst_n2) );
  AND2_X1 sbox_G_Inst_4__CF_Inst_U1 ( .A1(sbox_Rq2[2]), .A2(sbox_Rq2[3]), .ZN(
        sbox_G_CF_Out[4]) );
  XNOR2_X1 sbox_G_Inst_5__CF_Inst_U3 ( .A(sbox_Rq2[1]), .B(
        sbox_G_Inst_5__CF_Inst_n2), .ZN(sbox_G_CF_Out[5]) );
  NAND2_X1 sbox_G_Inst_5__CF_Inst_U2 ( .A1(sbox_Rq3[2]), .A2(
        sbox_G_Inst_5__CF_Inst_n1), .ZN(sbox_G_Inst_5__CF_Inst_n2) );
  INV_X1 sbox_G_Inst_5__CF_Inst_U1 ( .A(sbox_Rq2[3]), .ZN(
        sbox_G_Inst_5__CF_Inst_n1) );
  XNOR2_X1 sbox_G_Inst_6__CF_Inst_U2 ( .A(sbox_G_Inst_6__CF_Inst_n1), .B(
        sbox_Rq3[1]), .ZN(sbox_G_CF_Out[6]) );
  NAND2_X1 sbox_G_Inst_6__CF_Inst_U1 ( .A1(sbox_Rq1[2]), .A2(sbox_Rq3[3]), 
        .ZN(sbox_G_Inst_6__CF_Inst_n1) );
  AND2_X1 sbox_G_Inst_7__CF_Inst_U1 ( .A1(sbox_Rq2[2]), .A2(sbox_Rq3[3]), .ZN(
        sbox_G_CF_Out[7]) );
  NOR2_X1 sbox_G_Inst_8__CF_Inst_U2 ( .A1(sbox_Rq3[3]), .A2(
        sbox_G_Inst_8__CF_Inst_n2), .ZN(sbox_G_CF_Out[8]) );
  INV_X1 sbox_G_Inst_8__CF_Inst_U1 ( .A(sbox_Rq3[2]), .ZN(
        sbox_G_Inst_8__CF_Inst_n2) );
  XNOR2_X1 sbox_G_Inst_9__CF_Inst_U3 ( .A(sbox_Rq1[0]), .B(
        sbox_G_Inst_9__CF_Inst_n2), .ZN(sbox_G_CF_Out[9]) );
  NAND2_X1 sbox_G_Inst_9__CF_Inst_U2 ( .A1(sbox_Rq1[1]), .A2(
        sbox_G_Inst_9__CF_Inst_n1), .ZN(sbox_G_Inst_9__CF_Inst_n2) );
  INV_X1 sbox_G_Inst_9__CF_Inst_U1 ( .A(sbox_Rq1[3]), .ZN(
        sbox_G_Inst_9__CF_Inst_n1) );
  AND2_X1 sbox_G_Inst_10__CF_Inst_U1 ( .A1(sbox_Rq2[1]), .A2(sbox_Rq1[3]), 
        .ZN(sbox_G_CF_Out[10]) );
  XNOR2_X1 sbox_G_Inst_11__CF_Inst_U3 ( .A(sbox_Rq1[2]), .B(
        sbox_G_Inst_11__CF_Inst_n2), .ZN(sbox_G_CF_Out[11]) );
  NAND2_X1 sbox_G_Inst_11__CF_Inst_U2 ( .A1(sbox_Rq3[1]), .A2(
        sbox_G_Inst_11__CF_Inst_n1), .ZN(sbox_G_Inst_11__CF_Inst_n2) );
  INV_X1 sbox_G_Inst_11__CF_Inst_U1 ( .A(sbox_Rq1[3]), .ZN(
        sbox_G_Inst_11__CF_Inst_n1) );
  XNOR2_X1 sbox_G_Inst_12__CF_Inst_U3 ( .A(sbox_Rq2[0]), .B(
        sbox_G_Inst_12__CF_Inst_n2), .ZN(sbox_G_CF_Out[12]) );
  NAND2_X1 sbox_G_Inst_12__CF_Inst_U2 ( .A1(sbox_Rq1[1]), .A2(
        sbox_G_Inst_12__CF_Inst_n1), .ZN(sbox_G_Inst_12__CF_Inst_n2) );
  INV_X1 sbox_G_Inst_12__CF_Inst_U1 ( .A(sbox_Rq2[3]), .ZN(
        sbox_G_Inst_12__CF_Inst_n1) );
  AND2_X1 sbox_G_Inst_13__CF_Inst_U1 ( .A1(sbox_Rq2[1]), .A2(sbox_Rq2[3]), 
        .ZN(sbox_G_CF_Out[13]) );
  XNOR2_X1 sbox_G_Inst_14__CF_Inst_U2 ( .A(sbox_G_Inst_14__CF_Inst_n1), .B(
        sbox_Rq2[2]), .ZN(sbox_G_CF_Out[14]) );
  NAND2_X1 sbox_G_Inst_14__CF_Inst_U1 ( .A1(sbox_Rq3[1]), .A2(sbox_Rq2[3]), 
        .ZN(sbox_G_Inst_14__CF_Inst_n1) );
  XNOR2_X1 sbox_G_Inst_15__CF_Inst_U3 ( .A(sbox_G_Inst_15__CF_Inst_n2), .B(
        sbox_G_Inst_15__CF_Inst_n1), .ZN(sbox_G_CF_Out[15]) );
  NAND2_X1 sbox_G_Inst_15__CF_Inst_U2 ( .A1(sbox_Rq1[1]), .A2(sbox_Rq3[3]), 
        .ZN(sbox_G_Inst_15__CF_Inst_n1) );
  XOR2_X1 sbox_G_Inst_15__CF_Inst_U1 ( .A(sbox_Rq3[0]), .B(sbox_Rq3[2]), .Z(
        sbox_G_Inst_15__CF_Inst_n2) );
  AND2_X1 sbox_G_Inst_16__CF_Inst_U1 ( .A1(sbox_Rq2[1]), .A2(sbox_Rq3[3]), 
        .ZN(sbox_G_CF_Out[16]) );
  NOR2_X1 sbox_G_Inst_17__CF_Inst_U2 ( .A1(sbox_Rq3[3]), .A2(
        sbox_G_Inst_17__CF_Inst_n2), .ZN(sbox_G_CF_Out[17]) );
  INV_X1 sbox_G_Inst_17__CF_Inst_U1 ( .A(sbox_Rq3[1]), .ZN(
        sbox_G_Inst_17__CF_Inst_n2) );
  NAND2_X1 sbox_G_Inst_18__CF_Inst_U2 ( .A1(sbox_Rq1[3]), .A2(
        sbox_G_Inst_18__CF_Inst_n2), .ZN(sbox_G_CF_Out[18]) );
  INV_X1 sbox_G_Inst_18__CF_Inst_U1 ( .A(sbox_Rq1[2]), .ZN(
        sbox_G_Inst_18__CF_Inst_n2) );
  NOR2_X1 sbox_G_Inst_19__CF_Inst_U2 ( .A1(sbox_Rq1[3]), .A2(
        sbox_G_Inst_19__CF_Inst_n2), .ZN(sbox_G_CF_Out[19]) );
  INV_X1 sbox_G_Inst_19__CF_Inst_U1 ( .A(sbox_Rq2[2]), .ZN(
        sbox_G_Inst_19__CF_Inst_n2) );
  XNOR2_X1 sbox_G_Inst_20__CF_Inst_U3 ( .A(sbox_Rq1[1]), .B(
        sbox_G_Inst_20__CF_Inst_n2), .ZN(sbox_G_CF_Out[20]) );
  NAND2_X1 sbox_G_Inst_20__CF_Inst_U2 ( .A1(sbox_Rq3[2]), .A2(
        sbox_G_Inst_20__CF_Inst_n1), .ZN(sbox_G_Inst_20__CF_Inst_n2) );
  INV_X1 sbox_G_Inst_20__CF_Inst_U1 ( .A(sbox_Rq1[3]), .ZN(
        sbox_G_Inst_20__CF_Inst_n1) );
  OR2_X1 sbox_G_Inst_21__CF_Inst_U1 ( .A1(sbox_Rq2[3]), .A2(sbox_Rq1[2]), .ZN(
        sbox_G_CF_Out[21]) );
  AND2_X1 sbox_G_Inst_22__CF_Inst_U1 ( .A1(sbox_Rq2[2]), .A2(sbox_Rq2[3]), 
        .ZN(sbox_G_CF_Out[22]) );
  XNOR2_X1 sbox_G_Inst_23__CF_Inst_U3 ( .A(sbox_Rq2[1]), .B(
        sbox_G_Inst_23__CF_Inst_n2), .ZN(sbox_G_CF_Out[23]) );
  NAND2_X1 sbox_G_Inst_23__CF_Inst_U2 ( .A1(sbox_Rq3[2]), .A2(
        sbox_G_Inst_23__CF_Inst_n1), .ZN(sbox_G_Inst_23__CF_Inst_n2) );
  INV_X1 sbox_G_Inst_23__CF_Inst_U1 ( .A(sbox_Rq2[3]), .ZN(
        sbox_G_Inst_23__CF_Inst_n1) );
  XNOR2_X1 sbox_G_Inst_24__CF_Inst_U2 ( .A(sbox_G_Inst_24__CF_Inst_n1), .B(
        sbox_Rq3[1]), .ZN(sbox_G_CF_Out[24]) );
  NAND2_X1 sbox_G_Inst_24__CF_Inst_U1 ( .A1(sbox_Rq1[2]), .A2(sbox_Rq3[3]), 
        .ZN(sbox_G_Inst_24__CF_Inst_n1) );
  AND2_X1 sbox_G_Inst_25__CF_Inst_U1 ( .A1(sbox_Rq2[2]), .A2(sbox_Rq3[3]), 
        .ZN(sbox_G_CF_Out[25]) );
  OR2_X1 sbox_G_Inst_26__CF_Inst_U1 ( .A1(sbox_Rq3[3]), .A2(sbox_Rq3[2]), .ZN(
        sbox_G_CF_Out[26]) );
  XNOR2_X1 sbox_G_InstXOR_0__Compression1_U2 ( .A(
        sbox_G_InstXOR_0__Compression1_n3), .B(sbox_G_CF_Reg[2]), .ZN(
        sboxOut1[1]) );
  XNOR2_X1 sbox_G_InstXOR_0__Compression1_U1 ( .A(sbox_G_CF_Reg[0]), .B(
        sbox_G_CF_Reg[1]), .ZN(sbox_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 sbox_G_InstXOR_0__Compression2_U2 ( .A(
        sbox_G_InstXOR_0__Compression2_n3), .B(sbox_G_CF_Reg[5]), .ZN(
        sboxOut2[1]) );
  XNOR2_X1 sbox_G_InstXOR_0__Compression2_U1 ( .A(sbox_G_CF_Reg[3]), .B(
        sbox_G_CF_Reg[4]), .ZN(sbox_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 sbox_G_InstXOR_0__Compression3_U2 ( .A(
        sbox_G_InstXOR_0__Compression3_n3), .B(sbox_G_CF_Reg[8]), .ZN(
        sboxOut3[1]) );
  XNOR2_X1 sbox_G_InstXOR_0__Compression3_U1 ( .A(sbox_G_CF_Reg[6]), .B(
        sbox_G_CF_Reg[7]), .ZN(sbox_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 sbox_G_InstXOR_1__Compression1_U2 ( .A(
        sbox_G_InstXOR_1__Compression1_n3), .B(sbox_G_CF_Reg[11]), .ZN(
        sboxOut1[2]) );
  XNOR2_X1 sbox_G_InstXOR_1__Compression1_U1 ( .A(sbox_G_CF_Reg[9]), .B(
        sbox_G_CF_Reg[10]), .ZN(sbox_G_InstXOR_1__Compression1_n3) );
  XNOR2_X1 sbox_G_InstXOR_1__Compression2_U2 ( .A(
        sbox_G_InstXOR_1__Compression2_n3), .B(sbox_G_CF_Reg[14]), .ZN(
        sboxOut2[2]) );
  XNOR2_X1 sbox_G_InstXOR_1__Compression2_U1 ( .A(sbox_G_CF_Reg[12]), .B(
        sbox_G_CF_Reg[13]), .ZN(sbox_G_InstXOR_1__Compression2_n3) );
  XNOR2_X1 sbox_G_InstXOR_1__Compression3_U2 ( .A(
        sbox_G_InstXOR_1__Compression3_n3), .B(sbox_G_CF_Reg[17]), .ZN(
        sboxOut3[2]) );
  XNOR2_X1 sbox_G_InstXOR_1__Compression3_U1 ( .A(sbox_G_CF_Reg[15]), .B(
        sbox_G_CF_Reg[16]), .ZN(sbox_G_InstXOR_1__Compression3_n3) );
  XNOR2_X1 sbox_G_InstXOR_2__Compression1_U2 ( .A(
        sbox_G_InstXOR_2__Compression1_n3), .B(sbox_G_CF_Reg[20]), .ZN(
        sboxOut1[3]) );
  XNOR2_X1 sbox_G_InstXOR_2__Compression1_U1 ( .A(sbox_G_CF_Reg[18]), .B(
        sbox_G_CF_Reg[19]), .ZN(sbox_G_InstXOR_2__Compression1_n3) );
  XNOR2_X1 sbox_G_InstXOR_2__Compression2_U2 ( .A(
        sbox_G_InstXOR_2__Compression2_n3), .B(sbox_G_CF_Reg[23]), .ZN(
        sboxOut2[3]) );
  XNOR2_X1 sbox_G_InstXOR_2__Compression2_U1 ( .A(sbox_G_CF_Reg[21]), .B(
        sbox_G_CF_Reg[22]), .ZN(sbox_G_InstXOR_2__Compression2_n3) );
  XNOR2_X1 sbox_G_InstXOR_2__Compression3_U2 ( .A(
        sbox_G_InstXOR_2__Compression3_n3), .B(sbox_G_CF_Reg[26]), .ZN(
        sboxOut3[3]) );
  XNOR2_X1 sbox_G_InstXOR_2__Compression3_U1 ( .A(sbox_G_CF_Reg[24]), .B(
        sbox_G_CF_Reg[25]), .ZN(sbox_G_InstXOR_2__Compression3_n3) );
endmodule


