
module circuit ( ClkxCI, RstxBI, PTxDI, KxDI, Zmul1xDI, Zmul2xDI, Zmul3xDI, 
        Zinv1xDI, Zinv2xDI, Zinv3xDI, 
        StartxSI, DonexSO, CxDO );
  input [15:0] PTxDI;
  input [15:0] KxDI;
  input [3:0] Zmul1xDI;
  input [3:0] Zmul2xDI;
  input [3:0] Zmul3xDI;
  input [1:0] Zinv1xDI;
  input [1:0] Zinv2xDI;
  input [1:0] Zinv3xDI;
  output [15:0] CxDO;
  input ClkxCI, RstxBI, StartxSI;
  output DonexSO;
  wire   disableKeyRegsxS, ClkKeyRegxC, StateKEYSCHEDULExS, nextRCONxS,
         showRCONxS, FinishedxS, StateKEYADDITION1o3xS, LastRoundxS,
         doMixColumnsxS, n113, n114, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         aes_ctrl_lsfr_23_cycles_1_n24, aes_ctrl_lsfr_23_cycles_1_n23,
         aes_ctrl_lsfr_23_cycles_1_n22, aes_ctrl_lsfr_23_cycles_1_n21,
         aes_ctrl_lsfr_23_cycles_1_n20, aes_ctrl_lsfr_23_cycles_1_n19,
         aes_ctrl_lsfr_23_cycles_1_n18, aes_ctrl_lsfr_23_cycles_1_n17,
         aes_ctrl_lsfr_23_cycles_1_n16, aes_ctrl_lsfr_23_cycles_1_n15,
         aes_ctrl_lsfr_23_cycles_1_n14, aes_ctrl_lsfr_23_cycles_1_n13,
         aes_ctrl_lsfr_23_cycles_1_n11, aes_ctrl_lsfr_23_cycles_1_n10,
         aes_ctrl_lsfr_23_cycles_1_n8, aes_ctrl_lsfr_23_cycles_1_n7,
         aes_ctrl_lsfr_23_cycles_1_n5, aes_ctrl_lsfr_23_cycles_1_n3,
         aes_ctrl_lsfr_23_cycles_1_n1, aes_ctrl_lsfr_23_cycles_1_n39,
         aes_ctrl_lsfr_23_cycles_1_n38, aes_ctrl_lsfr_23_cycles_1_n37,
         aes_ctrl_lsfr_23_cycles_1_n36, aes_ctrl_lsfr_23_cycles_1_n35,
         aes_ctrl_lsfr_23_cycles_1_n12, aes_ctrl_lsfr_23_cycles_1_n9,
         aes_ctrl_lsfr_23_cycles_1_n6, aes_ctrl_lsfr_23_cycles_1_n4,
         aes_ctrl_lsfr_23_cycles_1_n2, aes_ctrl_lsfr_23_cycles_1_N83,
         aes_ctrl_lsfr_23_cycles_1_N66, aes_ctrl_lsfr_23_cycles_1_N16,
         rcon_1_n45, rcon_1_n44, rcon_1_n43, rcon_1_n42, rcon_1_n41,
         rcon_1_n40, rcon_1_n39, rcon_1_n38, rcon_1_n37, rcon_1_n36,
         rcon_1_n34, rcon_1_n33, rcon_1_n32, rcon_1_n31, rcon_1_n30,
         rcon_1_n29, rcon_1_n28, rcon_1_n16, rcon_1_n15, rcon_1_n14,
         rcon_1_n13, rcon_1_n12, rcon_1_n11, rcon_1_n35, rcon_1_n26,
         rcon_1_n25, rcon_1_n24, rcon_1_n23, rcon_1_n22, rcon_1_n21,
         rcon_1_n20, rcon_1_n19, rcon_1_n18, rcon_1_n17, rcon_1_n9, rcon_1_n4,
         aes_sbox_n28, aes_sbox_n27, aes_sbox_n26, aes_sbox_n25, aes_sbox_n8,
         aes_sbox_n7, aes_sbox_n6, aes_sbox_n5, aes_sbox_n40, aes_sbox_n39,
         aes_sbox_n38, aes_sbox_n37, aes_sbox_n36, aes_sbox_n35, aes_sbox_n34,
         aes_sbox_n33, aes_sbox_n24, aes_sbox_n23, aes_sbox_n22, aes_sbox_n21,
         aes_sbox_n20, aes_sbox_n19, aes_sbox_n18, aes_sbox_n17, aes_sbox_n16,
         aes_sbox_n15, aes_sbox_n14, aes_sbox_n13, aes_sbox_n12, aes_sbox_n11,
         aes_sbox_n10, aes_sbox_n9, aes_sbox_InverterOutxD_0__0_,
         aes_sbox_InverterOutxD_0__1_, aes_sbox_InverterOutxD_0__2_,
         aes_sbox_InverterOutxD_0__3_, aes_sbox_InverterOutxD_1__0_,
         aes_sbox_InverterOutxD_1__1_, aes_sbox_InverterOutxD_1__2_,
         aes_sbox_InverterOutxD_1__3_, aes_sbox_InvMappedxD_0__0_,
         aes_sbox_InvMappedxD_0__1_, aes_sbox_InvMappedxD_0__5_,
         aes_sbox_InvMappedxD_0__6_, aes_sbox_mappedxD_0__0_,
         aes_sbox_mappedxD_0__1_, aes_sbox_mappedxD_0__3_,
         aes_sbox_mappedxD_0__4_, aes_sbox_mappedxD_0__5_,
         aes_sbox_mappedxD_0__6_, aes_sbox_mappedxD_0__7_,
         aes_sbox_mappedxD_1__0_, aes_sbox_mappedxD_1__1_,
         aes_sbox_mappedxD_1__3_, aes_sbox_mappedxD_1__4_,
         aes_sbox_mappedxD_1__5_, aes_sbox_mappedxD_1__6_,
         aes_sbox_mappedxD_1__7_, aes_sbox_Y0xD_0__0_, aes_sbox_Y0xD_0__1_,
         aes_sbox_Y0xD_0__2_, aes_sbox_Y0xD_0__3_, aes_sbox_Y0xD_1__0_,
         aes_sbox_Y0xD_1__1_, aes_sbox_Y0xD_1__2_, aes_sbox_Y0xD_1__3_,
         aes_sbox_Y1xD_0__0_, aes_sbox_Y1xD_0__1_, aes_sbox_Y1xD_0__2_,
         aes_sbox_Y1xD_0__3_, aes_sbox_Y1xD_1__0_, aes_sbox_Y1xD_1__1_,
         aes_sbox_Y1xD_1__2_, aes_sbox_Y1xD_1__3_,
         aes_sbox_input_mapping_1_n23, aes_sbox_input_mapping_1_n22,
         aes_sbox_input_mapping_1_n21, aes_sbox_input_mapping_1_n20,
         aes_sbox_input_mapping_1_n19, aes_sbox_input_mapping_1_n18,
         aes_sbox_input_mapping_1_n17, aes_sbox_output_mapping_1_n9,
         aes_sbox_output_mapping_1_n8, aes_sbox_output_mapping_1_n7,
         aes_sbox_input_mapping_0_n23, aes_sbox_input_mapping_0_n22,
         aes_sbox_input_mapping_0_n21, aes_sbox_input_mapping_0_n20,
         aes_sbox_input_mapping_0_n19, aes_sbox_input_mapping_0_n18,
         aes_sbox_input_mapping_0_n17, aes_sbox_output_mapping_0_n9,
         aes_sbox_output_mapping_0_n8, aes_sbox_output_mapping_0_n7,
         aes_sbox_mul_y0y1_n16, aes_sbox_mul_y0y1_n15, aes_sbox_mul_y0y1_n14,
         aes_sbox_mul_y0y1_n13, aes_sbox_mul_y0y1_n12, aes_sbox_mul_y0y1_n11,
         aes_sbox_mul_y0y1_n10, aes_sbox_mul_y0y1_n9, aes_sbox_mul_y0y1_n8,
         aes_sbox_mul_y0y1_n7, aes_sbox_mul_y0y1_n6, aes_sbox_mul_y0y1_n5,
         aes_sbox_mul_y0y1_n4, aes_sbox_mul_y0y1_n3, aes_sbox_mul_y0y1_n2,
         aes_sbox_mul_y0y1_n1, aes_sbox_mul_y0y1_Xi_mul_Yj_1__0_,
         aes_sbox_mul_y0y1_Xi_mul_Yj_1__1_, aes_sbox_mul_y0y1_Xi_mul_Yj_1__2_,
         aes_sbox_mul_y0y1_Xi_mul_Yj_1__3_, aes_sbox_mul_y0y1_Xi_mul_Yj_2__0_,
         aes_sbox_mul_y0y1_Xi_mul_Yj_2__1_, aes_sbox_mul_y0y1_Xi_mul_Yj_2__2_,
         aes_sbox_mul_y0y1_Xi_mul_Yj_2__3_, aes_sbox_mul_y0y1_gf4_mul_1_1_n77,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n76, aes_sbox_mul_y0y1_gf4_mul_1_1_n75,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n74, aes_sbox_mul_y0y1_gf4_mul_1_1_n73,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n72, aes_sbox_mul_y0y1_gf4_mul_1_1_n71,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n70, aes_sbox_mul_y0y1_gf4_mul_1_1_n69,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n68, aes_sbox_mul_y0y1_gf4_mul_1_1_n67,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n66, aes_sbox_mul_y0y1_gf4_mul_1_1_n65,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n64, aes_sbox_mul_y0y1_gf4_mul_1_1_n63,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n62, aes_sbox_mul_y0y1_gf4_mul_1_1_n61,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n60, aes_sbox_mul_y0y1_gf4_mul_1_1_n58,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n57, aes_sbox_mul_y0y1_gf4_mul_1_1_n56,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n55, aes_sbox_mul_y0y1_gf4_mul_1_1_n54,
         aes_sbox_mul_y0y1_gf4_mul_1_1_n53, aes_sbox_mul_y0y1_gf4_mul_1_0_n76,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n75, aes_sbox_mul_y0y1_gf4_mul_1_0_n74,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n73, aes_sbox_mul_y0y1_gf4_mul_1_0_n72,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n71, aes_sbox_mul_y0y1_gf4_mul_1_0_n70,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n69, aes_sbox_mul_y0y1_gf4_mul_1_0_n68,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n67, aes_sbox_mul_y0y1_gf4_mul_1_0_n66,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n65, aes_sbox_mul_y0y1_gf4_mul_1_0_n64,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n63, aes_sbox_mul_y0y1_gf4_mul_1_0_n62,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n61, aes_sbox_mul_y0y1_gf4_mul_1_0_n60,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n59, aes_sbox_mul_y0y1_gf4_mul_1_0_n58,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n57, aes_sbox_mul_y0y1_gf4_mul_1_0_n56,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n55, aes_sbox_mul_y0y1_gf4_mul_1_0_n54,
         aes_sbox_mul_y0y1_gf4_mul_1_0_n53, aes_sbox_mul_y0y1_gf4_mul_0_1_n76,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n75, aes_sbox_mul_y0y1_gf4_mul_0_1_n74,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n73, aes_sbox_mul_y0y1_gf4_mul_0_1_n72,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n71, aes_sbox_mul_y0y1_gf4_mul_0_1_n70,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n69, aes_sbox_mul_y0y1_gf4_mul_0_1_n68,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n67, aes_sbox_mul_y0y1_gf4_mul_0_1_n66,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n65, aes_sbox_mul_y0y1_gf4_mul_0_1_n64,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n63, aes_sbox_mul_y0y1_gf4_mul_0_1_n62,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n61, aes_sbox_mul_y0y1_gf4_mul_0_1_n60,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n59, aes_sbox_mul_y0y1_gf4_mul_0_1_n58,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n57, aes_sbox_mul_y0y1_gf4_mul_0_1_n56,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n55, aes_sbox_mul_y0y1_gf4_mul_0_1_n54,
         aes_sbox_mul_y0y1_gf4_mul_0_1_n53, aes_sbox_mul_y0y1_gf4_mul_0_0_n77,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n76, aes_sbox_mul_y0y1_gf4_mul_0_0_n75,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n74, aes_sbox_mul_y0y1_gf4_mul_0_0_n73,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n72, aes_sbox_mul_y0y1_gf4_mul_0_0_n71,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n70, aes_sbox_mul_y0y1_gf4_mul_0_0_n69,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n68, aes_sbox_mul_y0y1_gf4_mul_0_0_n67,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n66, aes_sbox_mul_y0y1_gf4_mul_0_0_n65,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n64, aes_sbox_mul_y0y1_gf4_mul_0_0_n63,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n62, aes_sbox_mul_y0y1_gf4_mul_0_0_n61,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n60, aes_sbox_mul_y0y1_gf4_mul_0_0_n59,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n58, aes_sbox_mul_y0y1_gf4_mul_0_0_n57,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n56, aes_sbox_mul_y0y1_gf4_mul_0_0_n55,
         aes_sbox_mul_y0y1_gf4_mul_0_0_n54, aes_sbox_inverter_gf24_n2,
         aes_sbox_inverter_gf24_n1, aes_sbox_inverter_gf24_n8,
         aes_sbox_inverter_gf24_n7, aes_sbox_inverter_gf24_n6,
         aes_sbox_inverter_gf24_n5, aes_sbox_inverter_gf24_n4,
         aes_sbox_inverter_gf24_n3, aes_sbox_inverter_gf24_d_0__0_,
         aes_sbox_inverter_gf24_d_1__0_, aes_sbox_inverter_gf24_ExDP_0__0_,
         aes_sbox_inverter_gf24_ExDP_0__1_, aes_sbox_inverter_gf24_ExDP_1__0_,
         aes_sbox_inverter_gf24_ExDP_1__1_, aes_sbox_inverter_gf24_a_mul_b_n8,
         aes_sbox_inverter_gf24_a_mul_b_n7, aes_sbox_inverter_gf24_a_mul_b_n6,
         aes_sbox_inverter_gf24_a_mul_b_n5, aes_sbox_inverter_gf24_a_mul_b_n4,
         aes_sbox_inverter_gf24_a_mul_b_n3, aes_sbox_inverter_gf24_a_mul_b_n2,
         aes_sbox_inverter_gf24_a_mul_b_n1,
         aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_,
         aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_,
         aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_,
         aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n14,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n13,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n12,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n11,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n14,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n13,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n12,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n11,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n14,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n13,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n12,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n11,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n14,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n13,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n12,
         aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n11,
         aes_sbox_inverter_gf24_a_mul_e_n16,
         aes_sbox_inverter_gf24_a_mul_e_n15,
         aes_sbox_inverter_gf24_a_mul_e_n14,
         aes_sbox_inverter_gf24_a_mul_e_n13,
         aes_sbox_inverter_gf24_a_mul_e_n12,
         aes_sbox_inverter_gf24_a_mul_e_n11,
         aes_sbox_inverter_gf24_a_mul_e_n10, aes_sbox_inverter_gf24_a_mul_e_n9,
         aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_,
         aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_,
         aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_,
         aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n14,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n13,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n12,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n11,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n14,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n13,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n12,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n11,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n14,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n13,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n12,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n11,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n14,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n13,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n12,
         aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n11,
         aes_sbox_inverter_gf24_b_mul_e_n16,
         aes_sbox_inverter_gf24_b_mul_e_n15,
         aes_sbox_inverter_gf24_b_mul_e_n14,
         aes_sbox_inverter_gf24_b_mul_e_n13,
         aes_sbox_inverter_gf24_b_mul_e_n12,
         aes_sbox_inverter_gf24_b_mul_e_n11,
         aes_sbox_inverter_gf24_b_mul_e_n10, aes_sbox_inverter_gf24_b_mul_e_n9,
         aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_,
         aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_,
         aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_,
         aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n14,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n13,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n12,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n11,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n14,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n13,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n12,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n11,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n14,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n13,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n12,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n11,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n14,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n13,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n12,
         aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n11, aes_sbox_mult_msb_n16,
         aes_sbox_mult_msb_n15, aes_sbox_mult_msb_n14, aes_sbox_mult_msb_n13,
         aes_sbox_mult_msb_n12, aes_sbox_mult_msb_n11, aes_sbox_mult_msb_n10,
         aes_sbox_mult_msb_n9, aes_sbox_mult_msb_n8, aes_sbox_mult_msb_n7,
         aes_sbox_mult_msb_n6, aes_sbox_mult_msb_n5, aes_sbox_mult_msb_n4,
         aes_sbox_mult_msb_n3, aes_sbox_mult_msb_n2, aes_sbox_mult_msb_n1,
         aes_sbox_mult_msb_Xi_mul_Yj_1__0_, aes_sbox_mult_msb_Xi_mul_Yj_1__1_,
         aes_sbox_mult_msb_Xi_mul_Yj_1__2_, aes_sbox_mult_msb_Xi_mul_Yj_1__3_,
         aes_sbox_mult_msb_Xi_mul_Yj_2__0_, aes_sbox_mult_msb_Xi_mul_Yj_2__1_,
         aes_sbox_mult_msb_Xi_mul_Yj_2__2_, aes_sbox_mult_msb_Xi_mul_Yj_2__3_,
         aes_sbox_mult_msb_gf4_mul_1_1_n77, aes_sbox_mult_msb_gf4_mul_1_1_n76,
         aes_sbox_mult_msb_gf4_mul_1_1_n75, aes_sbox_mult_msb_gf4_mul_1_1_n74,
         aes_sbox_mult_msb_gf4_mul_1_1_n73, aes_sbox_mult_msb_gf4_mul_1_1_n72,
         aes_sbox_mult_msb_gf4_mul_1_1_n71, aes_sbox_mult_msb_gf4_mul_1_1_n70,
         aes_sbox_mult_msb_gf4_mul_1_1_n69, aes_sbox_mult_msb_gf4_mul_1_1_n68,
         aes_sbox_mult_msb_gf4_mul_1_1_n67, aes_sbox_mult_msb_gf4_mul_1_1_n66,
         aes_sbox_mult_msb_gf4_mul_1_1_n65, aes_sbox_mult_msb_gf4_mul_1_1_n64,
         aes_sbox_mult_msb_gf4_mul_1_1_n63, aes_sbox_mult_msb_gf4_mul_1_1_n62,
         aes_sbox_mult_msb_gf4_mul_1_1_n61, aes_sbox_mult_msb_gf4_mul_1_1_n60,
         aes_sbox_mult_msb_gf4_mul_1_1_n59, aes_sbox_mult_msb_gf4_mul_1_1_n58,
         aes_sbox_mult_msb_gf4_mul_1_1_n57, aes_sbox_mult_msb_gf4_mul_1_1_n56,
         aes_sbox_mult_msb_gf4_mul_1_1_n55, aes_sbox_mult_msb_gf4_mul_1_1_n54,
         aes_sbox_mult_msb_gf4_mul_1_0_n76, aes_sbox_mult_msb_gf4_mul_1_0_n75,
         aes_sbox_mult_msb_gf4_mul_1_0_n74, aes_sbox_mult_msb_gf4_mul_1_0_n73,
         aes_sbox_mult_msb_gf4_mul_1_0_n72, aes_sbox_mult_msb_gf4_mul_1_0_n71,
         aes_sbox_mult_msb_gf4_mul_1_0_n70, aes_sbox_mult_msb_gf4_mul_1_0_n69,
         aes_sbox_mult_msb_gf4_mul_1_0_n68, aes_sbox_mult_msb_gf4_mul_1_0_n67,
         aes_sbox_mult_msb_gf4_mul_1_0_n66, aes_sbox_mult_msb_gf4_mul_1_0_n65,
         aes_sbox_mult_msb_gf4_mul_1_0_n64, aes_sbox_mult_msb_gf4_mul_1_0_n63,
         aes_sbox_mult_msb_gf4_mul_1_0_n62, aes_sbox_mult_msb_gf4_mul_1_0_n61,
         aes_sbox_mult_msb_gf4_mul_1_0_n60, aes_sbox_mult_msb_gf4_mul_1_0_n59,
         aes_sbox_mult_msb_gf4_mul_1_0_n58, aes_sbox_mult_msb_gf4_mul_1_0_n57,
         aes_sbox_mult_msb_gf4_mul_1_0_n56, aes_sbox_mult_msb_gf4_mul_1_0_n55,
         aes_sbox_mult_msb_gf4_mul_1_0_n54, aes_sbox_mult_msb_gf4_mul_1_0_n53,
         aes_sbox_mult_msb_gf4_mul_0_1_n77, aes_sbox_mult_msb_gf4_mul_0_1_n76,
         aes_sbox_mult_msb_gf4_mul_0_1_n75, aes_sbox_mult_msb_gf4_mul_0_1_n74,
         aes_sbox_mult_msb_gf4_mul_0_1_n73, aes_sbox_mult_msb_gf4_mul_0_1_n72,
         aes_sbox_mult_msb_gf4_mul_0_1_n71, aes_sbox_mult_msb_gf4_mul_0_1_n70,
         aes_sbox_mult_msb_gf4_mul_0_1_n69, aes_sbox_mult_msb_gf4_mul_0_1_n68,
         aes_sbox_mult_msb_gf4_mul_0_1_n67, aes_sbox_mult_msb_gf4_mul_0_1_n66,
         aes_sbox_mult_msb_gf4_mul_0_1_n65, aes_sbox_mult_msb_gf4_mul_0_1_n64,
         aes_sbox_mult_msb_gf4_mul_0_1_n63, aes_sbox_mult_msb_gf4_mul_0_1_n62,
         aes_sbox_mult_msb_gf4_mul_0_1_n61, aes_sbox_mult_msb_gf4_mul_0_1_n60,
         aes_sbox_mult_msb_gf4_mul_0_1_n59, aes_sbox_mult_msb_gf4_mul_0_1_n58,
         aes_sbox_mult_msb_gf4_mul_0_1_n57, aes_sbox_mult_msb_gf4_mul_0_1_n56,
         aes_sbox_mult_msb_gf4_mul_0_1_n55, aes_sbox_mult_msb_gf4_mul_0_1_n54,
         aes_sbox_mult_msb_gf4_mul_0_0_n76, aes_sbox_mult_msb_gf4_mul_0_0_n75,
         aes_sbox_mult_msb_gf4_mul_0_0_n74, aes_sbox_mult_msb_gf4_mul_0_0_n73,
         aes_sbox_mult_msb_gf4_mul_0_0_n72, aes_sbox_mult_msb_gf4_mul_0_0_n71,
         aes_sbox_mult_msb_gf4_mul_0_0_n70, aes_sbox_mult_msb_gf4_mul_0_0_n69,
         aes_sbox_mult_msb_gf4_mul_0_0_n68, aes_sbox_mult_msb_gf4_mul_0_0_n67,
         aes_sbox_mult_msb_gf4_mul_0_0_n66, aes_sbox_mult_msb_gf4_mul_0_0_n65,
         aes_sbox_mult_msb_gf4_mul_0_0_n64, aes_sbox_mult_msb_gf4_mul_0_0_n63,
         aes_sbox_mult_msb_gf4_mul_0_0_n62, aes_sbox_mult_msb_gf4_mul_0_0_n61,
         aes_sbox_mult_msb_gf4_mul_0_0_n60, aes_sbox_mult_msb_gf4_mul_0_0_n59,
         aes_sbox_mult_msb_gf4_mul_0_0_n58, aes_sbox_mult_msb_gf4_mul_0_0_n57,
         aes_sbox_mult_msb_gf4_mul_0_0_n56, aes_sbox_mult_msb_gf4_mul_0_0_n55,
         aes_sbox_mult_msb_gf4_mul_0_0_n54, aes_sbox_mult_msb_gf4_mul_0_0_n53,
         aes_sbox_mult_lsb_n16, aes_sbox_mult_lsb_n15, aes_sbox_mult_lsb_n14,
         aes_sbox_mult_lsb_n13, aes_sbox_mult_lsb_n12, aes_sbox_mult_lsb_n11,
         aes_sbox_mult_lsb_n10, aes_sbox_mult_lsb_n9, aes_sbox_mult_lsb_n8,
         aes_sbox_mult_lsb_n7, aes_sbox_mult_lsb_n6, aes_sbox_mult_lsb_n5,
         aes_sbox_mult_lsb_n4, aes_sbox_mult_lsb_n3, aes_sbox_mult_lsb_n2,
         aes_sbox_mult_lsb_n1, aes_sbox_mult_lsb_Xi_mul_Yj_1__0_,
         aes_sbox_mult_lsb_Xi_mul_Yj_1__1_, aes_sbox_mult_lsb_Xi_mul_Yj_1__2_,
         aes_sbox_mult_lsb_Xi_mul_Yj_1__3_, aes_sbox_mult_lsb_Xi_mul_Yj_2__0_,
         aes_sbox_mult_lsb_Xi_mul_Yj_2__1_, aes_sbox_mult_lsb_Xi_mul_Yj_2__2_,
         aes_sbox_mult_lsb_Xi_mul_Yj_2__3_, aes_sbox_mult_lsb_gf4_mul_1_1_n76,
         aes_sbox_mult_lsb_gf4_mul_1_1_n75, aes_sbox_mult_lsb_gf4_mul_1_1_n74,
         aes_sbox_mult_lsb_gf4_mul_1_1_n73, aes_sbox_mult_lsb_gf4_mul_1_1_n72,
         aes_sbox_mult_lsb_gf4_mul_1_1_n71, aes_sbox_mult_lsb_gf4_mul_1_1_n70,
         aes_sbox_mult_lsb_gf4_mul_1_1_n69, aes_sbox_mult_lsb_gf4_mul_1_1_n68,
         aes_sbox_mult_lsb_gf4_mul_1_1_n67, aes_sbox_mult_lsb_gf4_mul_1_1_n66,
         aes_sbox_mult_lsb_gf4_mul_1_1_n65, aes_sbox_mult_lsb_gf4_mul_1_1_n64,
         aes_sbox_mult_lsb_gf4_mul_1_1_n63, aes_sbox_mult_lsb_gf4_mul_1_1_n62,
         aes_sbox_mult_lsb_gf4_mul_1_1_n61, aes_sbox_mult_lsb_gf4_mul_1_1_n60,
         aes_sbox_mult_lsb_gf4_mul_1_1_n59, aes_sbox_mult_lsb_gf4_mul_1_1_n58,
         aes_sbox_mult_lsb_gf4_mul_1_1_n57, aes_sbox_mult_lsb_gf4_mul_1_1_n56,
         aes_sbox_mult_lsb_gf4_mul_1_1_n55, aes_sbox_mult_lsb_gf4_mul_1_1_n54,
         aes_sbox_mult_lsb_gf4_mul_1_1_n53, aes_sbox_mult_lsb_gf4_mul_1_0_n76,
         aes_sbox_mult_lsb_gf4_mul_1_0_n75, aes_sbox_mult_lsb_gf4_mul_1_0_n74,
         aes_sbox_mult_lsb_gf4_mul_1_0_n73, aes_sbox_mult_lsb_gf4_mul_1_0_n72,
         aes_sbox_mult_lsb_gf4_mul_1_0_n71, aes_sbox_mult_lsb_gf4_mul_1_0_n70,
         aes_sbox_mult_lsb_gf4_mul_1_0_n69, aes_sbox_mult_lsb_gf4_mul_1_0_n68,
         aes_sbox_mult_lsb_gf4_mul_1_0_n67, aes_sbox_mult_lsb_gf4_mul_1_0_n66,
         aes_sbox_mult_lsb_gf4_mul_1_0_n65, aes_sbox_mult_lsb_gf4_mul_1_0_n64,
         aes_sbox_mult_lsb_gf4_mul_1_0_n63, aes_sbox_mult_lsb_gf4_mul_1_0_n62,
         aes_sbox_mult_lsb_gf4_mul_1_0_n61, aes_sbox_mult_lsb_gf4_mul_1_0_n60,
         aes_sbox_mult_lsb_gf4_mul_1_0_n59, aes_sbox_mult_lsb_gf4_mul_1_0_n58,
         aes_sbox_mult_lsb_gf4_mul_1_0_n57, aes_sbox_mult_lsb_gf4_mul_1_0_n56,
         aes_sbox_mult_lsb_gf4_mul_1_0_n55, aes_sbox_mult_lsb_gf4_mul_1_0_n54,
         aes_sbox_mult_lsb_gf4_mul_1_0_n53, aes_sbox_mult_lsb_gf4_mul_0_1_n76,
         aes_sbox_mult_lsb_gf4_mul_0_1_n75, aes_sbox_mult_lsb_gf4_mul_0_1_n74,
         aes_sbox_mult_lsb_gf4_mul_0_1_n73, aes_sbox_mult_lsb_gf4_mul_0_1_n72,
         aes_sbox_mult_lsb_gf4_mul_0_1_n71, aes_sbox_mult_lsb_gf4_mul_0_1_n70,
         aes_sbox_mult_lsb_gf4_mul_0_1_n69, aes_sbox_mult_lsb_gf4_mul_0_1_n68,
         aes_sbox_mult_lsb_gf4_mul_0_1_n67, aes_sbox_mult_lsb_gf4_mul_0_1_n66,
         aes_sbox_mult_lsb_gf4_mul_0_1_n65, aes_sbox_mult_lsb_gf4_mul_0_1_n64,
         aes_sbox_mult_lsb_gf4_mul_0_1_n63, aes_sbox_mult_lsb_gf4_mul_0_1_n62,
         aes_sbox_mult_lsb_gf4_mul_0_1_n61, aes_sbox_mult_lsb_gf4_mul_0_1_n60,
         aes_sbox_mult_lsb_gf4_mul_0_1_n59, aes_sbox_mult_lsb_gf4_mul_0_1_n58,
         aes_sbox_mult_lsb_gf4_mul_0_1_n57, aes_sbox_mult_lsb_gf4_mul_0_1_n56,
         aes_sbox_mult_lsb_gf4_mul_0_1_n55, aes_sbox_mult_lsb_gf4_mul_0_1_n54,
         aes_sbox_mult_lsb_gf4_mul_0_1_n53, aes_sbox_mult_lsb_gf4_mul_0_0_n76,
         aes_sbox_mult_lsb_gf4_mul_0_0_n75, aes_sbox_mult_lsb_gf4_mul_0_0_n74,
         aes_sbox_mult_lsb_gf4_mul_0_0_n73, aes_sbox_mult_lsb_gf4_mul_0_0_n72,
         aes_sbox_mult_lsb_gf4_mul_0_0_n71, aes_sbox_mult_lsb_gf4_mul_0_0_n70,
         aes_sbox_mult_lsb_gf4_mul_0_0_n69, aes_sbox_mult_lsb_gf4_mul_0_0_n68,
         aes_sbox_mult_lsb_gf4_mul_0_0_n67, aes_sbox_mult_lsb_gf4_mul_0_0_n66,
         aes_sbox_mult_lsb_gf4_mul_0_0_n65, aes_sbox_mult_lsb_gf4_mul_0_0_n64,
         aes_sbox_mult_lsb_gf4_mul_0_0_n63, aes_sbox_mult_lsb_gf4_mul_0_0_n62,
         aes_sbox_mult_lsb_gf4_mul_0_0_n61, aes_sbox_mult_lsb_gf4_mul_0_0_n60,
         aes_sbox_mult_lsb_gf4_mul_0_0_n59, aes_sbox_mult_lsb_gf4_mul_0_0_n58,
         aes_sbox_mult_lsb_gf4_mul_0_0_n57, aes_sbox_mult_lsb_gf4_mul_0_0_n56,
         aes_sbox_mult_lsb_gf4_mul_0_0_n55, aes_sbox_mult_lsb_gf4_mul_0_0_n54,
         aes_sbox_mult_lsb_gf4_mul_0_0_n53, aes_key_regs_1_n4,
         aes_key_regs_1_K02xDP_0_, aes_key_regs_1_K02xDP_1_,
         aes_key_regs_1_K02xDP_2_, aes_key_regs_1_K02xDP_3_,
         aes_key_regs_1_K02xDP_4_, aes_key_regs_1_K02xDP_5_,
         aes_key_regs_1_K02xDP_6_, aes_key_regs_1_K02xDP_7_,
         aes_key_regs_1_K01xDP_0_, aes_key_regs_1_K01xDP_1_,
         aes_key_regs_1_K01xDP_2_, aes_key_regs_1_K01xDP_3_,
         aes_key_regs_1_K01xDP_4_, aes_key_regs_1_K01xDP_5_,
         aes_key_regs_1_K01xDP_6_, aes_key_regs_1_K01xDP_7_,
         aes_state_regs_1_n113, aes_state_regs_1_n112, aes_state_regs_1_n111,
         aes_state_regs_1_n110, aes_state_regs_1_n109, aes_state_regs_1_n108,
         aes_state_regs_1_n107, aes_state_regs_1_n106, aes_state_regs_1_n81,
         aes_state_regs_1_n80, aes_state_regs_1_n79, aes_state_regs_1_n78,
         aes_state_regs_1_n77, aes_state_regs_1_n76, aes_state_regs_1_n75,
         aes_state_regs_1_n74, aes_state_regs_1_n73, aes_state_regs_1_n72,
         aes_state_regs_1_n71, aes_state_regs_1_n70, aes_state_regs_1_n69,
         aes_state_regs_1_n68, aes_state_regs_1_n67, aes_state_regs_1_n66,
         aes_state_regs_1_n65, aes_state_regs_1_n64, aes_state_regs_1_n63,
         aes_state_regs_1_n56, aes_state_regs_1_n46, aes_state_regs_1_n45,
         aes_state_regs_1_n105, aes_state_regs_1_n104, aes_state_regs_1_n103,
         aes_state_regs_1_n102, aes_state_regs_1_n101, aes_state_regs_1_n100,
         aes_state_regs_1_n99, aes_state_regs_1_n98, aes_state_regs_1_n97,
         aes_state_regs_1_n96, aes_state_regs_1_n95, aes_state_regs_1_n94,
         aes_state_regs_1_n93, aes_state_regs_1_n92, aes_state_regs_1_n91,
         aes_state_regs_1_n90, aes_state_regs_1_n89, aes_state_regs_1_n88,
         aes_state_regs_1_n87, aes_state_regs_1_n86, aes_state_regs_1_n85,
         aes_state_regs_1_n84, aes_state_regs_1_n83, aes_state_regs_1_n82,
         aes_state_regs_1_n62, aes_state_regs_1_n61, aes_state_regs_1_n60,
         aes_state_regs_1_n59, aes_state_regs_1_n58, aes_state_regs_1_n57,
         aes_state_regs_1_n55, aes_state_regs_1_n54, aes_state_regs_1_n53,
         aes_state_regs_1_n52, aes_state_regs_1_n51, aes_state_regs_1_n50,
         aes_state_regs_1_n49, aes_state_regs_1_n48, aes_state_regs_1_n47,
         aes_state_regs_1_n38, aes_state_regs_1_n37, aes_state_regs_1_n36,
         aes_state_regs_1_n35, aes_state_regs_1_n34, aes_state_regs_1_n33,
         aes_state_regs_1_n32, aes_state_regs_1_n31, aes_state_regs_1_n30,
         aes_state_regs_1_n29, aes_state_regs_1_n28, aes_state_regs_1_n27,
         aes_state_regs_1_n26, aes_state_regs_1_n25, aes_state_regs_1_n24,
         aes_state_regs_1_n23, aes_state_regs_1_n22, aes_state_regs_1_n21,
         aes_state_regs_1_n20, aes_state_regs_1_n19, aes_state_regs_1_n18,
         aes_state_regs_1_n17, aes_state_regs_1_n16, aes_state_regs_1_n15,
         aes_state_regs_1_n14, aes_state_regs_1_n13, aes_state_regs_1_n12,
         aes_state_regs_1_n11, aes_state_regs_1_n10, aes_state_regs_1_n9,
         aes_state_regs_1_n8, aes_state_regs_1_n7, aes_state_regs_1_n6,
         aes_state_regs_1_n5, aes_state_regs_1_n4, aes_state_regs_1_n3,
         aes_state_regs_1_n2, aes_state_regs_1_n1, aes_state_regs_1_S03xDP_0_,
         aes_state_regs_1_S02xDP_0_, aes_state_regs_1_S02xDP_1_,
         aes_state_regs_1_S02xDP_2_, aes_state_regs_1_S02xDP_3_,
         aes_state_regs_1_S02xDP_4_, aes_state_regs_1_S02xDP_5_,
         aes_state_regs_1_S02xDP_6_, aes_state_regs_1_S02xDP_7_,
         aes_state_regs_1_S31xDP_0_, aes_state_regs_1_S30xDP_0_,
         aes_state_regs_1_S30xDP_1_, aes_state_regs_1_S30xDP_2_,
         aes_state_regs_1_S30xDP_3_, aes_state_regs_1_S30xDP_4_,
         aes_state_regs_1_S30xDP_5_, aes_state_regs_1_S30xDP_6_,
         aes_state_regs_1_S30xDP_7_, aes_state_regs_1_S20xDP_0_,
         aes_state_regs_1_S20xDP_1_, aes_state_regs_1_S20xDP_2_,
         aes_state_regs_1_S20xDP_3_, aes_state_regs_1_S20xDP_4_,
         aes_state_regs_1_S20xDP_5_, aes_state_regs_1_S20xDP_6_,
         aes_state_regs_1_S20xDP_7_, aes_state_regs_1_S23xDP_0_,
         aes_state_regs_1_S23xDP_1_, aes_state_regs_1_S23xDP_2_,
         aes_state_regs_1_S23xDP_3_, aes_state_regs_1_S23xDP_4_,
         aes_state_regs_1_S23xDP_5_, aes_state_regs_1_S23xDP_6_,
         aes_state_regs_1_S23xDP_7_, aes_state_regs_1_S22xDP_0_,
         aes_state_regs_1_S10xDP_0_, aes_state_regs_1_S10xDP_1_,
         aes_state_regs_1_S10xDP_2_, aes_state_regs_1_S10xDP_3_,
         aes_state_regs_1_S10xDP_4_, aes_state_regs_1_S10xDP_5_,
         aes_state_regs_1_S10xDP_6_, aes_state_regs_1_S10xDP_7_,
         aes_state_regs_1_S01xDO_0_, aes_state_regs_1_S01xDO_1_,
         aes_state_regs_1_S01xDO_2_, aes_state_regs_1_S01xDO_3_,
         aes_state_regs_1_S01xDO_4_, aes_state_regs_1_S01xDO_5_,
         aes_state_regs_1_S01xDO_6_, aes_state_regs_1_S01xDO_7_,
         aes_state_regs_1_mix_columns_1_n245,
         aes_state_regs_1_mix_columns_1_n244,
         aes_state_regs_1_mix_columns_1_n243,
         aes_state_regs_1_mix_columns_1_n242,
         aes_state_regs_1_mix_columns_1_n241,
         aes_state_regs_1_mix_columns_1_n240,
         aes_state_regs_1_mix_columns_1_n239,
         aes_state_regs_1_mix_columns_1_n238,
         aes_state_regs_1_mix_columns_1_n237,
         aes_state_regs_1_mix_columns_1_n236,
         aes_state_regs_1_mix_columns_1_n235,
         aes_state_regs_1_mix_columns_1_n234,
         aes_state_regs_1_mix_columns_1_n233,
         aes_state_regs_1_mix_columns_1_n232,
         aes_state_regs_1_mix_columns_1_n231,
         aes_state_regs_1_mix_columns_1_n230,
         aes_state_regs_1_mix_columns_1_n229,
         aes_state_regs_1_mix_columns_1_n228,
         aes_state_regs_1_mix_columns_1_n227,
         aes_state_regs_1_mix_columns_1_n226,
         aes_state_regs_1_mix_columns_1_n225,
         aes_state_regs_1_mix_columns_1_n224,
         aes_state_regs_1_mix_columns_1_n223,
         aes_state_regs_1_mix_columns_1_n222,
         aes_state_regs_1_mix_columns_1_n221,
         aes_state_regs_1_mix_columns_1_n220,
         aes_state_regs_1_mix_columns_1_n219,
         aes_state_regs_1_mix_columns_1_n218,
         aes_state_regs_1_mix_columns_1_n217,
         aes_state_regs_1_mix_columns_1_n216,
         aes_state_regs_1_mix_columns_1_n215,
         aes_state_regs_1_mix_columns_1_n214,
         aes_state_regs_1_mix_columns_1_n213,
         aes_state_regs_1_mix_columns_1_n212,
         aes_state_regs_1_mix_columns_1_n211,
         aes_state_regs_1_mix_columns_1_n210,
         aes_state_regs_1_mix_columns_1_n209,
         aes_state_regs_1_mix_columns_1_n208,
         aes_state_regs_1_mix_columns_1_n207,
         aes_state_regs_1_mix_columns_1_n206,
         aes_state_regs_1_mix_columns_1_n205,
         aes_state_regs_1_mix_columns_1_n204,
         aes_state_regs_1_mix_columns_1_n203,
         aes_state_regs_1_mix_columns_1_n202,
         aes_state_regs_1_mix_columns_1_n201,
         aes_state_regs_1_mix_columns_1_n200,
         aes_state_regs_1_mix_columns_1_n199,
         aes_state_regs_1_mix_columns_1_n198,
         aes_state_regs_1_mix_columns_1_n197,
         aes_state_regs_1_mix_columns_1_n196,
         aes_state_regs_1_mix_columns_1_n195,
         aes_state_regs_1_mix_columns_1_n194,
         aes_state_regs_1_mix_columns_1_n193,
         aes_state_regs_1_mix_columns_1_n192,
         aes_state_regs_1_mix_columns_1_n191,
         aes_state_regs_1_mix_columns_1_n190,
         aes_state_regs_1_mix_columns_1_n189,
         aes_state_regs_1_mix_columns_1_n188,
         aes_state_regs_1_mix_columns_1_n187,
         aes_state_regs_1_mix_columns_1_n186,
         aes_state_regs_1_mix_columns_1_n185,
         aes_state_regs_1_mix_columns_1_n184,
         aes_state_regs_1_mix_columns_1_n183,
         aes_state_regs_1_mix_columns_1_n182,
         aes_state_regs_1_mix_columns_1_n181,
         aes_state_regs_1_mix_columns_1_n180,
         aes_state_regs_1_mix_columns_1_n179,
         aes_state_regs_1_mix_columns_1_n178,
         aes_state_regs_1_mix_columns_1_n177,
         aes_state_regs_1_mix_columns_1_n176,
         aes_state_regs_1_mix_columns_1_n175,
         aes_state_regs_1_mix_columns_1_n174,
         aes_state_regs_1_mix_columns_1_n173,
         aes_state_regs_1_mix_columns_1_n172,
         aes_state_regs_1_mix_columns_1_n171,
         aes_state_regs_1_mix_columns_1_n170,
         aes_state_regs_1_mix_columns_1_n169,
         aes_state_regs_1_mix_columns_1_n168,
         aes_state_regs_1_mix_columns_1_n167,
         aes_state_regs_1_mix_columns_1_n166,
         aes_state_regs_1_mix_columns_1_n165,
         aes_state_regs_1_mix_columns_1_n164,
         aes_state_regs_1_mix_columns_1_n163,
         aes_state_regs_1_mix_columns_1_n162,
         aes_state_regs_1_mix_columns_1_n161,
         aes_state_regs_1_mix_columns_1_n160,
         aes_state_regs_1_mix_columns_1_n159, aes_key_regs_0_n4,
         aes_key_regs_0_K02xDP_0_, aes_key_regs_0_K02xDP_1_,
         aes_key_regs_0_K02xDP_2_, aes_key_regs_0_K02xDP_3_,
         aes_key_regs_0_K02xDP_4_, aes_key_regs_0_K02xDP_5_,
         aes_key_regs_0_K02xDP_6_, aes_key_regs_0_K02xDP_7_,
         aes_key_regs_0_K01xDP_0_, aes_key_regs_0_K01xDP_1_,
         aes_key_regs_0_K01xDP_2_, aes_key_regs_0_K01xDP_3_,
         aes_key_regs_0_K01xDP_4_, aes_key_regs_0_K01xDP_5_,
         aes_key_regs_0_K01xDP_6_, aes_key_regs_0_K01xDP_7_,
         aes_state_regs_0_n202, aes_state_regs_0_n201, aes_state_regs_0_n200,
         aes_state_regs_0_n199, aes_state_regs_0_n198, aes_state_regs_0_n197,
         aes_state_regs_0_n196, aes_state_regs_0_n195, aes_state_regs_0_n194,
         aes_state_regs_0_n193, aes_state_regs_0_n192, aes_state_regs_0_n191,
         aes_state_regs_0_n190, aes_state_regs_0_n189, aes_state_regs_0_n188,
         aes_state_regs_0_n187, aes_state_regs_0_n186, aes_state_regs_0_n185,
         aes_state_regs_0_n184, aes_state_regs_0_n183, aes_state_regs_0_n182,
         aes_state_regs_0_n181, aes_state_regs_0_n180, aes_state_regs_0_n179,
         aes_state_regs_0_n178, aes_state_regs_0_n177, aes_state_regs_0_n176,
         aes_state_regs_0_n175, aes_state_regs_0_n174, aes_state_regs_0_n51,
         aes_state_regs_0_n50, aes_state_regs_0_n49, aes_state_regs_0_n48,
         aes_state_regs_0_n47, aes_state_regs_0_n46, aes_state_regs_0_n45,
         aes_state_regs_0_n44, aes_state_regs_0_n43, aes_state_regs_0_n42,
         aes_state_regs_0_n41, aes_state_regs_0_n40, aes_state_regs_0_n39,
         aes_state_regs_0_n38, aes_state_regs_0_n37, aes_state_regs_0_n36,
         aes_state_regs_0_n35, aes_state_regs_0_n34, aes_state_regs_0_n33,
         aes_state_regs_0_n32, aes_state_regs_0_n31, aes_state_regs_0_n30,
         aes_state_regs_0_n29, aes_state_regs_0_n28, aes_state_regs_0_n173,
         aes_state_regs_0_n172, aes_state_regs_0_n171, aes_state_regs_0_n170,
         aes_state_regs_0_n169, aes_state_regs_0_n168, aes_state_regs_0_n167,
         aes_state_regs_0_n166, aes_state_regs_0_n165, aes_state_regs_0_n164,
         aes_state_regs_0_n163, aes_state_regs_0_n162, aes_state_regs_0_n161,
         aes_state_regs_0_n160, aes_state_regs_0_n159, aes_state_regs_0_n158,
         aes_state_regs_0_n157, aes_state_regs_0_n156, aes_state_regs_0_n155,
         aes_state_regs_0_n154, aes_state_regs_0_n153, aes_state_regs_0_n152,
         aes_state_regs_0_n151, aes_state_regs_0_n150, aes_state_regs_0_n149,
         aes_state_regs_0_n148, aes_state_regs_0_n147, aes_state_regs_0_n146,
         aes_state_regs_0_n145, aes_state_regs_0_n144, aes_state_regs_0_n143,
         aes_state_regs_0_n142, aes_state_regs_0_n141, aes_state_regs_0_n140,
         aes_state_regs_0_n139, aes_state_regs_0_n138, aes_state_regs_0_n137,
         aes_state_regs_0_n136, aes_state_regs_0_n127, aes_state_regs_0_n126,
         aes_state_regs_0_n125, aes_state_regs_0_n124, aes_state_regs_0_n123,
         aes_state_regs_0_n122, aes_state_regs_0_n121, aes_state_regs_0_n109,
         aes_state_regs_0_S03xDP_0_, aes_state_regs_0_S02xDP_0_,
         aes_state_regs_0_S02xDP_1_, aes_state_regs_0_S02xDP_2_,
         aes_state_regs_0_S02xDP_3_, aes_state_regs_0_S02xDP_4_,
         aes_state_regs_0_S02xDP_5_, aes_state_regs_0_S02xDP_6_,
         aes_state_regs_0_S02xDP_7_, aes_state_regs_0_S31xDP_0_,
         aes_state_regs_0_S30xDP_0_, aes_state_regs_0_S30xDP_1_,
         aes_state_regs_0_S30xDP_2_, aes_state_regs_0_S30xDP_3_,
         aes_state_regs_0_S30xDP_4_, aes_state_regs_0_S30xDP_5_,
         aes_state_regs_0_S30xDP_6_, aes_state_regs_0_S30xDP_7_,
         aes_state_regs_0_S20xDP_0_, aes_state_regs_0_S20xDP_1_,
         aes_state_regs_0_S20xDP_2_, aes_state_regs_0_S20xDP_3_,
         aes_state_regs_0_S20xDP_4_, aes_state_regs_0_S20xDP_5_,
         aes_state_regs_0_S20xDP_6_, aes_state_regs_0_S20xDP_7_,
         aes_state_regs_0_S23xDP_0_, aes_state_regs_0_S23xDP_1_,
         aes_state_regs_0_S23xDP_2_, aes_state_regs_0_S23xDP_3_,
         aes_state_regs_0_S23xDP_4_, aes_state_regs_0_S23xDP_5_,
         aes_state_regs_0_S23xDP_6_, aes_state_regs_0_S23xDP_7_,
         aes_state_regs_0_S22xDP_0_, aes_state_regs_0_S10xDP_0_,
         aes_state_regs_0_S10xDP_1_, aes_state_regs_0_S10xDP_2_,
         aes_state_regs_0_S10xDP_3_, aes_state_regs_0_S10xDP_4_,
         aes_state_regs_0_S10xDP_5_, aes_state_regs_0_S10xDP_6_,
         aes_state_regs_0_S10xDP_7_, aes_state_regs_0_S01xDO_0_,
         aes_state_regs_0_S01xDO_1_, aes_state_regs_0_S01xDO_2_,
         aes_state_regs_0_S01xDO_3_, aes_state_regs_0_S01xDO_4_,
         aes_state_regs_0_S01xDO_5_, aes_state_regs_0_S01xDO_6_,
         aes_state_regs_0_S01xDO_7_, aes_state_regs_0_mix_columns_1_n245,
         aes_state_regs_0_mix_columns_1_n244,
         aes_state_regs_0_mix_columns_1_n243,
         aes_state_regs_0_mix_columns_1_n242,
         aes_state_regs_0_mix_columns_1_n241,
         aes_state_regs_0_mix_columns_1_n240,
         aes_state_regs_0_mix_columns_1_n239,
         aes_state_regs_0_mix_columns_1_n238,
         aes_state_regs_0_mix_columns_1_n237,
         aes_state_regs_0_mix_columns_1_n236,
         aes_state_regs_0_mix_columns_1_n235,
         aes_state_regs_0_mix_columns_1_n234,
         aes_state_regs_0_mix_columns_1_n233,
         aes_state_regs_0_mix_columns_1_n232,
         aes_state_regs_0_mix_columns_1_n231,
         aes_state_regs_0_mix_columns_1_n230,
         aes_state_regs_0_mix_columns_1_n229,
         aes_state_regs_0_mix_columns_1_n228,
         aes_state_regs_0_mix_columns_1_n227,
         aes_state_regs_0_mix_columns_1_n226,
         aes_state_regs_0_mix_columns_1_n225,
         aes_state_regs_0_mix_columns_1_n224,
         aes_state_regs_0_mix_columns_1_n223,
         aes_state_regs_0_mix_columns_1_n222,
         aes_state_regs_0_mix_columns_1_n221,
         aes_state_regs_0_mix_columns_1_n220,
         aes_state_regs_0_mix_columns_1_n219,
         aes_state_regs_0_mix_columns_1_n218,
         aes_state_regs_0_mix_columns_1_n217,
         aes_state_regs_0_mix_columns_1_n216,
         aes_state_regs_0_mix_columns_1_n215,
         aes_state_regs_0_mix_columns_1_n214,
         aes_state_regs_0_mix_columns_1_n213,
         aes_state_regs_0_mix_columns_1_n212,
         aes_state_regs_0_mix_columns_1_n211,
         aes_state_regs_0_mix_columns_1_n210,
         aes_state_regs_0_mix_columns_1_n209,
         aes_state_regs_0_mix_columns_1_n208,
         aes_state_regs_0_mix_columns_1_n207,
         aes_state_regs_0_mix_columns_1_n206,
         aes_state_regs_0_mix_columns_1_n205,
         aes_state_regs_0_mix_columns_1_n204,
         aes_state_regs_0_mix_columns_1_n203,
         aes_state_regs_0_mix_columns_1_n202,
         aes_state_regs_0_mix_columns_1_n201,
         aes_state_regs_0_mix_columns_1_n200,
         aes_state_regs_0_mix_columns_1_n199,
         aes_state_regs_0_mix_columns_1_n198,
         aes_state_regs_0_mix_columns_1_n197,
         aes_state_regs_0_mix_columns_1_n196,
         aes_state_regs_0_mix_columns_1_n195,
         aes_state_regs_0_mix_columns_1_n194,
         aes_state_regs_0_mix_columns_1_n193,
         aes_state_regs_0_mix_columns_1_n192,
         aes_state_regs_0_mix_columns_1_n191,
         aes_state_regs_0_mix_columns_1_n190,
         aes_state_regs_0_mix_columns_1_n189,
         aes_state_regs_0_mix_columns_1_n188,
         aes_state_regs_0_mix_columns_1_n187,
         aes_state_regs_0_mix_columns_1_n186,
         aes_state_regs_0_mix_columns_1_n185,
         aes_state_regs_0_mix_columns_1_n184,
         aes_state_regs_0_mix_columns_1_n183,
         aes_state_regs_0_mix_columns_1_n182,
         aes_state_regs_0_mix_columns_1_n181,
         aes_state_regs_0_mix_columns_1_n180,
         aes_state_regs_0_mix_columns_1_n179,
         aes_state_regs_0_mix_columns_1_n178,
         aes_state_regs_0_mix_columns_1_n177,
         aes_state_regs_0_mix_columns_1_n176,
         aes_state_regs_0_mix_columns_1_n175,
         aes_state_regs_0_mix_columns_1_n174,
         aes_state_regs_0_mix_columns_1_n173,
         aes_state_regs_0_mix_columns_1_n172,
         aes_state_regs_0_mix_columns_1_n171,
         aes_state_regs_0_mix_columns_1_n170,
         aes_state_regs_0_mix_columns_1_n169,
         aes_state_regs_0_mix_columns_1_n168,
         aes_state_regs_0_mix_columns_1_n167,
         aes_state_regs_0_mix_columns_1_n166,
         aes_state_regs_0_mix_columns_1_n165,
         aes_state_regs_0_mix_columns_1_n164,
         aes_state_regs_0_mix_columns_1_n163,
         aes_state_regs_0_mix_columns_1_n162,
         aes_state_regs_0_mix_columns_1_n161,
         aes_state_regs_0_mix_columns_1_n160,
         aes_state_regs_0_mix_columns_1_n159;
  wire   [15:0] KeyToSboxOutxD;
  wire   [15:0] KeyInxD;
  wire   [15:0] StateOutxD;
  wire   [15:0] StateInxD;
  wire   [15:0] KeyOutxD;
  wire   [15:0] K03xD;
  wire   [7:0] RCONxD;
  wire   [15:0] aes_sbox_InvUnmappedxD;
  wire   [7:0] aes_sbox_Y0mulY1xD;
  wire   [5:0] aes_sbox_Y0xorY1xD;
  wire   [7:0] aes_sbox_Y0xorY12xD;
  wire   [7:0] aes_sbox_Y1_4xDP;
  wire   [7:0] aes_sbox_Y1_3xDP;
  wire   [7:0] aes_sbox_Y1_2xDP;
  wire   [7:0] aes_sbox_Y1_1xDP;
  wire   [7:0] aes_sbox_Y1_0xDP;
  wire   [7:0] aes_sbox_Y0_4xDP;
  wire   [7:0] aes_sbox_Y0_3xDP;
  wire   [7:0] aes_sbox_Y0_2xDP;
  wire   [7:0] aes_sbox_Y0_1xDP;
  wire   [7:0] aes_sbox_Y0_0xDP;
  wire   [7:0] aes_sbox_InverterInxD;
  wire   [7:0] aes_sbox_InverterInxDP;
  wire   [15:0] aes_sbox_mul_y0y1_FFxDN;
  wire   [3:0] aes_sbox_inverter_gf24_AmulBxD;
  wire   [3:0] aes_sbox_inverter_gf24_ExD;
  wire   [3:0] aes_sbox_inverter_gf24_pipelinedBxDP;
  wire   [3:0] aes_sbox_inverter_gf24_pipelinedAxDP;
  wire   [3:0] aes_sbox_inverter_gf24_BxDP;
  wire   [3:0] aes_sbox_inverter_gf24_AxDP;
  wire   [7:0] aes_sbox_inverter_gf24_a_mul_b_FFxDN;
  wire   [7:0] aes_sbox_inverter_gf24_a_mul_e_FFxDN;
  wire   [7:0] aes_sbox_inverter_gf24_b_mul_e_FFxDN;
  wire   [15:0] aes_sbox_mult_msb_FFxDN;
  wire   [15:0] aes_sbox_mult_lsb_FFxDN;
  wire   [7:0] aes_key_regs_1_K23xDN;
  wire   [7:0] aes_key_regs_1_K22xDN;
  wire   [7:0] aes_key_regs_1_K21xDN;
  wire   [7:0] aes_key_regs_1_K20xDN;
  wire   [7:0] aes_key_regs_1_K13xDN;
  wire   [7:0] aes_key_regs_1_K12xDN;
  wire   [7:0] aes_key_regs_1_K11xDN;
  wire   [7:0] aes_key_regs_1_K10xDN;
  wire   [7:0] aes_key_regs_1_K02xDN;
  wire   [7:0] aes_key_regs_1_K01xDN;
  wire   [7:0] aes_key_regs_1_K00xDN;
  wire   [7:0] aes_state_regs_1_MixColumnsS3xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS2xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS1xD;
  wire   [7:0] aes_state_regs_1_MixColumnsS0xD;
  wire   [7:0] aes_state_regs_1_S20xDN;
  wire   [7:1] aes_state_regs_1_S21xDP;
  wire   [7:0] aes_state_regs_1_S10xDN;
  wire   [7:0] aes_state_regs_1_S03xDN;
  wire   [7:0] aes_state_regs_1_S02xDN;
  wire   [7:0] aes_state_regs_1_S01xDN;
  wire   [7:0] aes_state_regs_1_S00xDP;
  wire   [7:0] aes_key_regs_0_K23xDN;
  wire   [7:0] aes_key_regs_0_K22xDN;
  wire   [7:0] aes_key_regs_0_K21xDN;
  wire   [7:0] aes_key_regs_0_K20xDN;
  wire   [7:0] aes_key_regs_0_K13xDN;
  wire   [7:0] aes_key_regs_0_K12xDN;
  wire   [7:0] aes_key_regs_0_K11xDN;
  wire   [7:0] aes_key_regs_0_K10xDN;
  wire   [7:0] aes_key_regs_0_K02xDN;
  wire   [7:0] aes_key_regs_0_K01xDN;
  wire   [7:0] aes_key_regs_0_K00xDN;
  wire   [7:0] aes_state_regs_0_MixColumnsS3xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS2xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS1xD;
  wire   [7:0] aes_state_regs_0_MixColumnsS0xD;
  wire   [7:0] aes_state_regs_0_S20xDN;
  wire   [7:1] aes_state_regs_0_S21xDP;
  wire   [7:0] aes_state_regs_0_S10xDN;
  wire   [7:0] aes_state_regs_0_S03xDN;
  wire   [7:0] aes_state_regs_0_S02xDN;
  wire   [7:0] aes_state_regs_0_S01xDN;
  wire   [7:0] aes_state_regs_0_S00xDP;

  DFFR_X1 disableKeyRegsxSP_reg ( .D(n113), .CK(ClkxCI), .RN(RstxBI), .Q(), 
        .QN(n226) );
  OAI22_X1 U296 ( .A1(StateOutxD[5]), .A2(n338), .B1(PTxDI[5]), .B2(n337), 
        .ZN(n290) );
  OAI22_X1 U297 ( .A1(StateOutxD[13]), .A2(n338), .B1(PTxDI[13]), .B2(n337), 
        .ZN(n323) );
  OAI22_X1 U298 ( .A1(StateOutxD[14]), .A2(n338), .B1(PTxDI[14]), .B2(n337), 
        .ZN(n328) );
  NOR2_X1 U299 ( .A1(StateKEYSCHEDULExS), .A2(nextRCONxS), .ZN(n257) );
  OAI22_X1 U300 ( .A1(K03xD[13]), .A2(n334), .B1(StateInxD[13]), .B2(n333), 
        .ZN(n322) );
  AOI22_X1 U301 ( .A1(FinishedxS), .A2(KxDI[14]), .B1(KeyOutxD[14]), .B2(n326), 
        .ZN(n327) );
  OAI22_X1 U302 ( .A1(K03xD[14]), .A2(n334), .B1(StateInxD[14]), .B2(n333), 
        .ZN(n326) );
  INV_X1 U303 ( .A(n332), .ZN(n334) );
  NOR2_X1 U304 ( .A1(FinishedxS), .A2(n252), .ZN(n331) );
  INV_X1 U305 ( .A(StateKEYADDITION1o3xS), .ZN(n252) );
  INV_X1 U306 ( .A(n331), .ZN(n333) );
  INV_X1 U307 ( .A(n336), .ZN(n338) );
  NAND2_X2 U308 ( .A1(FinishedxS), .A2(n257), .ZN(n337) );
  INV_X1 U309 ( .A(n337), .ZN(n335) );
  OAI21_X1 U310 ( .B1(n264), .B2(KeyInxD[1]), .A(n263), .ZN(CxDO[1]) );
  AOI22_X1 U311 ( .A1(KeyToSboxOutxD[1]), .A2(n114), .B1(n262), .B2(KeyInxD[1]), .ZN(n263) );
  OAI22_X1 U312 ( .A1(StateOutxD[1]), .A2(n338), .B1(PTxDI[1]), .B2(n337), 
        .ZN(n262) );
  OAI21_X1 U313 ( .B1(n271), .B2(KeyInxD[2]), .A(n270), .ZN(CxDO[2]) );
  AOI22_X1 U314 ( .A1(n336), .A2(StateOutxD[2]), .B1(n335), .B2(PTxDI[2]), 
        .ZN(n271) );
  AOI22_X1 U315 ( .A1(KeyToSboxOutxD[2]), .A2(n114), .B1(n269), .B2(KeyInxD[2]), .ZN(n270) );
  OAI22_X1 U316 ( .A1(StateOutxD[2]), .A2(n338), .B1(PTxDI[2]), .B2(n337), 
        .ZN(n269) );
  OAI21_X1 U317 ( .B1(n278), .B2(KeyInxD[3]), .A(n277), .ZN(CxDO[3]) );
  AOI22_X1 U318 ( .A1(n336), .A2(StateOutxD[3]), .B1(n335), .B2(PTxDI[3]), 
        .ZN(n278) );
  AOI22_X1 U319 ( .A1(KeyToSboxOutxD[3]), .A2(n114), .B1(n276), .B2(KeyInxD[3]), .ZN(n277) );
  OAI22_X1 U320 ( .A1(StateOutxD[3]), .A2(n338), .B1(PTxDI[3]), .B2(n337), 
        .ZN(n276) );
  OAI21_X1 U321 ( .B1(n285), .B2(KeyInxD[4]), .A(n284), .ZN(CxDO[4]) );
  AOI22_X1 U322 ( .A1(KeyToSboxOutxD[4]), .A2(n114), .B1(n283), .B2(KeyInxD[4]), .ZN(n284) );
  OAI22_X1 U323 ( .A1(StateOutxD[4]), .A2(n338), .B1(PTxDI[4]), .B2(n337), 
        .ZN(n283) );
  OAI21_X1 U324 ( .B1(n292), .B2(KeyInxD[5]), .A(n291), .ZN(CxDO[5]) );
  AOI22_X1 U325 ( .A1(KeyToSboxOutxD[5]), .A2(n114), .B1(n290), .B2(KeyInxD[5]), .ZN(n291) );
  OAI21_X1 U326 ( .B1(n299), .B2(KeyInxD[6]), .A(n298), .ZN(CxDO[6]) );
  OAI22_X1 U327 ( .A1(StateOutxD[6]), .A2(n338), .B1(PTxDI[6]), .B2(n337), 
        .ZN(n297) );
  OAI21_X1 U328 ( .B1(n306), .B2(KeyInxD[7]), .A(n305), .ZN(CxDO[7]) );
  AOI22_X1 U329 ( .A1(KeyToSboxOutxD[7]), .A2(n114), .B1(n304), .B2(KeyInxD[7]), .ZN(n305) );
  OAI22_X1 U330 ( .A1(StateOutxD[7]), .A2(n338), .B1(PTxDI[7]), .B2(n337), 
        .ZN(n304) );
  OAI21_X1 U331 ( .B1(n312), .B2(KeyInxD[9]), .A(n311), .ZN(CxDO[9]) );
  AOI22_X1 U332 ( .A1(n336), .A2(StateOutxD[9]), .B1(n335), .B2(PTxDI[9]), 
        .ZN(n312) );
  AOI22_X1 U333 ( .A1(KeyToSboxOutxD[9]), .A2(n114), .B1(n310), .B2(KeyInxD[9]), .ZN(n311) );
  OAI22_X1 U334 ( .A1(StateOutxD[9]), .A2(n338), .B1(PTxDI[9]), .B2(n337), 
        .ZN(n310) );
  OAI21_X1 U335 ( .B1(n315), .B2(KeyInxD[10]), .A(n314), .ZN(CxDO[10]) );
  AOI22_X1 U336 ( .A1(n336), .A2(StateOutxD[10]), .B1(n335), .B2(PTxDI[10]), 
        .ZN(n315) );
  AOI22_X1 U337 ( .A1(KeyToSboxOutxD[10]), .A2(n114), .B1(n313), .B2(
        KeyInxD[10]), .ZN(n314) );
  OAI22_X1 U338 ( .A1(StateOutxD[10]), .A2(n338), .B1(PTxDI[10]), .B2(n337), 
        .ZN(n313) );
  OAI21_X1 U339 ( .B1(n318), .B2(KeyInxD[11]), .A(n317), .ZN(CxDO[11]) );
  AOI22_X1 U340 ( .A1(n336), .A2(StateOutxD[11]), .B1(n335), .B2(PTxDI[11]), 
        .ZN(n318) );
  AOI22_X1 U341 ( .A1(KeyToSboxOutxD[11]), .A2(n114), .B1(n316), .B2(
        KeyInxD[11]), .ZN(n317) );
  OAI22_X1 U342 ( .A1(StateOutxD[11]), .A2(n338), .B1(PTxDI[11]), .B2(n337), 
        .ZN(n316) );
  OAI21_X1 U343 ( .B1(n321), .B2(KeyInxD[12]), .A(n320), .ZN(CxDO[12]) );
  AOI22_X1 U344 ( .A1(n336), .A2(StateOutxD[12]), .B1(n335), .B2(PTxDI[12]), 
        .ZN(n321) );
  AOI22_X1 U345 ( .A1(KeyToSboxOutxD[12]), .A2(n114), .B1(n319), .B2(
        KeyInxD[12]), .ZN(n320) );
  OAI22_X1 U346 ( .A1(StateOutxD[12]), .A2(n338), .B1(PTxDI[12]), .B2(n337), 
        .ZN(n319) );
  OAI21_X1 U347 ( .B1(n325), .B2(KeyInxD[13]), .A(n324), .ZN(CxDO[13]) );
  AOI22_X1 U348 ( .A1(n336), .A2(StateOutxD[13]), .B1(n335), .B2(PTxDI[13]), 
        .ZN(n325) );
  AOI22_X1 U349 ( .A1(KeyToSboxOutxD[13]), .A2(n114), .B1(n323), .B2(
        KeyInxD[13]), .ZN(n324) );
  OAI21_X1 U350 ( .B1(n330), .B2(KeyInxD[14]), .A(n329), .ZN(CxDO[14]) );
  AOI22_X1 U351 ( .A1(n336), .A2(StateOutxD[14]), .B1(n335), .B2(PTxDI[14]), 
        .ZN(n330) );
  AOI22_X1 U352 ( .A1(KeyToSboxOutxD[14]), .A2(n114), .B1(n328), .B2(
        KeyInxD[14]), .ZN(n329) );
  OAI21_X1 U353 ( .B1(n341), .B2(KeyInxD[15]), .A(n340), .ZN(CxDO[15]) );
  AOI22_X1 U354 ( .A1(n336), .A2(StateOutxD[15]), .B1(n335), .B2(PTxDI[15]), 
        .ZN(n341) );
  AOI22_X1 U355 ( .A1(KeyToSboxOutxD[15]), .A2(n114), .B1(n339), .B2(
        KeyInxD[15]), .ZN(n340) );
  OAI22_X1 U356 ( .A1(StateOutxD[15]), .A2(n338), .B1(PTxDI[15]), .B2(n337), 
        .ZN(n339) );
  AND2_X1 U357 ( .A1(LastRoundxS), .A2(showRCONxS), .ZN(DonexSO) );
  OAI21_X1 U358 ( .B1(n333), .B2(n256), .A(n255), .ZN(KeyInxD[0]) );
  XNOR2_X1 U359 ( .A(StateInxD[0]), .B(n253), .ZN(n256) );
  AOI22_X1 U360 ( .A1(FinishedxS), .A2(KxDI[0]), .B1(n332), .B2(n254), .ZN(
        n255) );
  XOR2_X1 U361 ( .A(KeyOutxD[0]), .B(RCONxD[0]), .Z(n253) );
  XOR2_X1 U362 ( .A(KeyOutxD[0]), .B(K03xD[0]), .Z(n254) );
  OAI21_X1 U363 ( .B1(n333), .B2(n261), .A(n260), .ZN(KeyInxD[1]) );
  XNOR2_X1 U364 ( .A(StateInxD[1]), .B(n258), .ZN(n261) );
  AOI22_X1 U365 ( .A1(FinishedxS), .A2(KxDI[1]), .B1(n332), .B2(n259), .ZN(
        n260) );
  XOR2_X1 U366 ( .A(KeyOutxD[1]), .B(RCONxD[1]), .Z(n258) );
  XOR2_X1 U367 ( .A(KeyOutxD[1]), .B(K03xD[1]), .Z(n259) );
  OAI21_X1 U368 ( .B1(n333), .B2(n268), .A(n267), .ZN(KeyInxD[2]) );
  XNOR2_X1 U369 ( .A(StateInxD[2]), .B(n265), .ZN(n268) );
  AOI22_X1 U370 ( .A1(FinishedxS), .A2(KxDI[2]), .B1(n332), .B2(n266), .ZN(
        n267) );
  XOR2_X1 U371 ( .A(KeyOutxD[2]), .B(RCONxD[2]), .Z(n265) );
  XOR2_X1 U372 ( .A(KeyOutxD[2]), .B(K03xD[2]), .Z(n266) );
  OAI21_X1 U373 ( .B1(n333), .B2(n275), .A(n274), .ZN(KeyInxD[3]) );
  XNOR2_X1 U374 ( .A(StateInxD[3]), .B(n272), .ZN(n275) );
  AOI22_X1 U375 ( .A1(FinishedxS), .A2(KxDI[3]), .B1(n332), .B2(n273), .ZN(
        n274) );
  XOR2_X1 U376 ( .A(KeyOutxD[3]), .B(RCONxD[3]), .Z(n272) );
  XOR2_X1 U377 ( .A(KeyOutxD[3]), .B(K03xD[3]), .Z(n273) );
  OAI21_X1 U378 ( .B1(n333), .B2(n282), .A(n281), .ZN(KeyInxD[4]) );
  XNOR2_X1 U379 ( .A(StateInxD[4]), .B(n279), .ZN(n282) );
  AOI22_X1 U380 ( .A1(FinishedxS), .A2(KxDI[4]), .B1(n332), .B2(n280), .ZN(
        n281) );
  XOR2_X1 U381 ( .A(KeyOutxD[4]), .B(RCONxD[4]), .Z(n279) );
  XOR2_X1 U382 ( .A(KeyOutxD[4]), .B(K03xD[4]), .Z(n280) );
  OAI21_X1 U383 ( .B1(n333), .B2(n289), .A(n288), .ZN(KeyInxD[5]) );
  AOI22_X1 U384 ( .A1(FinishedxS), .A2(KxDI[5]), .B1(n332), .B2(n287), .ZN(
        n288) );
  XOR2_X1 U385 ( .A(KeyOutxD[5]), .B(RCONxD[5]), .Z(n286) );
  XOR2_X1 U386 ( .A(KeyOutxD[5]), .B(K03xD[5]), .Z(n287) );
  OAI21_X1 U387 ( .B1(n333), .B2(n296), .A(n295), .ZN(KeyInxD[6]) );
  XNOR2_X1 U388 ( .A(StateInxD[6]), .B(n293), .ZN(n296) );
  AOI22_X1 U389 ( .A1(FinishedxS), .A2(KxDI[6]), .B1(n332), .B2(n294), .ZN(
        n295) );
  XOR2_X1 U390 ( .A(KeyOutxD[6]), .B(RCONxD[6]), .Z(n293) );
  XOR2_X1 U391 ( .A(KeyOutxD[6]), .B(K03xD[6]), .Z(n294) );
  OAI21_X1 U392 ( .B1(n333), .B2(n303), .A(n302), .ZN(KeyInxD[7]) );
  XNOR2_X1 U393 ( .A(StateInxD[7]), .B(n300), .ZN(n303) );
  AOI22_X1 U394 ( .A1(FinishedxS), .A2(KxDI[7]), .B1(n332), .B2(n301), .ZN(
        n302) );
  XOR2_X1 U395 ( .A(KeyOutxD[7]), .B(RCONxD[7]), .Z(n300) );
  XOR2_X1 U396 ( .A(KeyOutxD[7]), .B(K03xD[7]), .Z(n301) );
  OAI21_X1 U397 ( .B1(KeyOutxD[8]), .B2(n309), .A(n308), .ZN(KeyInxD[8]) );
  AOI22_X1 U398 ( .A1(n332), .A2(K03xD[8]), .B1(n331), .B2(StateInxD[8]), .ZN(
        n309) );
  AOI22_X1 U399 ( .A1(FinishedxS), .A2(KxDI[8]), .B1(KeyOutxD[8]), .B2(n307), 
        .ZN(n308) );
  OAI22_X1 U400 ( .A1(K03xD[8]), .A2(n334), .B1(StateInxD[8]), .B2(n333), .ZN(
        n307) );
  AOI22_X1 U401 ( .A1(n331), .A2(StateInxD[9]), .B1(n332), .B2(K03xD[9]), .ZN(
        n227) );
  OAI22_X1 U402 ( .A1(n333), .A2(StateInxD[9]), .B1(n334), .B2(K03xD[9]), .ZN(
        n228) );
  AOI22_X1 U403 ( .A1(FinishedxS), .A2(KxDI[9]), .B1(KeyOutxD[9]), .B2(n228), 
        .ZN(n229) );
  OAI21_X1 U404 ( .B1(KeyOutxD[9]), .B2(n227), .A(n229), .ZN(KeyInxD[9]) );
  AOI22_X1 U405 ( .A1(n331), .A2(StateInxD[10]), .B1(n332), .B2(K03xD[10]), 
        .ZN(n230) );
  OAI22_X1 U406 ( .A1(n333), .A2(StateInxD[10]), .B1(n334), .B2(K03xD[10]), 
        .ZN(n231) );
  AOI22_X1 U407 ( .A1(FinishedxS), .A2(KxDI[10]), .B1(KeyOutxD[10]), .B2(n231), 
        .ZN(n232) );
  OAI21_X1 U408 ( .B1(KeyOutxD[10]), .B2(n230), .A(n232), .ZN(KeyInxD[10]) );
  AOI22_X1 U409 ( .A1(n331), .A2(StateInxD[11]), .B1(n332), .B2(K03xD[11]), 
        .ZN(n233) );
  OAI22_X1 U410 ( .A1(n333), .A2(StateInxD[11]), .B1(n334), .B2(K03xD[11]), 
        .ZN(n234) );
  AOI22_X1 U411 ( .A1(FinishedxS), .A2(KxDI[11]), .B1(KeyOutxD[11]), .B2(n234), 
        .ZN(n235) );
  OAI21_X1 U412 ( .B1(KeyOutxD[11]), .B2(n233), .A(n235), .ZN(KeyInxD[11]) );
  AOI22_X1 U413 ( .A1(n331), .A2(StateInxD[12]), .B1(n332), .B2(K03xD[12]), 
        .ZN(n236) );
  OAI22_X1 U414 ( .A1(n333), .A2(StateInxD[12]), .B1(n334), .B2(K03xD[12]), 
        .ZN(n237) );
  AOI22_X1 U415 ( .A1(FinishedxS), .A2(KxDI[12]), .B1(KeyOutxD[12]), .B2(n237), 
        .ZN(n238) );
  OAI21_X1 U416 ( .B1(KeyOutxD[12]), .B2(n236), .A(n238), .ZN(KeyInxD[12]) );
  AOI22_X1 U417 ( .A1(K03xD[13]), .A2(n332), .B1(StateInxD[13]), .B2(n331), 
        .ZN(n239) );
  AOI22_X1 U418 ( .A1(FinishedxS), .A2(KxDI[13]), .B1(KeyOutxD[13]), .B2(n322), 
        .ZN(n240) );
  OAI21_X1 U419 ( .B1(KeyOutxD[13]), .B2(n239), .A(n240), .ZN(KeyInxD[13]) );
  AOI22_X1 U420 ( .A1(n331), .A2(StateInxD[15]), .B1(n332), .B2(K03xD[15]), 
        .ZN(n241) );
  OAI22_X1 U421 ( .A1(n333), .A2(StateInxD[15]), .B1(n334), .B2(K03xD[15]), 
        .ZN(n242) );
  AOI22_X1 U422 ( .A1(FinishedxS), .A2(KxDI[15]), .B1(KeyOutxD[15]), .B2(n242), 
        .ZN(n243) );
  OAI21_X1 U423 ( .B1(KeyOutxD[15]), .B2(n241), .A(n243), .ZN(KeyInxD[15]) );
  AOI22_X1 U424 ( .A1(n336), .A2(StateOutxD[0]), .B1(n335), .B2(PTxDI[0]), 
        .ZN(n244) );
  OAI22_X1 U425 ( .A1(n337), .A2(PTxDI[0]), .B1(n338), .B2(StateOutxD[0]), 
        .ZN(n245) );
  AOI22_X1 U426 ( .A1(n114), .A2(KeyToSboxOutxD[0]), .B1(KeyInxD[0]), .B2(n245), .ZN(n246) );
  OAI21_X1 U427 ( .B1(KeyInxD[0]), .B2(n244), .A(n246), .ZN(CxDO[0]) );
  INV_X1 U428 ( .A(ClkxCI), .ZN(n251) );
  AOI22_X1 U429 ( .A1(n336), .A2(StateOutxD[8]), .B1(n335), .B2(PTxDI[8]), 
        .ZN(n247) );
  OAI22_X1 U430 ( .A1(n337), .A2(PTxDI[8]), .B1(n338), .B2(StateOutxD[8]), 
        .ZN(n248) );
  AOI22_X1 U431 ( .A1(n114), .A2(KeyToSboxOutxD[8]), .B1(KeyInxD[8]), .B2(n248), .ZN(n249) );
  OAI21_X1 U432 ( .B1(KeyInxD[8]), .B2(n247), .A(n249), .ZN(CxDO[8]) );
  AOI22_X1 U433 ( .A1(n331), .A2(StateInxD[14]), .B1(K03xD[14]), .B2(n332), 
        .ZN(n250) );
  OAI21_X1 U434 ( .B1(KeyOutxD[14]), .B2(n250), .A(n327), .ZN(KeyInxD[14]) );
  INV_X1 U435 ( .A(disableKeyRegsxS), .ZN(n113) );
  NOR2_X4 U436 ( .A1(FinishedxS), .A2(n114), .ZN(n336) );
  INV_X4 U437 ( .A(n257), .ZN(n114) );
  NOR2_X4 U438 ( .A1(FinishedxS), .A2(StateKEYADDITION1o3xS), .ZN(n332) );
  NOR2_X1 U439 ( .A1(n226), .A2(n251), .ZN(ClkKeyRegxC) );
  AOI22_X1 U440 ( .A1(n336), .A2(StateOutxD[1]), .B1(n335), .B2(PTxDI[1]), 
        .ZN(n264) );
  AOI22_X1 U441 ( .A1(n336), .A2(StateOutxD[4]), .B1(n335), .B2(PTxDI[4]), 
        .ZN(n285) );
  XNOR2_X1 U442 ( .A(StateInxD[5]), .B(n286), .ZN(n289) );
  AOI22_X1 U443 ( .A1(n336), .A2(StateOutxD[5]), .B1(n335), .B2(PTxDI[5]), 
        .ZN(n292) );
  AOI22_X1 U444 ( .A1(n336), .A2(StateOutxD[6]), .B1(n335), .B2(PTxDI[6]), 
        .ZN(n299) );
  AOI22_X1 U445 ( .A1(KeyToSboxOutxD[6]), .A2(n114), .B1(n297), .B2(KeyInxD[6]), .ZN(n298) );
  AOI22_X1 U446 ( .A1(n336), .A2(StateOutxD[7]), .B1(n335), .B2(PTxDI[7]), 
        .ZN(n306) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U31 ( .A1(aes_ctrl_lsfr_23_cycles_1_n23), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n17), .ZN(nextRCONxS) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U30 ( .A1(aes_ctrl_lsfr_23_cycles_1_n6), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n17), .ZN(disableKeyRegsxS) );
  OAI22_X1 aes_ctrl_lsfr_23_cycles_1_U29 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n23), .B1(aes_ctrl_lsfr_23_cycles_1_n3), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n24), .ZN(aes_ctrl_lsfr_23_cycles_1_n39)
         );
  AOI221_X1 aes_ctrl_lsfr_23_cycles_1_U28 ( .B1(StartxSI), .B2(
        aes_ctrl_lsfr_23_cycles_1_n22), .C1(aes_ctrl_lsfr_23_cycles_1_n21), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n22), .A(aes_ctrl_lsfr_23_cycles_1_n8), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n3) );
  XNOR2_X1 aes_ctrl_lsfr_23_cycles_1_U27 ( .A(aes_ctrl_lsfr_23_cycles_1_n1), 
        .B(aes_ctrl_lsfr_23_cycles_1_n5), .ZN(aes_ctrl_lsfr_23_cycles_1_n36)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U26 ( .A1(aes_ctrl_lsfr_23_cycles_1_n22), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n19), .ZN(aes_ctrl_lsfr_23_cycles_1_n1)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U25 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_N16)
         );
  AOI211_X1 aes_ctrl_lsfr_23_cycles_1_U24 ( .C1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n11), .A(aes_ctrl_lsfr_23_cycles_1_n13), 
        .B(aes_ctrl_lsfr_23_cycles_1_n7), .ZN(aes_ctrl_lsfr_23_cycles_1_N66)
         );
  OAI22_X1 aes_ctrl_lsfr_23_cycles_1_U23 ( .A1(aes_ctrl_lsfr_23_cycles_1_n7), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n15), .B1(aes_ctrl_lsfr_23_cycles_1_n17), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_N83)
         );
  AOI22_X1 aes_ctrl_lsfr_23_cycles_1_U22 ( .A1(aes_ctrl_lsfr_23_cycles_1_n20), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .B1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n23), .ZN(aes_ctrl_lsfr_23_cycles_1_n37)
         );
  OAI221_X1 aes_ctrl_lsfr_23_cycles_1_U21 ( .B1(aes_ctrl_lsfr_23_cycles_1_n20), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n4), .C1(aes_ctrl_lsfr_23_cycles_1_n23), 
        .C2(aes_ctrl_lsfr_23_cycles_1_n18), .A(aes_ctrl_lsfr_23_cycles_1_n22), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n35) );
  XNOR2_X1 aes_ctrl_lsfr_23_cycles_1_U20 ( .A(aes_ctrl_lsfr_23_cycles_1_n24), 
        .B(aes_ctrl_lsfr_23_cycles_1_n9), .ZN(aes_ctrl_lsfr_23_cycles_1_n38)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U19 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .ZN(aes_ctrl_lsfr_23_cycles_1_n18)
         );
  NAND3_X1 aes_ctrl_lsfr_23_cycles_1_U18 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n9), .A3(aes_ctrl_lsfr_23_cycles_1_n6), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n14) );
  OAI21_X1 aes_ctrl_lsfr_23_cycles_1_U17 ( .B1(aes_ctrl_lsfr_23_cycles_1_n10), 
        .B2(aes_ctrl_lsfr_23_cycles_1_n8), .A(aes_ctrl_lsfr_23_cycles_1_n5), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n11) );
  NOR2_X2 aes_ctrl_lsfr_23_cycles_1_U16 ( .A1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n11), .ZN(aes_ctrl_lsfr_23_cycles_1_n13)
         );
  INV_X1 aes_ctrl_lsfr_23_cycles_1_U15 ( .A(aes_ctrl_lsfr_23_cycles_1_n13), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n15) );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U14 ( .A1(aes_ctrl_lsfr_23_cycles_1_n4), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n7), .ZN(aes_ctrl_lsfr_23_cycles_1_n17)
         );
  AND2_X1 aes_ctrl_lsfr_23_cycles_1_U13 ( .A1(aes_ctrl_lsfr_23_cycles_1_n8), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n22), .ZN(aes_ctrl_lsfr_23_cycles_1_n24)
         );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U12 ( .A1(aes_ctrl_lsfr_23_cycles_1_n19), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n5), .ZN(aes_ctrl_lsfr_23_cycles_1_n23)
         );
  OR2_X1 aes_ctrl_lsfr_23_cycles_1_U11 ( .A1(aes_ctrl_lsfr_23_cycles_1_n2), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n4), .ZN(aes_ctrl_lsfr_23_cycles_1_n22)
         );
  OR3_X1 aes_ctrl_lsfr_23_cycles_1_U10 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n10), .A3(aes_ctrl_lsfr_23_cycles_1_n5), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n21) );
  INV_X1 aes_ctrl_lsfr_23_cycles_1_U9 ( .A(aes_ctrl_lsfr_23_cycles_1_n23), 
        .ZN(aes_ctrl_lsfr_23_cycles_1_n20) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U8 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n9), .ZN(aes_ctrl_lsfr_23_cycles_1_n19)
         );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U7 ( .A1(aes_ctrl_lsfr_23_cycles_1_n17), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n16), .ZN(StateKEYSCHEDULExS) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U6 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n21), .ZN(showRCONxS) );
  NOR4_X1 aes_ctrl_lsfr_23_cycles_1_U5 ( .A1(aes_ctrl_lsfr_23_cycles_1_n12), 
        .A2(LastRoundxS), .A3(aes_ctrl_lsfr_23_cycles_1_n7), .A4(
        aes_ctrl_lsfr_23_cycles_1_n10), .ZN(doMixColumnsxS) );
  NOR2_X1 aes_ctrl_lsfr_23_cycles_1_U4 ( .A1(aes_ctrl_lsfr_23_cycles_1_n18), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n16), .ZN(StateKEYADDITION1o3xS) );
  NAND2_X1 aes_ctrl_lsfr_23_cycles_1_U3 ( .A1(aes_ctrl_lsfr_23_cycles_1_n11), 
        .A2(aes_ctrl_lsfr_23_cycles_1_n14), .ZN(aes_ctrl_lsfr_23_cycles_1_n16)
         );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_2_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n36), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n5), .QN(aes_ctrl_lsfr_23_cycles_1_n6) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_1_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n38), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n10), .QN(aes_ctrl_lsfr_23_cycles_1_n9) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_3_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n35), .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(
        aes_ctrl_lsfr_23_cycles_1_n4) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_4_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n37), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n7), .QN(aes_ctrl_lsfr_23_cycles_1_n2) );
  DFFR_X1 aes_ctrl_lsfr_23_cycles_1_LSFRxDP_reg_0_ ( .D(
        aes_ctrl_lsfr_23_cycles_1_n39), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_ctrl_lsfr_23_cycles_1_n8), .QN(aes_ctrl_lsfr_23_cycles_1_n12) );
  INV_X1 rcon_1_U37 ( .A(nextRCONxS), .ZN(rcon_1_n39) );
  AOI211_X1 rcon_1_U36 ( .C1(rcon_1_n9), .C2(rcon_1_n28), .A(rcon_1_n43), .B(
        rcon_1_n29), .ZN(rcon_1_n22) );
  OAI22_X1 rcon_1_U35 ( .A1(rcon_1_n38), .A2(rcon_1_n4), .B1(rcon_1_n9), .B2(
        rcon_1_n42), .ZN(rcon_1_n29) );
  INV_X1 rcon_1_U34 ( .A(rcon_1_n44), .ZN(rcon_1_n28) );
  INV_X1 rcon_1_U32 ( .A(rcon_1_n38), .ZN(rcon_1_n16) );
  INV_X1 rcon_1_U31 ( .A(rcon_1_n35), .ZN(rcon_1_n15) );
  OAI211_X1 rcon_1_U30 ( .C1(rcon_1_n38), .C2(rcon_1_n17), .A(rcon_1_n44), .B(
        rcon_1_n14), .ZN(rcon_1_n25) );
  INV_X1 rcon_1_U29 ( .A(rcon_1_n43), .ZN(rcon_1_n14) );
  AOI211_X1 rcon_1_U28 ( .C1(rcon_1_n39), .C2(rcon_1_n34), .A(rcon_1_n43), .B(
        rcon_1_n13), .ZN(rcon_1_n24) );
  AOI22_X1 rcon_1_U27 ( .A1(rcon_1_n37), .A2(rcon_1_n44), .B1(rcon_1_n42), 
        .B2(rcon_1_n17), .ZN(rcon_1_n13) );
  OAI21_X1 rcon_1_U26 ( .B1(rcon_1_n38), .B2(rcon_1_n33), .A(rcon_1_n12), .ZN(
        rcon_1_n21) );
  OAI211_X1 rcon_1_U25 ( .C1(rcon_1_n35), .C2(rcon_1_n4), .A(rcon_1_n38), .B(
        rcon_1_n11), .ZN(rcon_1_n12) );
  OAI21_X1 rcon_1_U24 ( .B1(rcon_1_n35), .B2(rcon_1_n36), .A(rcon_1_n4), .ZN(
        rcon_1_n11) );
  OAI22_X1 rcon_1_U23 ( .A1(rcon_1_n26), .A2(rcon_1_n38), .B1(rcon_1_n30), 
        .B2(rcon_1_n41), .ZN(rcon_1_n19) );
  OAI22_X1 rcon_1_U22 ( .A1(rcon_1_n38), .A2(rcon_1_n30), .B1(rcon_1_n33), 
        .B2(rcon_1_n41), .ZN(rcon_1_n20) );
  OAI22_X1 rcon_1_U21 ( .A1(rcon_1_n38), .A2(rcon_1_n31), .B1(rcon_1_n34), 
        .B2(rcon_1_n41), .ZN(rcon_1_n23) );
  NOR2_X1 rcon_1_U20 ( .A1(rcon_1_n32), .A2(rcon_1_n40), .ZN(RCONxD[7]) );
  NOR2_X1 rcon_1_U19 ( .A1(rcon_1_n26), .A2(rcon_1_n40), .ZN(RCONxD[6]) );
  NOR2_X1 rcon_1_U18 ( .A1(rcon_1_n30), .A2(rcon_1_n40), .ZN(RCONxD[5]) );
  NOR2_X1 rcon_1_U17 ( .A1(rcon_1_n33), .A2(rcon_1_n40), .ZN(RCONxD[4]) );
  AND2_X1 rcon_1_U16 ( .A1(rcon_1_n4), .A2(showRCONxS), .ZN(RCONxD[3]) );
  NOR2_X1 rcon_1_U15 ( .A1(rcon_1_n31), .A2(rcon_1_n40), .ZN(RCONxD[2]) );
  NOR2_X1 rcon_1_U14 ( .A1(rcon_1_n34), .A2(rcon_1_n40), .ZN(RCONxD[1]) );
  NOR2_X1 rcon_1_U13 ( .A1(rcon_1_n17), .A2(rcon_1_n40), .ZN(RCONxD[0]) );
  NAND2_X1 rcon_1_U12 ( .A1(rcon_1_n38), .A2(rcon_1_n45), .ZN(rcon_1_n41) );
  INV_X1 rcon_1_U11 ( .A(rcon_1_n39), .ZN(rcon_1_n38) );
  NOR2_X1 rcon_1_U10 ( .A1(rcon_1_n45), .A2(rcon_1_n39), .ZN(rcon_1_n43) );
  NAND2_X1 rcon_1_U9 ( .A1(rcon_1_n38), .A2(rcon_1_n35), .ZN(rcon_1_n44) );
  NAND2_X1 rcon_1_U8 ( .A1(rcon_1_n38), .A2(rcon_1_n32), .ZN(rcon_1_n42) );
  INV_X2 rcon_1_U7 ( .A(rcon_1_n45), .ZN(FinishedxS) );
  INV_X1 rcon_1_U6 ( .A(showRCONxS), .ZN(rcon_1_n40) );
  NOR2_X1 rcon_1_U5 ( .A1(rcon_1_n30), .A2(rcon_1_n31), .ZN(LastRoundxS) );
  NAND2_X1 rcon_1_U4 ( .A1(rcon_1_n36), .A2(rcon_1_n4), .ZN(rcon_1_n45) );
  OAI33_X1 rcon_1_U3 ( .A1(1'b0), .A2(rcon_1_n38), .A3(rcon_1_n15), .B1(
        rcon_1_n16), .B2(rcon_1_n26), .B3(rcon_1_n4), .ZN(rcon_1_n18) );
  DFFR_X1 rcon_1_RCONxDP_reg_4_ ( .D(rcon_1_n21), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(rcon_1_n33) );
  DFFR_X1 rcon_1_RCONxDP_reg_1_ ( .D(rcon_1_n24), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(rcon_1_n34) );
  DFFR_X1 rcon_1_RCONxDP_reg_0_ ( .D(rcon_1_n25), .CK(ClkxCI), .RN(RstxBI), 
        .Q(rcon_1_n37), .QN(rcon_1_n17) );
  DFFR_X1 rcon_1_RCONxDP_reg_7_ ( .D(rcon_1_n18), .CK(ClkxCI), .RN(RstxBI), 
        .Q(rcon_1_n35), .QN(rcon_1_n32) );
  DFFS_X1 rcon_1_RCONxDP_reg_3_ ( .D(rcon_1_n22), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n4), .QN() );
  DFFS_X1 rcon_1_RCONxDP_reg_2_ ( .D(rcon_1_n23), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n9), .QN(rcon_1_n31) );
  DFFS_X1 rcon_1_RCONxDP_reg_5_ ( .D(rcon_1_n20), .CK(ClkxCI), .SN(RstxBI), 
        .Q(), .QN(rcon_1_n30) );
  DFFS_X1 rcon_1_RCONxDP_reg_6_ ( .D(rcon_1_n19), .CK(ClkxCI), .SN(RstxBI), 
        .Q(rcon_1_n36), .QN(rcon_1_n26) );
  MUX2_X1 aes_sbox_U30 ( .A(aes_sbox_n6), .B(aes_sbox_Y0xorY12xD[6]), .S(
        RstxBI), .Z(aes_sbox_n39) );
  MUX2_X1 aes_sbox_U29 ( .A(aes_sbox_n8), .B(aes_sbox_Y0xorY12xD[4]), .S(
        RstxBI), .Z(aes_sbox_n37) );
  MUX2_X1 aes_sbox_U28 ( .A(aes_sbox_n28), .B(aes_sbox_Y0xorY12xD[0]), .S(
        RstxBI), .Z(aes_sbox_n33) );
  XOR2_X1 aes_sbox_U27 ( .A(aes_sbox_n23), .B(aes_sbox_n24), .Z(
        aes_sbox_Y0xorY1xD[5]) );
  XOR2_X1 aes_sbox_U26 ( .A(aes_sbox_n19), .B(aes_sbox_n20), .Z(
        aes_sbox_Y0xorY1xD[3]) );
  XOR2_X1 aes_sbox_U25 ( .A(aes_sbox_n17), .B(aes_sbox_n18), .Z(
        aes_sbox_Y0xorY12xD[4]) );
  XOR2_X1 aes_sbox_U24 ( .A(aes_sbox_n11), .B(aes_sbox_n12), .Z(
        aes_sbox_Y0xorY1xD[0]) );
  XOR2_X1 aes_sbox_U23 ( .A(aes_sbox_n10), .B(aes_sbox_n9), .Z(
        aes_sbox_Y0xorY12xD[0]) );
  XOR2_X1 aes_sbox_U22 ( .A(aes_sbox_n5), .B(aes_sbox_Y0mulY1xD[7]), .Z(
        aes_sbox_InverterInxD[7]) );
  XOR2_X1 aes_sbox_U21 ( .A(aes_sbox_n6), .B(aes_sbox_Y0mulY1xD[6]), .Z(
        aes_sbox_InverterInxD[6]) );
  XOR2_X1 aes_sbox_U20 ( .A(aes_sbox_n7), .B(aes_sbox_Y0mulY1xD[5]), .Z(
        aes_sbox_InverterInxD[5]) );
  XOR2_X1 aes_sbox_U19 ( .A(aes_sbox_n8), .B(aes_sbox_Y0mulY1xD[4]), .Z(
        aes_sbox_InverterInxD[4]) );
  XOR2_X1 aes_sbox_U18 ( .A(aes_sbox_n25), .B(aes_sbox_Y0mulY1xD[3]), .Z(
        aes_sbox_InverterInxD[3]) );
  XOR2_X1 aes_sbox_U17 ( .A(aes_sbox_n26), .B(aes_sbox_Y0mulY1xD[2]), .Z(
        aes_sbox_InverterInxD[2]) );
  XOR2_X1 aes_sbox_U16 ( .A(aes_sbox_n27), .B(aes_sbox_Y0mulY1xD[1]), .Z(
        aes_sbox_InverterInxD[1]) );
  XOR2_X1 aes_sbox_U15 ( .A(aes_sbox_n28), .B(aes_sbox_Y0mulY1xD[0]), .Z(
        aes_sbox_InverterInxD[0]) );
  MUX2_X1 aes_sbox_U14 ( .A(aes_sbox_n7), .B(aes_sbox_Y0xorY12xD[5]), .S(
        RstxBI), .Z(aes_sbox_n38) );
  MUX2_X1 aes_sbox_U13 ( .A(aes_sbox_n27), .B(aes_sbox_Y0xorY12xD[1]), .S(
        RstxBI), .Z(aes_sbox_n34) );
  INV_X1 aes_sbox_U12 ( .A(aes_sbox_InvMappedxD_0__0_), .ZN(StateInxD[0]) );
  INV_X1 aes_sbox_U11 ( .A(aes_sbox_InvMappedxD_0__6_), .ZN(StateInxD[6]) );
  XOR2_X1 aes_sbox_U10 ( .A(aes_sbox_n15), .B(aes_sbox_n16), .Z(
        aes_sbox_Y0xorY1xD[2]) );
  MUX2_X1 aes_sbox_U9 ( .A(aes_sbox_n26), .B(aes_sbox_Y0xorY12xD[2]), .S(
        RstxBI), .Z(aes_sbox_n35) );
  INV_X1 aes_sbox_U8 ( .A(aes_sbox_InvMappedxD_0__1_), .ZN(StateInxD[1]) );
  XOR2_X1 aes_sbox_U7 ( .A(aes_sbox_n21), .B(aes_sbox_n22), .Z(
        aes_sbox_Y0xorY1xD[4]) );
  MUX2_X1 aes_sbox_U6 ( .A(aes_sbox_n5), .B(aes_sbox_Y0xorY12xD[7]), .S(RstxBI), .Z(aes_sbox_n40) );
  XOR2_X1 aes_sbox_U5 ( .A(aes_sbox_n13), .B(aes_sbox_n14), .Z(
        aes_sbox_Y0xorY1xD[1]) );
  MUX2_X1 aes_sbox_U4 ( .A(aes_sbox_n25), .B(aes_sbox_Y0xorY12xD[3]), .S(
        RstxBI), .Z(aes_sbox_n36) );
  INV_X1 aes_sbox_U3 ( .A(aes_sbox_InvMappedxD_0__5_), .ZN(StateInxD[5]) );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_0__0_ ( .D(aes_sbox_Y1_3xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_0__0_ ( .D(aes_sbox_Y1_2xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_0__1_ ( .D(aes_sbox_Y1_3xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_0__1_ ( .D(aes_sbox_Y1_2xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_0__2_ ( .D(aes_sbox_Y1_3xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_0__2_ ( .D(aes_sbox_Y1_2xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_0__3_ ( .D(aes_sbox_Y1_3xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_0__3_ ( .D(aes_sbox_Y1_2xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_1__0_ ( .D(aes_sbox_Y1_3xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_1__0_ ( .D(aes_sbox_Y1_2xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_1__1_ ( .D(aes_sbox_Y1_3xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_1__1_ ( .D(aes_sbox_Y1_2xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_1__2_ ( .D(aes_sbox_Y1_3xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_1__2_ ( .D(aes_sbox_Y1_2xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y1_4xDP_reg_1__3_ ( .D(aes_sbox_Y1_3xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_4xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y1_3xDP_reg_1__3_ ( .D(aes_sbox_Y1_2xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_3xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_0__0_ ( .D(aes_sbox_Y1_1xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_0__1_ ( .D(aes_sbox_Y1_1xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_0__2_ ( .D(aes_sbox_Y1_1xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_0__3_ ( .D(aes_sbox_Y1_1xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_1__0_ ( .D(aes_sbox_Y1_1xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_1__1_ ( .D(aes_sbox_Y1_1xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_1__2_ ( .D(aes_sbox_Y1_1xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y1_2xDP_reg_1__3_ ( .D(aes_sbox_Y1_1xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_2xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_0__0_ ( .D(aes_sbox_Y1_0xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_0__1_ ( .D(aes_sbox_Y1_0xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_0__2_ ( .D(aes_sbox_Y1_0xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_0__3_ ( .D(aes_sbox_Y1_0xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_1__0_ ( .D(aes_sbox_Y1_0xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_1__1_ ( .D(aes_sbox_Y1_0xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_1__2_ ( .D(aes_sbox_Y1_0xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y1_1xDP_reg_1__3_ ( .D(aes_sbox_Y1_0xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_1xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_0__0_ ( .D(aes_sbox_Y1xD_0__0_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_0__1_ ( .D(aes_sbox_Y1xD_0__1_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_0__2_ ( .D(aes_sbox_Y1xD_0__2_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_0__3_ ( .D(aes_sbox_Y1xD_0__3_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_1__0_ ( .D(aes_sbox_Y1xD_1__0_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_1__1_ ( .D(aes_sbox_Y1xD_1__1_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_1__2_ ( .D(aes_sbox_Y1xD_1__2_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y1_0xDP_reg_1__3_ ( .D(aes_sbox_Y1xD_1__3_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y1_0xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_0__0_ ( .D(aes_sbox_Y0_3xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_0__1_ ( .D(aes_sbox_Y0_3xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_0__2_ ( .D(aes_sbox_Y0_3xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_0__3_ ( .D(aes_sbox_Y0_3xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_1__0_ ( .D(aes_sbox_Y0_3xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_1__1_ ( .D(aes_sbox_Y0_3xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_1__2_ ( .D(aes_sbox_Y0_3xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y0_4xDP_reg_1__3_ ( .D(aes_sbox_Y0_3xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_4xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_0__0_ ( .D(aes_sbox_Y0_2xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_0__1_ ( .D(aes_sbox_Y0_2xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_0__2_ ( .D(aes_sbox_Y0_2xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_0__3_ ( .D(aes_sbox_Y0_2xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_1__0_ ( .D(aes_sbox_Y0_2xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_1__1_ ( .D(aes_sbox_Y0_2xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_1__2_ ( .D(aes_sbox_Y0_2xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y0_3xDP_reg_1__3_ ( .D(aes_sbox_Y0_2xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_3xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_0__0_ ( .D(aes_sbox_Y0_1xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_0__1_ ( .D(aes_sbox_Y0_1xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_0__2_ ( .D(aes_sbox_Y0_1xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_0__3_ ( .D(aes_sbox_Y0_1xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_1__0_ ( .D(aes_sbox_Y0_1xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_1__1_ ( .D(aes_sbox_Y0_1xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_1__2_ ( .D(aes_sbox_Y0_1xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y0_2xDP_reg_1__3_ ( .D(aes_sbox_Y0_1xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_2xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_0__0_ ( .D(aes_sbox_Y0_0xDP[0]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_0__1_ ( .D(aes_sbox_Y0_0xDP[1]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_0__2_ ( .D(aes_sbox_Y0_0xDP[2]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_0__3_ ( .D(aes_sbox_Y0_0xDP[3]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_1__0_ ( .D(aes_sbox_Y0_0xDP[4]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_1__1_ ( .D(aes_sbox_Y0_0xDP[5]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_1__2_ ( .D(aes_sbox_Y0_0xDP[6]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y0_1xDP_reg_1__3_ ( .D(aes_sbox_Y0_0xDP[7]), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_1xDP[7]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_0__0_ ( .D(aes_sbox_Y0xD_0__0_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[0]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_0__1_ ( .D(aes_sbox_Y0xD_0__1_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[1]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_0__2_ ( .D(aes_sbox_Y0xD_0__2_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[2]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_0__3_ ( .D(aes_sbox_Y0xD_0__3_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[3]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_1__0_ ( .D(aes_sbox_Y0xD_1__0_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[4]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_1__1_ ( .D(aes_sbox_Y0xD_1__1_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[5]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_1__2_ ( .D(aes_sbox_Y0xD_1__2_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[6]), .QN() );
  DFFR_X1 aes_sbox_Y0_0xDP_reg_1__3_ ( .D(aes_sbox_Y0xD_1__3_), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_sbox_Y0_0xDP[7]), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_0__0_ ( .D(aes_sbox_InverterInxD[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[0]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_0__0_ ( .D(aes_sbox_n33), .CK(ClkxCI), .Q(
        aes_sbox_n28), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_0__1_ ( .D(aes_sbox_InverterInxD[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[1]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_0__1_ ( .D(aes_sbox_n34), .CK(ClkxCI), .Q(
        aes_sbox_n27), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_0__2_ ( .D(aes_sbox_InverterInxD[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[2]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_0__2_ ( .D(aes_sbox_n35), .CK(ClkxCI), .Q(
        aes_sbox_n26), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_0__3_ ( .D(aes_sbox_InverterInxD[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[3]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_0__3_ ( .D(aes_sbox_n36), .CK(ClkxCI), .Q(
        aes_sbox_n25), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_1__0_ ( .D(aes_sbox_InverterInxD[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[4]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_1__0_ ( .D(aes_sbox_n37), .CK(ClkxCI), .Q(
        aes_sbox_n8), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_1__1_ ( .D(aes_sbox_InverterInxD[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[5]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_1__1_ ( .D(aes_sbox_n38), .CK(ClkxCI), .Q(
        aes_sbox_n7), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_1__2_ ( .D(aes_sbox_InverterInxD[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[6]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_1__2_ ( .D(aes_sbox_n39), .CK(ClkxCI), .Q(
        aes_sbox_n6), .QN() );
  DFFR_X1 aes_sbox_InverterInxDP_reg_1__3_ ( .D(aes_sbox_InverterInxD[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_InverterInxDP[7]), .QN() );
  DFF_X1 aes_sbox_Y0xorY12xDP_reg_1__3_ ( .D(aes_sbox_n40), .CK(ClkxCI), .Q(
        aes_sbox_n5), .QN() );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__0_ ( .D(aes_sbox_mappedxD_0__0_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y0xD_0__0_), .QN(aes_sbox_n9) );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__1_ ( .D(aes_sbox_mappedxD_0__1_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y0xD_0__1_), .QN(aes_sbox_n11) );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__2_ ( .D(CxDO[0]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(aes_sbox_Y0xD_0__2_), .QN(aes_sbox_n13) );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__3_ ( .D(aes_sbox_mappedxD_0__3_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y0xD_0__3_), .QN(aes_sbox_n15) );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__4_ ( .D(aes_sbox_mappedxD_0__4_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_0__0_), .QN(aes_sbox_n10) );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__5_ ( .D(aes_sbox_mappedxD_0__5_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_0__1_), .QN(aes_sbox_n12) );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__6_ ( .D(aes_sbox_mappedxD_0__6_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_0__2_), .QN(aes_sbox_n14) );
  DFFR_X1 aes_sbox_mappedxDP_reg_0__7_ ( .D(aes_sbox_mappedxD_0__7_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_0__3_), .QN(aes_sbox_n16) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__0_ ( .D(aes_sbox_mappedxD_1__0_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y0xD_1__0_), .QN(aes_sbox_n17) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__1_ ( .D(aes_sbox_mappedxD_1__1_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y0xD_1__1_), .QN(aes_sbox_n19) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__2_ ( .D(CxDO[8]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(aes_sbox_Y0xD_1__2_), .QN(aes_sbox_n21) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__3_ ( .D(aes_sbox_mappedxD_1__3_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y0xD_1__3_), .QN(aes_sbox_n23) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__4_ ( .D(aes_sbox_mappedxD_1__4_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_1__0_), .QN(aes_sbox_n18) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__5_ ( .D(aes_sbox_mappedxD_1__5_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_1__1_), .QN(aes_sbox_n20) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__6_ ( .D(aes_sbox_mappedxD_1__6_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_1__2_), .QN(aes_sbox_n22) );
  DFFR_X1 aes_sbox_mappedxDP_reg_1__7_ ( .D(aes_sbox_mappedxD_1__7_), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_sbox_Y1xD_1__3_), .QN(aes_sbox_n24) );
  XNOR2_X1 aes_sbox_input_mapping_1_U14 ( .A(aes_sbox_input_mapping_1_n20), 
        .B(aes_sbox_input_mapping_1_n19), .ZN(aes_sbox_mappedxD_1__3_) );
  XNOR2_X1 aes_sbox_input_mapping_1_U13 ( .A(aes_sbox_input_mapping_1_n18), 
        .B(CxDO[11]), .ZN(aes_sbox_input_mapping_1_n19) );
  XNOR2_X1 aes_sbox_input_mapping_1_U12 ( .A(CxDO[15]), .B(CxDO[12]), .ZN(
        aes_sbox_input_mapping_1_n18) );
  XNOR2_X1 aes_sbox_input_mapping_1_U11 ( .A(aes_sbox_input_mapping_1_n17), 
        .B(CxDO[11]), .ZN(aes_sbox_mappedxD_1__0_) );
  XNOR2_X1 aes_sbox_input_mapping_1_U10 ( .A(aes_sbox_input_mapping_1_n23), 
        .B(CxDO[14]), .ZN(aes_sbox_input_mapping_1_n17) );
  XNOR2_X1 aes_sbox_input_mapping_1_U9 ( .A(aes_sbox_input_mapping_1_n23), .B(
        aes_sbox_input_mapping_1_n22), .ZN(aes_sbox_mappedxD_1__7_) );
  XOR2_X1 aes_sbox_input_mapping_1_U8 ( .A(CxDO[12]), .B(
        aes_sbox_mappedxD_1__1_), .Z(aes_sbox_mappedxD_1__6_) );
  XNOR2_X1 aes_sbox_input_mapping_1_U7 ( .A(aes_sbox_input_mapping_1_n21), .B(
        aes_sbox_input_mapping_1_n20), .ZN(aes_sbox_mappedxD_1__5_) );
  XNOR2_X1 aes_sbox_input_mapping_1_U6 ( .A(CxDO[8]), .B(
        aes_sbox_input_mapping_1_n22), .ZN(aes_sbox_mappedxD_1__4_) );
  XOR2_X1 aes_sbox_input_mapping_1_U5 ( .A(CxDO[8]), .B(
        aes_sbox_input_mapping_1_n21), .Z(aes_sbox_mappedxD_1__1_) );
  XNOR2_X1 aes_sbox_input_mapping_1_U4 ( .A(CxDO[10]), .B(
        aes_sbox_input_mapping_1_n20), .ZN(aes_sbox_input_mapping_1_n23) );
  XNOR2_X1 aes_sbox_input_mapping_1_U3 ( .A(CxDO[15]), .B(
        aes_sbox_input_mapping_1_n21), .ZN(aes_sbox_input_mapping_1_n22) );
  XOR2_X1 aes_sbox_input_mapping_1_U2 ( .A(CxDO[14]), .B(CxDO[13]), .Z(
        aes_sbox_input_mapping_1_n21) );
  XNOR2_X1 aes_sbox_input_mapping_1_U1 ( .A(CxDO[8]), .B(CxDO[9]), .ZN(
        aes_sbox_input_mapping_1_n20) );
  XOR2_X1 aes_sbox_square_scaler_gf24_1_U3 ( .A(aes_sbox_Y0xorY1xD[3]), .B(
        aes_sbox_Y0xorY1xD[5]), .Z(aes_sbox_Y0xorY12xD[6]) );
  XOR2_X1 aes_sbox_square_scaler_gf24_1_U2 ( .A(aes_sbox_Y0xorY12xD[4]), .B(
        aes_sbox_Y0xorY1xD[3]), .Z(aes_sbox_Y0xorY12xD[5]) );
  XOR2_X1 aes_sbox_square_scaler_gf24_1_U1 ( .A(aes_sbox_Y0xorY12xD[4]), .B(
        aes_sbox_Y0xorY1xD[4]), .Z(aes_sbox_Y0xorY12xD[7]) );
  XNOR2_X1 aes_sbox_output_mapping_1_U11 ( .A(aes_sbox_output_mapping_1_n8), 
        .B(aes_sbox_InvUnmappedxD[9]), .ZN(StateInxD[9]) );
  XNOR2_X1 aes_sbox_output_mapping_1_U10 ( .A(aes_sbox_InvUnmappedxD[13]), .B(
        aes_sbox_InvUnmappedxD[12]), .ZN(aes_sbox_output_mapping_1_n8) );
  XOR2_X1 aes_sbox_output_mapping_1_U9 ( .A(aes_sbox_InvUnmappedxD[14]), .B(
        aes_sbox_InvUnmappedxD[8]), .Z(StateInxD[13]) );
  XNOR2_X1 aes_sbox_output_mapping_1_U8 ( .A(aes_sbox_output_mapping_1_n7), 
        .B(StateInxD[13]), .ZN(StateInxD[10]) );
  XNOR2_X1 aes_sbox_output_mapping_1_U7 ( .A(StateInxD[15]), .B(
        aes_sbox_InvUnmappedxD[10]), .ZN(aes_sbox_output_mapping_1_n7) );
  XNOR2_X1 aes_sbox_output_mapping_1_U6 ( .A(aes_sbox_InvUnmappedxD[9]), .B(
        aes_sbox_output_mapping_1_n9), .ZN(StateInxD[8]) );
  XNOR2_X1 aes_sbox_output_mapping_1_U5 ( .A(StateInxD[12]), .B(
        aes_sbox_output_mapping_1_n9), .ZN(StateInxD[11]) );
  XOR2_X1 aes_sbox_output_mapping_1_U4 ( .A(StateInxD[15]), .B(
        aes_sbox_InvUnmappedxD[15]), .Z(StateInxD[12]) );
  XOR2_X1 aes_sbox_output_mapping_1_U3 ( .A(aes_sbox_InvUnmappedxD[11]), .B(
        aes_sbox_InvUnmappedxD[15]), .Z(StateInxD[14]) );
  XOR2_X1 aes_sbox_output_mapping_1_U2 ( .A(aes_sbox_InvUnmappedxD[11]), .B(
        aes_sbox_InvUnmappedxD[13]), .Z(StateInxD[15]) );
  XNOR2_X1 aes_sbox_output_mapping_1_U1 ( .A(aes_sbox_InvUnmappedxD[14]), .B(
        aes_sbox_InvUnmappedxD[12]), .ZN(aes_sbox_output_mapping_1_n9) );
  XNOR2_X1 aes_sbox_input_mapping_0_U14 ( .A(aes_sbox_input_mapping_0_n20), 
        .B(aes_sbox_input_mapping_0_n19), .ZN(aes_sbox_mappedxD_0__3_) );
  XNOR2_X1 aes_sbox_input_mapping_0_U13 ( .A(aes_sbox_input_mapping_0_n18), 
        .B(CxDO[3]), .ZN(aes_sbox_input_mapping_0_n19) );
  XNOR2_X1 aes_sbox_input_mapping_0_U12 ( .A(CxDO[7]), .B(CxDO[4]), .ZN(
        aes_sbox_input_mapping_0_n18) );
  XNOR2_X1 aes_sbox_input_mapping_0_U11 ( .A(aes_sbox_input_mapping_0_n17), 
        .B(CxDO[3]), .ZN(aes_sbox_mappedxD_0__0_) );
  XNOR2_X1 aes_sbox_input_mapping_0_U10 ( .A(aes_sbox_input_mapping_0_n23), 
        .B(CxDO[6]), .ZN(aes_sbox_input_mapping_0_n17) );
  XNOR2_X1 aes_sbox_input_mapping_0_U9 ( .A(aes_sbox_input_mapping_0_n23), .B(
        aes_sbox_input_mapping_0_n22), .ZN(aes_sbox_mappedxD_0__7_) );
  XOR2_X1 aes_sbox_input_mapping_0_U8 ( .A(CxDO[4]), .B(
        aes_sbox_mappedxD_0__1_), .Z(aes_sbox_mappedxD_0__6_) );
  XNOR2_X1 aes_sbox_input_mapping_0_U7 ( .A(aes_sbox_input_mapping_0_n21), .B(
        aes_sbox_input_mapping_0_n20), .ZN(aes_sbox_mappedxD_0__5_) );
  XNOR2_X1 aes_sbox_input_mapping_0_U6 ( .A(CxDO[0]), .B(
        aes_sbox_input_mapping_0_n22), .ZN(aes_sbox_mappedxD_0__4_) );
  XOR2_X1 aes_sbox_input_mapping_0_U5 ( .A(CxDO[0]), .B(
        aes_sbox_input_mapping_0_n21), .Z(aes_sbox_mappedxD_0__1_) );
  XNOR2_X1 aes_sbox_input_mapping_0_U4 ( .A(CxDO[2]), .B(
        aes_sbox_input_mapping_0_n20), .ZN(aes_sbox_input_mapping_0_n23) );
  XNOR2_X1 aes_sbox_input_mapping_0_U3 ( .A(CxDO[7]), .B(
        aes_sbox_input_mapping_0_n21), .ZN(aes_sbox_input_mapping_0_n22) );
  XOR2_X1 aes_sbox_input_mapping_0_U2 ( .A(CxDO[6]), .B(CxDO[5]), .Z(
        aes_sbox_input_mapping_0_n21) );
  XNOR2_X1 aes_sbox_input_mapping_0_U1 ( .A(CxDO[0]), .B(CxDO[1]), .ZN(
        aes_sbox_input_mapping_0_n20) );
  XOR2_X1 aes_sbox_square_scaler_gf24_0_U3 ( .A(aes_sbox_Y0xorY12xD[0]), .B(
        aes_sbox_Y0xorY1xD[0]), .Z(aes_sbox_Y0xorY12xD[1]) );
  XOR2_X1 aes_sbox_square_scaler_gf24_0_U2 ( .A(aes_sbox_Y0xorY1xD[0]), .B(
        aes_sbox_Y0xorY1xD[2]), .Z(aes_sbox_Y0xorY12xD[2]) );
  XOR2_X1 aes_sbox_square_scaler_gf24_0_U1 ( .A(aes_sbox_Y0xorY12xD[0]), .B(
        aes_sbox_Y0xorY1xD[1]), .Z(aes_sbox_Y0xorY12xD[3]) );
  XNOR2_X1 aes_sbox_output_mapping_0_U11 ( .A(aes_sbox_InvUnmappedxD[1]), .B(
        aes_sbox_output_mapping_0_n9), .ZN(aes_sbox_InvMappedxD_0__0_) );
  XOR2_X1 aes_sbox_output_mapping_0_U10 ( .A(aes_sbox_InvUnmappedxD[3]), .B(
        aes_sbox_InvUnmappedxD[7]), .Z(aes_sbox_InvMappedxD_0__6_) );
  XNOR2_X1 aes_sbox_output_mapping_0_U9 ( .A(aes_sbox_output_mapping_0_n8), 
        .B(aes_sbox_InvUnmappedxD[1]), .ZN(aes_sbox_InvMappedxD_0__1_) );
  XNOR2_X1 aes_sbox_output_mapping_0_U8 ( .A(aes_sbox_InvUnmappedxD[4]), .B(
        aes_sbox_InvUnmappedxD[5]), .ZN(aes_sbox_output_mapping_0_n8) );
  XNOR2_X1 aes_sbox_output_mapping_0_U7 ( .A(aes_sbox_output_mapping_0_n7), 
        .B(aes_sbox_InvUnmappedxD[2]), .ZN(StateInxD[2]) );
  XNOR2_X1 aes_sbox_output_mapping_0_U6 ( .A(aes_sbox_InvMappedxD_0__5_), .B(
        StateInxD[7]), .ZN(aes_sbox_output_mapping_0_n7) );
  XOR2_X1 aes_sbox_output_mapping_0_U5 ( .A(aes_sbox_InvUnmappedxD[6]), .B(
        aes_sbox_InvUnmappedxD[0]), .Z(aes_sbox_InvMappedxD_0__5_) );
  XNOR2_X1 aes_sbox_output_mapping_0_U4 ( .A(StateInxD[4]), .B(
        aes_sbox_output_mapping_0_n9), .ZN(StateInxD[3]) );
  XOR2_X1 aes_sbox_output_mapping_0_U3 ( .A(StateInxD[7]), .B(
        aes_sbox_InvUnmappedxD[7]), .Z(StateInxD[4]) );
  XOR2_X1 aes_sbox_output_mapping_0_U2 ( .A(aes_sbox_InvUnmappedxD[3]), .B(
        aes_sbox_InvUnmappedxD[5]), .Z(StateInxD[7]) );
  XNOR2_X1 aes_sbox_output_mapping_0_U1 ( .A(aes_sbox_InvUnmappedxD[6]), .B(
        aes_sbox_InvUnmappedxD[4]), .ZN(aes_sbox_output_mapping_0_n9) );
  XOR2_X1 aes_sbox_mul_y0y1_U18 ( .A(aes_sbox_mul_y0y1_n2), .B(
        aes_sbox_mul_y0y1_n1), .Z(aes_sbox_Y0mulY1xD[7]) );
  XOR2_X1 aes_sbox_mul_y0y1_U17 ( .A(aes_sbox_mul_y0y1_n4), .B(
        aes_sbox_mul_y0y1_n3), .Z(aes_sbox_Y0mulY1xD[6]) );
  XOR2_X1 aes_sbox_mul_y0y1_U16 ( .A(aes_sbox_mul_y0y1_n6), .B(
        aes_sbox_mul_y0y1_n5), .Z(aes_sbox_Y0mulY1xD[5]) );
  XOR2_X1 aes_sbox_mul_y0y1_U15 ( .A(aes_sbox_mul_y0y1_n8), .B(
        aes_sbox_mul_y0y1_n7), .Z(aes_sbox_Y0mulY1xD[4]) );
  XOR2_X1 aes_sbox_mul_y0y1_U14 ( .A(aes_sbox_mul_y0y1_n10), .B(
        aes_sbox_mul_y0y1_n9), .Z(aes_sbox_Y0mulY1xD[3]) );
  XOR2_X1 aes_sbox_mul_y0y1_U13 ( .A(aes_sbox_mul_y0y1_n12), .B(
        aes_sbox_mul_y0y1_n11), .Z(aes_sbox_Y0mulY1xD[2]) );
  XOR2_X1 aes_sbox_mul_y0y1_U12 ( .A(aes_sbox_mul_y0y1_n14), .B(
        aes_sbox_mul_y0y1_n13), .Z(aes_sbox_Y0mulY1xD[1]) );
  XOR2_X1 aes_sbox_mul_y0y1_U11 ( .A(aes_sbox_mul_y0y1_n16), .B(
        aes_sbox_mul_y0y1_n15), .Z(aes_sbox_Y0mulY1xD[0]) );
  XOR2_X1 aes_sbox_mul_y0y1_U10 ( .A(Zmul1xDI[0]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__0_), .Z(aes_sbox_mul_y0y1_FFxDN[8]) );
  XOR2_X1 aes_sbox_mul_y0y1_U9 ( .A(Zmul1xDI[3]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__3_), .Z(aes_sbox_mul_y0y1_FFxDN[11]) );
  XOR2_X1 aes_sbox_mul_y0y1_U8 ( .A(Zmul1xDI[3]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__3_), .Z(aes_sbox_mul_y0y1_FFxDN[7]) );
  XOR2_X1 aes_sbox_mul_y0y1_U7 ( .A(Zmul1xDI[2]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__2_), .Z(aes_sbox_mul_y0y1_FFxDN[10]) );
  XOR2_X1 aes_sbox_mul_y0y1_U6 ( .A(Zmul1xDI[1]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__1_), .Z(aes_sbox_mul_y0y1_FFxDN[9]) );
  XOR2_X1 aes_sbox_mul_y0y1_U5 ( .A(Zmul1xDI[2]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__2_), .Z(aes_sbox_mul_y0y1_FFxDN[6]) );
  XOR2_X1 aes_sbox_mul_y0y1_U4 ( .A(Zmul1xDI[1]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__1_), .Z(aes_sbox_mul_y0y1_FFxDN[5]) );
  XOR2_X1 aes_sbox_mul_y0y1_U3 ( .A(Zmul1xDI[0]), .B(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__0_), .Z(aes_sbox_mul_y0y1_FFxDN[4]) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_0__0_ ( .D(aes_sbox_mul_y0y1_FFxDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n15) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_0__1_ ( .D(aes_sbox_mul_y0y1_FFxDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n13) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_0__2_ ( .D(aes_sbox_mul_y0y1_FFxDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n11) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_0__3_ ( .D(aes_sbox_mul_y0y1_FFxDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n9) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_1__0_ ( .D(aes_sbox_mul_y0y1_FFxDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n16) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_1__1_ ( .D(aes_sbox_mul_y0y1_FFxDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n14) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_1__2_ ( .D(aes_sbox_mul_y0y1_FFxDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n12) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_1__3_ ( .D(aes_sbox_mul_y0y1_FFxDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n10) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_2__0_ ( .D(aes_sbox_mul_y0y1_FFxDN[8]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n7) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_2__1_ ( .D(aes_sbox_mul_y0y1_FFxDN[9]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n5) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_2__2_ ( .D(aes_sbox_mul_y0y1_FFxDN[10]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n3) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_2__3_ ( .D(aes_sbox_mul_y0y1_FFxDN[11]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n1) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_3__0_ ( .D(aes_sbox_mul_y0y1_FFxDN[12]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n8) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_3__1_ ( .D(aes_sbox_mul_y0y1_FFxDN[13]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n6) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_3__2_ ( .D(aes_sbox_mul_y0y1_FFxDN[14]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n4) );
  DFFR_X1 aes_sbox_mul_y0y1_FFxDP_reg_3__3_ ( .D(aes_sbox_mul_y0y1_FFxDN[15]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mul_y0y1_n2) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U29 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n67), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n68), .ZN(aes_sbox_mul_y0y1_FFxDN[15])
         );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U28 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n77), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n76), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n68) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U27 ( .A1(aes_sbox_Y0xD_1__3_), .A2(
        aes_sbox_Y1xD_1__3_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n67) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U26 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n65), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n66), .ZN(aes_sbox_mul_y0y1_FFxDN[14])
         );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U25 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n76), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n75), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n66) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U24 ( .A1(aes_sbox_Y1xD_1__2_), .A2(
        aes_sbox_Y0xD_1__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n65) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U23 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n63), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n64), .ZN(aes_sbox_mul_y0y1_FFxDN[13])
         );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U22 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n77), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n74), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n64) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U21 ( .A1(aes_sbox_Y0xD_1__1_), .A2(
        aes_sbox_Y1xD_1__1_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n63) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U20 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n61), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n62), .ZN(aes_sbox_mul_y0y1_FFxDN[12])
         );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U19 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n74), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n75), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n62) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U18 ( .A1(aes_sbox_Y1xD_1__0_), .A2(
        aes_sbox_Y0xD_1__0_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n61) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U17 ( .B1(aes_sbox_Y1xD_1__3_), .B2(
        aes_sbox_Y1xD_1__2_), .C1(aes_sbox_Y0xD_1__3_), .C2(
        aes_sbox_Y0xD_1__2_), .A(aes_sbox_mul_y0y1_gf4_mul_1_1_n60), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n76) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U16 ( .A1(aes_sbox_Y1xD_1__3_), .A2(
        aes_sbox_Y1xD_1__2_), .B1(aes_sbox_Y0xD_1__2_), .B2(
        aes_sbox_Y0xD_1__3_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n60) );
  INV_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U14 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n72), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n58) );
  INV_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U13 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n70), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n57) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U12 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n55), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n71), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n56) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U11 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n72), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n73), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n55) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U10 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n53), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n54), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n75) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U9 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n70), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n72), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n54) );
  NOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U8 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n73), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n71), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n53) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U7 ( .A1(aes_sbox_Y0xD_1__0_), .A2(
        aes_sbox_Y0xD_1__1_), .B1(aes_sbox_Y1xD_1__1_), .B2(
        aes_sbox_Y1xD_1__0_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n69) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U6 ( .B1(aes_sbox_Y0xD_1__0_), .B2(
        aes_sbox_Y0xD_1__1_), .C1(aes_sbox_Y1xD_1__0_), .C2(
        aes_sbox_Y1xD_1__1_), .A(aes_sbox_mul_y0y1_gf4_mul_1_1_n69), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n74) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U5 ( .A(aes_sbox_Y1xD_1__0_), .B(
        aes_sbox_Y1xD_1__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n71) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U4 ( .A(aes_sbox_Y1xD_1__1_), .B(
        aes_sbox_Y1xD_1__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_1_1_n72) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U3 ( .A(aes_sbox_Y0xD_1__0_), .B(
        aes_sbox_Y0xD_1__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_1_n73) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U2 ( .A(aes_sbox_Y0xD_1__1_), .B(
        aes_sbox_Y0xD_1__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_1_1_n70) );
  OAI33_X1 aes_sbox_mul_y0y1_gf4_mul_1_1_U1 ( .A1(1'b0), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n56), .A3(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n57), .B1(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n70), .B2(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n73), .B3(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n58), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_1_n77) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U28 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n63), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n62), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n74) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U27 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n60), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n61), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__0_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U26 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n74), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n72), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n61) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U25 ( .A1(aes_sbox_Y0xD_0__0_), .A2(
        aes_sbox_Y1xD_1__0_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n60) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U24 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n58), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n59), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__3_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U23 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n76), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n75), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n59) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U22 ( .A1(aes_sbox_Y0xD_0__3_), .A2(
        aes_sbox_Y1xD_1__3_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n58) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U21 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n56), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n57), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__2_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U20 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n75), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n74), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n57) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U19 ( .A1(aes_sbox_Y0xD_0__2_), .A2(
        aes_sbox_Y1xD_1__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n56) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U18 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n54), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n55), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_2__1_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U17 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n76), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n72), .Z(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n55) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U16 ( .A1(aes_sbox_Y0xD_0__1_), .A2(
        aes_sbox_Y1xD_1__1_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n54) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U15 ( .B1(aes_sbox_Y1xD_1__1_), .B2(
        aes_sbox_Y1xD_1__0_), .C1(aes_sbox_Y0xD_0__1_), .C2(
        aes_sbox_Y0xD_0__0_), .A(aes_sbox_mul_y0y1_gf4_mul_1_0_n53), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n72) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U14 ( .A1(aes_sbox_Y1xD_1__1_), .A2(
        aes_sbox_Y1xD_1__0_), .B1(aes_sbox_Y0xD_0__0_), .B2(
        aes_sbox_Y0xD_0__1_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n53) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U13 ( .A1(aes_sbox_Y0xD_0__2_), .A2(
        aes_sbox_Y0xD_0__3_), .B1(aes_sbox_Y1xD_1__3_), .B2(
        aes_sbox_Y1xD_1__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n73) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U12 ( .B1(aes_sbox_Y0xD_0__2_), .B2(
        aes_sbox_Y0xD_0__3_), .C1(aes_sbox_Y1xD_1__2_), .C2(
        aes_sbox_Y1xD_1__3_), .A(aes_sbox_mul_y0y1_gf4_mul_1_0_n73), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n75) );
  INV_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U11 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n64), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n71) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U10 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n67), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n69), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n65) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U9 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n67), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n71), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n68) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U8 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n66), .B(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n65), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n70) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U7 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n71), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n70), .B1(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n69), .B2(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n68), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n76) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U6 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n67), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n64), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n62) );
  NOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U5 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n69), .A2(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n66), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_1_0_n63) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U4 ( .A(aes_sbox_Y1xD_1__0_), .B(
        aes_sbox_Y1xD_1__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n66) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U3 ( .A(aes_sbox_Y1xD_1__1_), .B(
        aes_sbox_Y1xD_1__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_1_0_n67) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U2 ( .A(aes_sbox_Y0xD_0__0_), .B(
        aes_sbox_Y0xD_0__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_1_0_n69) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_1_0_U1 ( .A(aes_sbox_Y0xD_0__1_), .B(
        aes_sbox_Y0xD_0__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_1_0_n64) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U28 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n63), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n62), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n74) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U27 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n59), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n60), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__3_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U26 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n76), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n75), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n60) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U25 ( .A1(aes_sbox_Y0xD_1__3_), .A2(
        aes_sbox_Y1xD_0__3_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n59) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U24 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n57), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n58), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__2_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U23 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n74), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n75), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n58) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U22 ( .A1(aes_sbox_Y0xD_1__2_), .A2(
        aes_sbox_Y1xD_0__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n57) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U21 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n55), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n56), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__1_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U20 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n76), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n72), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n56) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U19 ( .A1(aes_sbox_Y0xD_1__1_), .A2(
        aes_sbox_Y1xD_0__1_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n55) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U18 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n53), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n54), .ZN(
        aes_sbox_mul_y0y1_Xi_mul_Yj_1__0_) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U17 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n72), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n74), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n54) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U16 ( .A1(aes_sbox_Y0xD_1__0_), .A2(
        aes_sbox_Y1xD_0__0_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n53) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U15 ( .A1(aes_sbox_Y0xD_1__2_), .A2(
        aes_sbox_Y0xD_1__3_), .B1(aes_sbox_Y1xD_0__3_), .B2(
        aes_sbox_Y1xD_0__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n73) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U14 ( .B1(aes_sbox_Y0xD_1__2_), .B2(
        aes_sbox_Y0xD_1__3_), .C1(aes_sbox_Y1xD_0__2_), .C2(
        aes_sbox_Y1xD_0__3_), .A(aes_sbox_mul_y0y1_gf4_mul_0_1_n73), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n75) );
  INV_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U13 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n64), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n71) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U12 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n67), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n69), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n65) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U11 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n67), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n71), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n68) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U10 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n66), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n65), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n70) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U9 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n71), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n70), .B1(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n69), .B2(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n68), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n76) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U8 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n67), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n64), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n62) );
  NOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U7 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n69), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n66), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n63) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U6 ( .A1(aes_sbox_Y0xD_1__0_), .A2(
        aes_sbox_Y0xD_1__1_), .B1(aes_sbox_Y1xD_0__1_), .B2(
        aes_sbox_Y1xD_0__0_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n61) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U5 ( .B1(aes_sbox_Y0xD_1__0_), .B2(
        aes_sbox_Y0xD_1__1_), .C1(aes_sbox_Y1xD_0__0_), .C2(
        aes_sbox_Y1xD_0__1_), .A(aes_sbox_mul_y0y1_gf4_mul_0_1_n61), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_1_n72) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U4 ( .A(aes_sbox_Y1xD_0__0_), .B(
        aes_sbox_Y1xD_0__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n66) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U3 ( .A(aes_sbox_Y1xD_0__1_), .B(
        aes_sbox_Y1xD_0__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_0_1_n67) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U2 ( .A(aes_sbox_Y0xD_1__0_), .B(
        aes_sbox_Y0xD_1__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_1_n69) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_1_U1 ( .A(aes_sbox_Y0xD_1__1_), .B(
        aes_sbox_Y0xD_1__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_0_1_n64) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U29 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n69), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n68), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n75) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U28 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n66), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n67), .ZN(aes_sbox_mul_y0y1_FFxDN[3]) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U27 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n77), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n76), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n67) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U26 ( .A1(aes_sbox_Y0xD_0__3_), .A2(
        aes_sbox_Y1xD_0__3_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n66) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U25 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n64), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n65), .ZN(aes_sbox_mul_y0y1_FFxDN[0]) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U24 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n74), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n75), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n65) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U23 ( .A1(aes_sbox_Y1xD_0__0_), .A2(
        aes_sbox_Y0xD_0__0_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n64) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U22 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n62), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n63), .ZN(aes_sbox_mul_y0y1_FFxDN[1]) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U21 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n77), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n74), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n63) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U20 ( .A1(aes_sbox_Y0xD_0__1_), .A2(
        aes_sbox_Y1xD_0__1_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n62) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U19 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n60), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n61), .ZN(aes_sbox_mul_y0y1_FFxDN[2]) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U18 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n76), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n75), .Z(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n61) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U17 ( .A1(aes_sbox_Y1xD_0__2_), .A2(
        aes_sbox_Y0xD_0__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n60) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U16 ( .B1(aes_sbox_Y1xD_0__3_), .B2(
        aes_sbox_Y1xD_0__2_), .C1(aes_sbox_Y0xD_0__3_), .C2(
        aes_sbox_Y0xD_0__2_), .A(aes_sbox_mul_y0y1_gf4_mul_0_0_n59), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n76) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U15 ( .A1(aes_sbox_Y1xD_0__3_), .A2(
        aes_sbox_Y1xD_0__2_), .B1(aes_sbox_Y0xD_0__2_), .B2(
        aes_sbox_Y0xD_0__3_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n59) );
  AOI221_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U14 ( .B1(aes_sbox_Y1xD_0__1_), .B2(
        aes_sbox_Y1xD_0__0_), .C1(aes_sbox_Y0xD_0__1_), .C2(
        aes_sbox_Y0xD_0__0_), .A(aes_sbox_mul_y0y1_gf4_mul_0_0_n58), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n74) );
  OAI22_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U13 ( .A1(aes_sbox_Y1xD_0__1_), .A2(
        aes_sbox_Y1xD_0__0_), .B1(aes_sbox_Y0xD_0__0_), .B2(
        aes_sbox_Y0xD_0__1_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n58) );
  INV_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U12 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n72), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n57) );
  INV_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U11 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n70), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n56) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U10 ( .A(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n54), .B(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n71), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n55) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U9 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n72), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n73), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n54) );
  NAND2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U7 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n72), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n70), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n68) );
  NOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U6 ( .A1(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n73), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n71), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n69) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U5 ( .A(aes_sbox_Y1xD_0__0_), .B(
        aes_sbox_Y1xD_0__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n71) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U4 ( .A(aes_sbox_Y1xD_0__1_), .B(
        aes_sbox_Y1xD_0__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_0_0_n72) );
  XNOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U3 ( .A(aes_sbox_Y0xD_0__0_), .B(
        aes_sbox_Y0xD_0__2_), .ZN(aes_sbox_mul_y0y1_gf4_mul_0_0_n73) );
  XOR2_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U2 ( .A(aes_sbox_Y0xD_0__1_), .B(
        aes_sbox_Y0xD_0__3_), .Z(aes_sbox_mul_y0y1_gf4_mul_0_0_n70) );
  OAI33_X1 aes_sbox_mul_y0y1_gf4_mul_0_0_U1 ( .A1(1'b0), .A2(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n55), .A3(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n56), .B1(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n70), .B2(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n73), .B3(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n57), .ZN(
        aes_sbox_mul_y0y1_gf4_mul_0_0_n77) );
  XNOR2_X1 aes_sbox_inverter_gf24_U12 ( .A(aes_sbox_inverter_gf24_AmulBxD[2]), 
        .B(aes_sbox_inverter_gf24_n3), .ZN(aes_sbox_inverter_gf24_ExD[3]) );
  XNOR2_X1 aes_sbox_inverter_gf24_U11 ( .A(aes_sbox_inverter_gf24_AmulBxD[3]), 
        .B(aes_sbox_inverter_gf24_n4), .ZN(aes_sbox_inverter_gf24_ExD[2]) );
  XNOR2_X1 aes_sbox_inverter_gf24_U10 ( .A(aes_sbox_inverter_gf24_AmulBxD[0]), 
        .B(aes_sbox_inverter_gf24_n5), .ZN(aes_sbox_inverter_gf24_ExD[1]) );
  XNOR2_X1 aes_sbox_inverter_gf24_U9 ( .A(aes_sbox_inverter_gf24_AmulBxD[1]), 
        .B(aes_sbox_inverter_gf24_n6), .ZN(aes_sbox_inverter_gf24_ExD[0]) );
  XNOR2_X1 aes_sbox_inverter_gf24_U8 ( .A(aes_sbox_inverter_gf24_n2), .B(
        aes_sbox_InverterInxDP[6]), .ZN(aes_sbox_inverter_gf24_n7) );
  XNOR2_X1 aes_sbox_inverter_gf24_U7 ( .A(aes_sbox_inverter_gf24_d_1__0_), .B(
        aes_sbox_InverterInxDP[4]), .ZN(aes_sbox_inverter_gf24_n2) );
  XNOR2_X1 aes_sbox_inverter_gf24_U6 ( .A(aes_sbox_inverter_gf24_n1), .B(
        aes_sbox_InverterInxDP[2]), .ZN(aes_sbox_inverter_gf24_n8) );
  XNOR2_X1 aes_sbox_inverter_gf24_U5 ( .A(aes_sbox_inverter_gf24_d_0__0_), .B(
        aes_sbox_InverterInxDP[0]), .ZN(aes_sbox_inverter_gf24_n1) );
  XOR2_X1 aes_sbox_inverter_gf24_U4 ( .A(aes_sbox_InverterInxDP[5]), .B(
        aes_sbox_InverterInxDP[7]), .Z(aes_sbox_inverter_gf24_d_1__0_) );
  XOR2_X1 aes_sbox_inverter_gf24_U3 ( .A(aes_sbox_InverterInxDP[1]), .B(
        aes_sbox_InverterInxDP[3]), .Z(aes_sbox_inverter_gf24_d_0__0_) );
  DFFR_X1 aes_sbox_inverter_gf24_ExDP_reg_0__0_ ( .D(
        aes_sbox_inverter_gf24_ExD[0]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_ExDP_0__0_), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_ExDP_reg_0__1_ ( .D(
        aes_sbox_inverter_gf24_ExD[1]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_ExDP_0__1_), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_ExDP_reg_1__0_ ( .D(
        aes_sbox_inverter_gf24_ExD[2]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_ExDP_1__0_), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_ExDP_reg_1__1_ ( .D(
        aes_sbox_inverter_gf24_ExD[3]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_ExDP_1__1_), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_CxDP_reg_0__0_ ( .D(aes_sbox_inverter_gf24_n8), .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_inverter_gf24_n5) );
  DFFR_X1 aes_sbox_inverter_gf24_CxDP_reg_0__1_ ( .D(
        aes_sbox_inverter_gf24_d_0__0_), .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(
        aes_sbox_inverter_gf24_n6) );
  DFFR_X1 aes_sbox_inverter_gf24_CxDP_reg_1__0_ ( .D(aes_sbox_inverter_gf24_n7), .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_inverter_gf24_n3) );
  DFFR_X1 aes_sbox_inverter_gf24_CxDP_reg_1__1_ ( .D(
        aes_sbox_inverter_gf24_d_1__0_), .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(
        aes_sbox_inverter_gf24_n4) );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedBxDP_reg_0__0_ ( .D(
        aes_sbox_inverter_gf24_BxDP[0]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedBxDP[0]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_BxDP_reg_0__0_ ( .D(aes_sbox_InverterInxDP[0]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_BxDP[0]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedBxDP_reg_0__1_ ( .D(
        aes_sbox_inverter_gf24_BxDP[1]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedBxDP[1]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_BxDP_reg_0__1_ ( .D(aes_sbox_InverterInxDP[1]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_BxDP[1]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedBxDP_reg_1__0_ ( .D(
        aes_sbox_inverter_gf24_BxDP[2]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedBxDP[2]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_BxDP_reg_1__0_ ( .D(aes_sbox_InverterInxDP[4]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_BxDP[2]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedBxDP_reg_1__1_ ( .D(
        aes_sbox_inverter_gf24_BxDP[3]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedBxDP[3]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_BxDP_reg_1__1_ ( .D(aes_sbox_InverterInxDP[5]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_BxDP[3]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedAxDP_reg_0__0_ ( .D(
        aes_sbox_inverter_gf24_AxDP[0]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedAxDP[0]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_AxDP_reg_0__0_ ( .D(aes_sbox_InverterInxDP[2]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_AxDP[0]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedAxDP_reg_0__1_ ( .D(
        aes_sbox_inverter_gf24_AxDP[1]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedAxDP[1]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_AxDP_reg_0__1_ ( .D(aes_sbox_InverterInxDP[3]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_AxDP[1]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedAxDP_reg_1__0_ ( .D(
        aes_sbox_inverter_gf24_AxDP[2]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedAxDP[2]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_AxDP_reg_1__0_ ( .D(aes_sbox_InverterInxDP[6]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_AxDP[2]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_pipelinedAxDP_reg_1__1_ ( .D(
        aes_sbox_inverter_gf24_AxDP[3]), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_sbox_inverter_gf24_pipelinedAxDP[3]), .QN() );
  DFFR_X1 aes_sbox_inverter_gf24_AxDP_reg_1__1_ ( .D(aes_sbox_InverterInxDP[7]), .CK(ClkxCI), .RN(RstxBI), .Q(aes_sbox_inverter_gf24_AxDP[3]), .QN() );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U10 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_n2), .B(
        aes_sbox_inverter_gf24_a_mul_b_n1), .Z(
        aes_sbox_inverter_gf24_AmulBxD[3]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U9 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_n4), .B(
        aes_sbox_inverter_gf24_a_mul_b_n3), .Z(
        aes_sbox_inverter_gf24_AmulBxD[2]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U8 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_n6), .B(
        aes_sbox_inverter_gf24_a_mul_b_n5), .Z(
        aes_sbox_inverter_gf24_AmulBxD[1]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U7 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_n8), .B(
        aes_sbox_inverter_gf24_a_mul_b_n7), .Z(
        aes_sbox_inverter_gf24_AmulBxD[0]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U6 ( .A(Zinv1xDI[1]), .B(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_), .Z(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[5]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U5 ( .A(Zinv1xDI[1]), .B(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_), .Z(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[3]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U4 ( .A(Zinv1xDI[0]), .B(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_), .Z(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[4]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_b_U3 ( .A(Zinv1xDI[0]), .B(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_), .Z(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[2]) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_0__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[0]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n7) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_0__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[1]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n5) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_1__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[2]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n8) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_1__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[3]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n6) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_2__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[4]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n3) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_2__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[5]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n1) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_3__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[6]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n4) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_b_FFxDP_reg_3__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[7]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_b_n2) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n13), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[7]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_U5 ( .A1(
        aes_sbox_InverterInxDP[7]), .A2(aes_sbox_InverterInxDP[5]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n12), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[6]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_U3 ( .A1(
        aes_sbox_InverterInxDP[6]), .A2(aes_sbox_InverterInxDP[4]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_U2 ( .B1(
        aes_sbox_InverterInxDP[6]), .B2(aes_sbox_InverterInxDP[7]), .C1(
        aes_sbox_InverterInxDP[5]), .C2(aes_sbox_InverterInxDP[4]), .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_U1 ( .A1(
        aes_sbox_InverterInxDP[6]), .A2(aes_sbox_InverterInxDP[7]), .B1(
        aes_sbox_InverterInxDP[4]), .B2(aes_sbox_InverterInxDP[5]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_1_n11) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n13), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_U5 ( .A1(
        aes_sbox_InverterInxDP[7]), .A2(aes_sbox_InverterInxDP[1]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n12), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_U3 ( .A1(
        aes_sbox_InverterInxDP[6]), .A2(aes_sbox_InverterInxDP[0]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_U2 ( .B1(
        aes_sbox_InverterInxDP[6]), .B2(aes_sbox_InverterInxDP[7]), .C1(
        aes_sbox_InverterInxDP[1]), .C2(aes_sbox_InverterInxDP[0]), .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_U1 ( .A1(
        aes_sbox_InverterInxDP[6]), .A2(aes_sbox_InverterInxDP[7]), .B1(
        aes_sbox_InverterInxDP[0]), .B2(aes_sbox_InverterInxDP[1]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_1_0_n11) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n13), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_U5 ( .A1(
        aes_sbox_InverterInxDP[3]), .A2(aes_sbox_InverterInxDP[5]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n12), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_U3 ( .A1(
        aes_sbox_InverterInxDP[2]), .A2(aes_sbox_InverterInxDP[4]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_U2 ( .B1(
        aes_sbox_InverterInxDP[2]), .B2(aes_sbox_InverterInxDP[3]), .C1(
        aes_sbox_InverterInxDP[5]), .C2(aes_sbox_InverterInxDP[4]), .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_U1 ( .A1(
        aes_sbox_InverterInxDP[2]), .A2(aes_sbox_InverterInxDP[3]), .B1(
        aes_sbox_InverterInxDP[4]), .B2(aes_sbox_InverterInxDP[5]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_1_n11) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n13), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[1]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_U5 ( .A1(
        aes_sbox_InverterInxDP[3]), .A2(aes_sbox_InverterInxDP[1]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n12), .B(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_FFxDN[0]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_U3 ( .A1(
        aes_sbox_InverterInxDP[2]), .A2(aes_sbox_InverterInxDP[0]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_U2 ( .B1(
        aes_sbox_InverterInxDP[2]), .B2(aes_sbox_InverterInxDP[3]), .C1(
        aes_sbox_InverterInxDP[1]), .C2(aes_sbox_InverterInxDP[0]), .A(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_U1 ( .A1(
        aes_sbox_InverterInxDP[2]), .A2(aes_sbox_InverterInxDP[3]), .B1(
        aes_sbox_InverterInxDP[0]), .B2(aes_sbox_InverterInxDP[1]), .ZN(
        aes_sbox_inverter_gf24_a_mul_b_gf2_mul_0_0_n11) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_e_U10 ( .A(Zinv2xDI[1]), .B(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_), .Z(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[5]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_e_U9 ( .A(Zinv2xDI[0]), .B(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_), .Z(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[2]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_e_U8 ( .A(Zinv2xDI[0]), .B(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_), .Z(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[4]) );
  XOR2_X1 aes_sbox_inverter_gf24_a_mul_e_U7 ( .A(Zinv2xDI[1]), .B(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_), .Z(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[3]) );
  XOR2_X2 aes_sbox_inverter_gf24_a_mul_e_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_n9), .B(
        aes_sbox_inverter_gf24_a_mul_e_n10), .Z(aes_sbox_InverterOutxD_0__0_)
         );
  XOR2_X2 aes_sbox_inverter_gf24_a_mul_e_U5 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_n11), .B(
        aes_sbox_inverter_gf24_a_mul_e_n12), .Z(aes_sbox_InverterOutxD_0__1_)
         );
  XOR2_X2 aes_sbox_inverter_gf24_a_mul_e_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_n13), .B(
        aes_sbox_inverter_gf24_a_mul_e_n14), .Z(aes_sbox_InverterOutxD_1__0_)
         );
  XOR2_X2 aes_sbox_inverter_gf24_a_mul_e_U3 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_n15), .B(
        aes_sbox_inverter_gf24_a_mul_e_n16), .Z(aes_sbox_InverterOutxD_1__1_)
         );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_0__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[0]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n10) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_0__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[1]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n12) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_1__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[2]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n9) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_1__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[3]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n11) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_2__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[4]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n14) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_2__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[5]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n16) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_3__0_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[6]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n13) );
  DFFR_X1 aes_sbox_inverter_gf24_a_mul_e_FFxDP_reg_3__1_ ( .D(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[7]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_a_mul_e_n15) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n13), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[7]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_U5 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[3]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n12), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[6]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_U3 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[2]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__0_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_U2 ( .B1(
        aes_sbox_inverter_gf24_pipelinedAxDP[2]), .B2(
        aes_sbox_inverter_gf24_pipelinedAxDP[3]), .C1(
        aes_sbox_inverter_gf24_ExDP_1__1_), .C2(
        aes_sbox_inverter_gf24_ExDP_1__0_), .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_U1 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[2]), .A2(
        aes_sbox_inverter_gf24_pipelinedAxDP[3]), .B1(
        aes_sbox_inverter_gf24_ExDP_1__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_1_n11) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n13), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_U5 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[3]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n12), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_U3 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[2]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__0_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_U2 ( .B1(
        aes_sbox_inverter_gf24_pipelinedAxDP[2]), .B2(
        aes_sbox_inverter_gf24_pipelinedAxDP[3]), .C1(
        aes_sbox_inverter_gf24_ExDP_0__1_), .C2(
        aes_sbox_inverter_gf24_ExDP_0__0_), .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_U1 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[2]), .A2(
        aes_sbox_inverter_gf24_pipelinedAxDP[3]), .B1(
        aes_sbox_inverter_gf24_ExDP_0__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_1_0_n11) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n13), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_U5 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[0]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__0_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n12), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_U3 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[1]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_U2 ( .B1(
        aes_sbox_inverter_gf24_pipelinedAxDP[0]), .B2(
        aes_sbox_inverter_gf24_pipelinedAxDP[1]), .C1(
        aes_sbox_inverter_gf24_ExDP_1__1_), .C2(
        aes_sbox_inverter_gf24_ExDP_1__0_), .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_U1 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[0]), .A2(
        aes_sbox_inverter_gf24_pipelinedAxDP[1]), .B1(
        aes_sbox_inverter_gf24_ExDP_1__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_1_n11) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_U6 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n13), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[0]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_U5 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[0]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__0_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_U4 ( .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n12), .B(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n14), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_FFxDN[1]) );
  NAND2_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_U3 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[1]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_U2 ( .B1(
        aes_sbox_inverter_gf24_pipelinedAxDP[0]), .B2(
        aes_sbox_inverter_gf24_pipelinedAxDP[1]), .C1(
        aes_sbox_inverter_gf24_ExDP_0__1_), .C2(
        aes_sbox_inverter_gf24_ExDP_0__0_), .A(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n11), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_U1 ( .A1(
        aes_sbox_inverter_gf24_pipelinedAxDP[0]), .A2(
        aes_sbox_inverter_gf24_pipelinedAxDP[1]), .B1(
        aes_sbox_inverter_gf24_ExDP_0__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .ZN(
        aes_sbox_inverter_gf24_a_mul_e_gf2_mul_0_0_n11) );
  XOR2_X1 aes_sbox_inverter_gf24_b_mul_e_U10 ( .A(Zinv3xDI[0]), .B(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_), .Z(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[4]) );
  XOR2_X1 aes_sbox_inverter_gf24_b_mul_e_U9 ( .A(Zinv3xDI[1]), .B(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_), .Z(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[5]) );
  XOR2_X1 aes_sbox_inverter_gf24_b_mul_e_U8 ( .A(Zinv3xDI[1]), .B(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_), .Z(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[3]) );
  XOR2_X1 aes_sbox_inverter_gf24_b_mul_e_U7 ( .A(Zinv3xDI[0]), .B(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_), .Z(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[2]) );
  XOR2_X2 aes_sbox_inverter_gf24_b_mul_e_U6 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_n13), .B(
        aes_sbox_inverter_gf24_b_mul_e_n14), .Z(aes_sbox_InverterOutxD_1__2_)
         );
  XOR2_X2 aes_sbox_inverter_gf24_b_mul_e_U5 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_n9), .B(
        aes_sbox_inverter_gf24_b_mul_e_n10), .Z(aes_sbox_InverterOutxD_0__2_)
         );
  XOR2_X2 aes_sbox_inverter_gf24_b_mul_e_U4 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_n15), .B(
        aes_sbox_inverter_gf24_b_mul_e_n16), .Z(aes_sbox_InverterOutxD_1__3_)
         );
  XOR2_X2 aes_sbox_inverter_gf24_b_mul_e_U3 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_n11), .B(
        aes_sbox_inverter_gf24_b_mul_e_n12), .Z(aes_sbox_InverterOutxD_0__3_)
         );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_0__0_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[0]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n10) );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_0__1_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[1]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n12) );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_1__0_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[2]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n9) );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_1__1_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[3]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n11) );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_2__0_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[4]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n14) );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_2__1_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[5]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n16) );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_3__0_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[6]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n13) );
  DFFR_X1 aes_sbox_inverter_gf24_b_mul_e_FFxDP_reg_3__1_ ( .D(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[7]), .CK(ClkxCI), .RN(RstxBI), 
        .Q(), .QN(aes_sbox_inverter_gf24_b_mul_e_n15) );
  AOI221_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_U6 ( .B1(
        aes_sbox_inverter_gf24_ExDP_1__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .C1(
        aes_sbox_inverter_gf24_pipelinedBxDP[3]), .C2(
        aes_sbox_inverter_gf24_pipelinedBxDP[2]), .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n13), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_U5 ( .A1(
        aes_sbox_inverter_gf24_ExDP_1__0_), .A2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .B1(
        aes_sbox_inverter_gf24_pipelinedBxDP[2]), .B2(
        aes_sbox_inverter_gf24_pipelinedBxDP[3]), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_U4 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n12), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n14), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[7]) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_U3 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[3]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n12) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_U2 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n11), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n14), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[6]) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_U1 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[2]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__0_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_1_n11) );
  AOI221_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_U6 ( .B1(
        aes_sbox_inverter_gf24_ExDP_0__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .C1(
        aes_sbox_inverter_gf24_pipelinedBxDP[3]), .C2(
        aes_sbox_inverter_gf24_pipelinedBxDP[2]), .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n13), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n14) );
  OAI22_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_U5 ( .A1(
        aes_sbox_inverter_gf24_ExDP_0__0_), .A2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .B1(
        aes_sbox_inverter_gf24_pipelinedBxDP[2]), .B2(
        aes_sbox_inverter_gf24_pipelinedBxDP[3]), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_U4 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n12), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n14), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_U3 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[2]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__0_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n12) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_U2 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n11), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n14), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_U1 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[3]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_1_0_n11) );
  AOI221_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_U6 ( .B1(
        aes_sbox_inverter_gf24_ExDP_1__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .C1(
        aes_sbox_inverter_gf24_pipelinedBxDP[1]), .C2(
        aes_sbox_inverter_gf24_pipelinedBxDP[0]), .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n13), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n14) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_U5 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n12), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n14), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_U4 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[1]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n12) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_U3 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n11), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n14), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_U2 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[0]), .A2(
        aes_sbox_inverter_gf24_ExDP_1__0_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n11) );
  OAI22_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_U1 ( .A1(
        aes_sbox_inverter_gf24_ExDP_1__0_), .A2(
        aes_sbox_inverter_gf24_ExDP_1__1_), .B1(
        aes_sbox_inverter_gf24_pipelinedBxDP[0]), .B2(
        aes_sbox_inverter_gf24_pipelinedBxDP[1]), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_1_n13) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_U6 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n14), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n13), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[1]) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_U5 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[1]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n14) );
  XNOR2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_U4 ( .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n12), .B(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n13), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_FFxDN[0]) );
  NAND2_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_U3 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[0]), .A2(
        aes_sbox_inverter_gf24_ExDP_0__0_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n12) );
  AOI221_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_U2 ( .B1(
        aes_sbox_inverter_gf24_pipelinedBxDP[0]), .B2(
        aes_sbox_inverter_gf24_pipelinedBxDP[1]), .C1(
        aes_sbox_inverter_gf24_ExDP_0__1_), .C2(
        aes_sbox_inverter_gf24_ExDP_0__0_), .A(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n11), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n13) );
  OAI22_X1 aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_U1 ( .A1(
        aes_sbox_inverter_gf24_pipelinedBxDP[0]), .A2(
        aes_sbox_inverter_gf24_pipelinedBxDP[1]), .B1(
        aes_sbox_inverter_gf24_ExDP_0__0_), .B2(
        aes_sbox_inverter_gf24_ExDP_0__1_), .ZN(
        aes_sbox_inverter_gf24_b_mul_e_gf2_mul_0_0_n11) );
  XOR2_X1 aes_sbox_mult_msb_U18 ( .A(aes_sbox_mult_msb_n2), .B(
        aes_sbox_mult_msb_n1), .Z(aes_sbox_InvUnmappedxD[15]) );
  XOR2_X1 aes_sbox_mult_msb_U17 ( .A(aes_sbox_mult_msb_n4), .B(
        aes_sbox_mult_msb_n3), .Z(aes_sbox_InvUnmappedxD[14]) );
  XOR2_X1 aes_sbox_mult_msb_U16 ( .A(aes_sbox_mult_msb_n6), .B(
        aes_sbox_mult_msb_n5), .Z(aes_sbox_InvUnmappedxD[13]) );
  XOR2_X1 aes_sbox_mult_msb_U15 ( .A(aes_sbox_mult_msb_n8), .B(
        aes_sbox_mult_msb_n7), .Z(aes_sbox_InvUnmappedxD[12]) );
  XOR2_X1 aes_sbox_mult_msb_U14 ( .A(aes_sbox_mult_msb_n10), .B(
        aes_sbox_mult_msb_n9), .Z(aes_sbox_InvUnmappedxD[7]) );
  XOR2_X1 aes_sbox_mult_msb_U13 ( .A(aes_sbox_mult_msb_n12), .B(
        aes_sbox_mult_msb_n11), .Z(aes_sbox_InvUnmappedxD[6]) );
  XOR2_X1 aes_sbox_mult_msb_U12 ( .A(aes_sbox_mult_msb_n14), .B(
        aes_sbox_mult_msb_n13), .Z(aes_sbox_InvUnmappedxD[5]) );
  XOR2_X1 aes_sbox_mult_msb_U11 ( .A(aes_sbox_mult_msb_n16), .B(
        aes_sbox_mult_msb_n15), .Z(aes_sbox_InvUnmappedxD[4]) );
  XOR2_X1 aes_sbox_mult_msb_U10 ( .A(Zmul2xDI[1]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_1__1_), .Z(aes_sbox_mult_msb_FFxDN[5]) );
  XOR2_X1 aes_sbox_mult_msb_U9 ( .A(Zmul2xDI[3]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_2__3_), .Z(aes_sbox_mult_msb_FFxDN[11]) );
  XOR2_X1 aes_sbox_mult_msb_U8 ( .A(Zmul2xDI[3]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_1__3_), .Z(aes_sbox_mult_msb_FFxDN[7]) );
  XOR2_X1 aes_sbox_mult_msb_U7 ( .A(Zmul2xDI[2]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_2__2_), .Z(aes_sbox_mult_msb_FFxDN[10]) );
  XOR2_X1 aes_sbox_mult_msb_U6 ( .A(Zmul2xDI[1]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_2__1_), .Z(aes_sbox_mult_msb_FFxDN[9]) );
  XOR2_X1 aes_sbox_mult_msb_U5 ( .A(Zmul2xDI[2]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_1__2_), .Z(aes_sbox_mult_msb_FFxDN[6]) );
  XOR2_X1 aes_sbox_mult_msb_U4 ( .A(Zmul2xDI[0]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_2__0_), .Z(aes_sbox_mult_msb_FFxDN[8]) );
  XOR2_X1 aes_sbox_mult_msb_U3 ( .A(Zmul2xDI[0]), .B(
        aes_sbox_mult_msb_Xi_mul_Yj_1__0_), .Z(aes_sbox_mult_msb_FFxDN[4]) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_0__0_ ( .D(aes_sbox_mult_msb_FFxDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n15) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_0__1_ ( .D(aes_sbox_mult_msb_FFxDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n13) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_0__2_ ( .D(aes_sbox_mult_msb_FFxDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n11) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_0__3_ ( .D(aes_sbox_mult_msb_FFxDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n9) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_1__0_ ( .D(aes_sbox_mult_msb_FFxDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n16) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_1__1_ ( .D(aes_sbox_mult_msb_FFxDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n14) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_1__2_ ( .D(aes_sbox_mult_msb_FFxDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n12) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_1__3_ ( .D(aes_sbox_mult_msb_FFxDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n10) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_2__0_ ( .D(aes_sbox_mult_msb_FFxDN[8]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n7) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_2__1_ ( .D(aes_sbox_mult_msb_FFxDN[9]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n5) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_2__2_ ( .D(aes_sbox_mult_msb_FFxDN[10]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n3) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_2__3_ ( .D(aes_sbox_mult_msb_FFxDN[11]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n1) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_3__0_ ( .D(aes_sbox_mult_msb_FFxDN[12]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n8) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_3__1_ ( .D(aes_sbox_mult_msb_FFxDN[13]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n6) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_3__2_ ( .D(aes_sbox_mult_msb_FFxDN[14]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n4) );
  DFFR_X1 aes_sbox_mult_msb_FFxDP_reg_3__3_ ( .D(aes_sbox_mult_msb_FFxDN[15]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_msb_n2) );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_1_1_U29 ( .B1(aes_sbox_Y0_4xDP[6]), .B2(
        aes_sbox_Y0_4xDP[7]), .C1(aes_sbox_InverterOutxD_1__2_), .C2(
        aes_sbox_InverterOutxD_1__3_), .A(aes_sbox_mult_msb_gf4_mul_1_1_n74), 
        .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n76) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_1_1_U28 ( .A1(aes_sbox_Y0_4xDP[6]), .A2(
        aes_sbox_Y0_4xDP[7]), .B1(aes_sbox_InverterOutxD_1__3_), .B2(
        aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n74)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U27 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n68), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n67), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n75) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U26 ( .A(aes_sbox_InverterOutxD_1__1_), 
        .B(aes_sbox_InverterOutxD_1__3_), .Z(aes_sbox_mult_msb_gf4_mul_1_1_n71) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U25 ( .A(aes_sbox_InverterOutxD_1__0_), .B(aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n70) );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_1_1_U24 ( .B1(aes_sbox_Y0_4xDP[4]), .B2(
        aes_sbox_Y0_4xDP[5]), .C1(aes_sbox_InverterOutxD_1__0_), .C2(
        aes_sbox_InverterOutxD_1__1_), .A(aes_sbox_mult_msb_gf4_mul_1_1_n66), 
        .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n73) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_1_1_U23 ( .A1(aes_sbox_Y0_4xDP[4]), .A2(
        aes_sbox_Y0_4xDP[5]), .B1(aes_sbox_InverterOutxD_1__1_), .B2(
        aes_sbox_InverterOutxD_1__0_), .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n66)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U22 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n64), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n65), .ZN(aes_sbox_mult_msb_FFxDN[15])
         );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U21 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n77), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n76), .Z(
        aes_sbox_mult_msb_gf4_mul_1_1_n65) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U20 ( .A1(aes_sbox_Y0_4xDP[7]), .A2(
        aes_sbox_InverterOutxD_1__3_), .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n64)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U19 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n62), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n63), .ZN(aes_sbox_mult_msb_FFxDN[14])
         );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U18 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n76), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n75), .Z(
        aes_sbox_mult_msb_gf4_mul_1_1_n63) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U17 ( .A1(
        aes_sbox_InverterOutxD_1__2_), .A2(aes_sbox_Y0_4xDP[6]), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n62) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U16 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n60), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n61), .ZN(aes_sbox_mult_msb_FFxDN[13])
         );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U15 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n77), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n73), .Z(
        aes_sbox_mult_msb_gf4_mul_1_1_n61) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U14 ( .A1(aes_sbox_Y0_4xDP[5]), .A2(
        aes_sbox_InverterOutxD_1__1_), .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n60)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U13 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n58), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n59), .ZN(aes_sbox_mult_msb_FFxDN[12])
         );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U12 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n73), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n75), .Z(
        aes_sbox_mult_msb_gf4_mul_1_1_n59) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U11 ( .A1(
        aes_sbox_InverterOutxD_1__0_), .A2(aes_sbox_Y0_4xDP[4]), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n58) );
  INV_X1 aes_sbox_mult_msb_gf4_mul_1_1_U10 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n71), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n57) );
  INV_X1 aes_sbox_mult_msb_gf4_mul_1_1_U9 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n69), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n56) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U8 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_1_n54), .B(
        aes_sbox_mult_msb_gf4_mul_1_1_n70), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n55) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U7 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_1_n71), .A2(
        aes_sbox_mult_msb_gf4_mul_1_1_n72), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n54) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U5 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_1_n71), .A2(
        aes_sbox_mult_msb_gf4_mul_1_1_n69), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n67) );
  NOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U4 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_1_n72), .A2(
        aes_sbox_mult_msb_gf4_mul_1_1_n70), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n68) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U3 ( .A(aes_sbox_Y0_4xDP[4]), .B(
        aes_sbox_Y0_4xDP[6]), .ZN(aes_sbox_mult_msb_gf4_mul_1_1_n72) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_1_U2 ( .A(aes_sbox_Y0_4xDP[5]), .B(
        aes_sbox_Y0_4xDP[7]), .Z(aes_sbox_mult_msb_gf4_mul_1_1_n69) );
  OAI33_X1 aes_sbox_mult_msb_gf4_mul_1_1_U1 ( .A1(1'b0), .A2(
        aes_sbox_mult_msb_gf4_mul_1_1_n55), .A3(
        aes_sbox_mult_msb_gf4_mul_1_1_n56), .B1(
        aes_sbox_mult_msb_gf4_mul_1_1_n69), .B2(
        aes_sbox_mult_msb_gf4_mul_1_1_n72), .B3(
        aes_sbox_mult_msb_gf4_mul_1_1_n57), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_1_n77) );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_1_0_U28 ( .B1(aes_sbox_Y0_4xDP[2]), .B2(
        aes_sbox_Y0_4xDP[3]), .C1(aes_sbox_InverterOutxD_1__2_), .C2(
        aes_sbox_InverterOutxD_1__3_), .A(aes_sbox_mult_msb_gf4_mul_1_0_n73), 
        .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n75) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_1_0_U27 ( .A1(aes_sbox_Y0_4xDP[2]), .A2(
        aes_sbox_Y0_4xDP[3]), .B1(aes_sbox_InverterOutxD_1__3_), .B2(
        aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n73)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U26 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n63), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n62), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n74) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U25 ( .A(aes_sbox_InverterOutxD_1__1_), 
        .B(aes_sbox_InverterOutxD_1__3_), .Z(aes_sbox_mult_msb_gf4_mul_1_0_n67) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U24 ( .A(aes_sbox_InverterOutxD_1__0_), .B(aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n66) );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_1_0_U23 ( .B1(aes_sbox_Y0_4xDP[0]), .B2(
        aes_sbox_Y0_4xDP[1]), .C1(aes_sbox_InverterOutxD_1__0_), .C2(
        aes_sbox_InverterOutxD_1__1_), .A(aes_sbox_mult_msb_gf4_mul_1_0_n61), 
        .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n72) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_1_0_U22 ( .A1(aes_sbox_Y0_4xDP[0]), .A2(
        aes_sbox_Y0_4xDP[1]), .B1(aes_sbox_InverterOutxD_1__1_), .B2(
        aes_sbox_InverterOutxD_1__0_), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n61)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U21 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n59), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n60), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_2__3_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U20 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n76), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n75), .Z(
        aes_sbox_mult_msb_gf4_mul_1_0_n60) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U19 ( .A1(aes_sbox_Y0_4xDP[3]), .A2(
        aes_sbox_InverterOutxD_1__3_), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n59)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U18 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n57), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n58), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_2__2_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U17 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n74), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n75), .Z(
        aes_sbox_mult_msb_gf4_mul_1_0_n58) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U16 ( .A1(aes_sbox_Y0_4xDP[2]), .A2(
        aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n57)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U15 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n55), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n56), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_2__1_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U14 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n76), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n72), .Z(
        aes_sbox_mult_msb_gf4_mul_1_0_n56) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U13 ( .A1(aes_sbox_Y0_4xDP[1]), .A2(
        aes_sbox_InverterOutxD_1__1_), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n55)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U12 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n53), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n54), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_2__0_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U11 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n72), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n74), .Z(
        aes_sbox_mult_msb_gf4_mul_1_0_n54) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U10 ( .A1(aes_sbox_Y0_4xDP[0]), .A2(
        aes_sbox_InverterOutxD_1__0_), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n53)
         );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U9 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_0_n67), .A2(
        aes_sbox_mult_msb_gf4_mul_1_0_n69), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n65) );
  INV_X1 aes_sbox_mult_msb_gf4_mul_1_0_U8 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n64), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n71) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U7 ( .A(
        aes_sbox_mult_msb_gf4_mul_1_0_n66), .B(
        aes_sbox_mult_msb_gf4_mul_1_0_n65), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n70) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U6 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_0_n67), .A2(
        aes_sbox_mult_msb_gf4_mul_1_0_n71), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n68) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_1_0_U5 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_0_n71), .A2(
        aes_sbox_mult_msb_gf4_mul_1_0_n70), .B1(
        aes_sbox_mult_msb_gf4_mul_1_0_n69), .B2(
        aes_sbox_mult_msb_gf4_mul_1_0_n68), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n76) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U4 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_0_n67), .A2(
        aes_sbox_mult_msb_gf4_mul_1_0_n64), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n62) );
  NOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U3 ( .A1(
        aes_sbox_mult_msb_gf4_mul_1_0_n69), .A2(
        aes_sbox_mult_msb_gf4_mul_1_0_n66), .ZN(
        aes_sbox_mult_msb_gf4_mul_1_0_n63) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U2 ( .A(aes_sbox_Y0_4xDP[0]), .B(
        aes_sbox_Y0_4xDP[2]), .ZN(aes_sbox_mult_msb_gf4_mul_1_0_n69) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_1_0_U1 ( .A(aes_sbox_Y0_4xDP[1]), .B(
        aes_sbox_Y0_4xDP[3]), .Z(aes_sbox_mult_msb_gf4_mul_1_0_n64) );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_0_1_U29 ( .B1(aes_sbox_Y0_4xDP[6]), .B2(
        aes_sbox_Y0_4xDP[7]), .C1(aes_sbox_InverterOutxD_0__2_), .C2(
        aes_sbox_InverterOutxD_0__3_), .A(aes_sbox_mult_msb_gf4_mul_0_1_n74), 
        .ZN(aes_sbox_mult_msb_gf4_mul_0_1_n76) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_0_1_U28 ( .A1(aes_sbox_Y0_4xDP[6]), .A2(
        aes_sbox_Y0_4xDP[7]), .B1(aes_sbox_InverterOutxD_0__3_), .B2(
        aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_msb_gf4_mul_0_1_n74)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U27 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n68), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n67), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n75) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U26 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n65), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n66), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_1__1_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U25 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n77), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n73), .Z(
        aes_sbox_mult_msb_gf4_mul_0_1_n66) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U24 ( .A1(aes_sbox_Y0_4xDP[5]), .A2(
        aes_sbox_InverterOutxD_0__1_), .ZN(aes_sbox_mult_msb_gf4_mul_0_1_n65)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U23 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n63), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n64), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_1__3_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U22 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n77), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n76), .Z(
        aes_sbox_mult_msb_gf4_mul_0_1_n64) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U21 ( .A1(aes_sbox_Y0_4xDP[7]), .A2(
        aes_sbox_InverterOutxD_0__3_), .ZN(aes_sbox_mult_msb_gf4_mul_0_1_n63)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U20 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n61), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n62), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_1__2_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U19 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n75), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n76), .Z(
        aes_sbox_mult_msb_gf4_mul_0_1_n62) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U18 ( .A1(aes_sbox_Y0_4xDP[6]), .A2(
        aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_msb_gf4_mul_0_1_n61)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U17 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n59), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n60), .ZN(
        aes_sbox_mult_msb_Xi_mul_Yj_1__0_) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U16 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n73), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n75), .Z(
        aes_sbox_mult_msb_gf4_mul_0_1_n60) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U15 ( .A1(aes_sbox_Y0_4xDP[4]), .A2(
        aes_sbox_InverterOutxD_0__0_), .ZN(aes_sbox_mult_msb_gf4_mul_0_1_n59)
         );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_0_1_U14 ( .B1(
        aes_sbox_InverterOutxD_0__1_), .B2(aes_sbox_InverterOutxD_0__0_), .C1(
        aes_sbox_Y0_4xDP[5]), .C2(aes_sbox_Y0_4xDP[4]), .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n58), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n73) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_0_1_U13 ( .A1(
        aes_sbox_InverterOutxD_0__1_), .A2(aes_sbox_InverterOutxD_0__0_), .B1(
        aes_sbox_Y0_4xDP[4]), .B2(aes_sbox_Y0_4xDP[5]), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n58) );
  INV_X1 aes_sbox_mult_msb_gf4_mul_0_1_U12 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n71), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n57) );
  INV_X1 aes_sbox_mult_msb_gf4_mul_0_1_U11 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n69), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n56) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U10 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_1_n54), .B(
        aes_sbox_mult_msb_gf4_mul_0_1_n70), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n55) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U9 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_1_n71), .A2(
        aes_sbox_mult_msb_gf4_mul_0_1_n72), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n54) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U7 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_1_n71), .A2(
        aes_sbox_mult_msb_gf4_mul_0_1_n69), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n67) );
  NOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U6 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_1_n72), .A2(
        aes_sbox_mult_msb_gf4_mul_0_1_n70), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n68) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U5 ( .A(aes_sbox_InverterOutxD_0__1_), 
        .B(aes_sbox_InverterOutxD_0__3_), .Z(aes_sbox_mult_msb_gf4_mul_0_1_n71) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U4 ( .A(aes_sbox_InverterOutxD_0__0_), 
        .B(aes_sbox_InverterOutxD_0__2_), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n70) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U3 ( .A(aes_sbox_Y0_4xDP[4]), .B(
        aes_sbox_Y0_4xDP[6]), .ZN(aes_sbox_mult_msb_gf4_mul_0_1_n72) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_1_U2 ( .A(aes_sbox_Y0_4xDP[5]), .B(
        aes_sbox_Y0_4xDP[7]), .Z(aes_sbox_mult_msb_gf4_mul_0_1_n69) );
  OAI33_X1 aes_sbox_mult_msb_gf4_mul_0_1_U1 ( .A1(1'b0), .A2(
        aes_sbox_mult_msb_gf4_mul_0_1_n55), .A3(
        aes_sbox_mult_msb_gf4_mul_0_1_n56), .B1(
        aes_sbox_mult_msb_gf4_mul_0_1_n69), .B2(
        aes_sbox_mult_msb_gf4_mul_0_1_n72), .B3(
        aes_sbox_mult_msb_gf4_mul_0_1_n57), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_1_n77) );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_0_0_U28 ( .B1(aes_sbox_Y0_4xDP[2]), .B2(
        aes_sbox_Y0_4xDP[3]), .C1(aes_sbox_InverterOutxD_0__2_), .C2(
        aes_sbox_InverterOutxD_0__3_), .A(aes_sbox_mult_msb_gf4_mul_0_0_n73), 
        .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n75) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_0_0_U27 ( .A1(aes_sbox_Y0_4xDP[2]), .A2(
        aes_sbox_Y0_4xDP[3]), .B1(aes_sbox_InverterOutxD_0__3_), .B2(
        aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n73)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U26 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n63), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n62), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n74) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U25 ( .A(aes_sbox_InverterOutxD_0__1_), 
        .B(aes_sbox_InverterOutxD_0__3_), .Z(aes_sbox_mult_msb_gf4_mul_0_0_n67) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U24 ( .A(aes_sbox_InverterOutxD_0__0_), .B(aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n66) );
  AOI221_X1 aes_sbox_mult_msb_gf4_mul_0_0_U23 ( .B1(aes_sbox_Y0_4xDP[0]), .B2(
        aes_sbox_Y0_4xDP[1]), .C1(aes_sbox_InverterOutxD_0__0_), .C2(
        aes_sbox_InverterOutxD_0__1_), .A(aes_sbox_mult_msb_gf4_mul_0_0_n61), 
        .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n72) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_0_0_U22 ( .A1(aes_sbox_Y0_4xDP[0]), .A2(
        aes_sbox_Y0_4xDP[1]), .B1(aes_sbox_InverterOutxD_0__1_), .B2(
        aes_sbox_InverterOutxD_0__0_), .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n61)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U21 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n59), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n60), .ZN(aes_sbox_mult_msb_FFxDN[2]) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U20 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n75), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n74), .Z(
        aes_sbox_mult_msb_gf4_mul_0_0_n60) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U19 ( .A1(
        aes_sbox_InverterOutxD_0__2_), .A2(aes_sbox_Y0_4xDP[2]), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n59) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U18 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n57), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n58), .ZN(aes_sbox_mult_msb_FFxDN[3]) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U17 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n76), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n75), .Z(
        aes_sbox_mult_msb_gf4_mul_0_0_n58) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U16 ( .A1(aes_sbox_Y0_4xDP[3]), .A2(
        aes_sbox_InverterOutxD_0__3_), .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n57)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U15 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n55), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n56), .ZN(aes_sbox_mult_msb_FFxDN[1]) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U14 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n76), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n72), .Z(
        aes_sbox_mult_msb_gf4_mul_0_0_n56) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U13 ( .A1(aes_sbox_Y0_4xDP[1]), .A2(
        aes_sbox_InverterOutxD_0__1_), .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n55)
         );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U12 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n53), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n54), .ZN(aes_sbox_mult_msb_FFxDN[0]) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U11 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n72), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n74), .Z(
        aes_sbox_mult_msb_gf4_mul_0_0_n54) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U10 ( .A1(
        aes_sbox_InverterOutxD_0__0_), .A2(aes_sbox_Y0_4xDP[0]), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n53) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U9 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_0_n67), .A2(
        aes_sbox_mult_msb_gf4_mul_0_0_n69), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n65) );
  INV_X1 aes_sbox_mult_msb_gf4_mul_0_0_U8 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n64), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n71) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U7 ( .A(
        aes_sbox_mult_msb_gf4_mul_0_0_n66), .B(
        aes_sbox_mult_msb_gf4_mul_0_0_n65), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n70) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U6 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_0_n67), .A2(
        aes_sbox_mult_msb_gf4_mul_0_0_n71), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n68) );
  OAI22_X1 aes_sbox_mult_msb_gf4_mul_0_0_U5 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_0_n71), .A2(
        aes_sbox_mult_msb_gf4_mul_0_0_n70), .B1(
        aes_sbox_mult_msb_gf4_mul_0_0_n69), .B2(
        aes_sbox_mult_msb_gf4_mul_0_0_n68), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n76) );
  NAND2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U4 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_0_n67), .A2(
        aes_sbox_mult_msb_gf4_mul_0_0_n64), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n62) );
  NOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U3 ( .A1(
        aes_sbox_mult_msb_gf4_mul_0_0_n69), .A2(
        aes_sbox_mult_msb_gf4_mul_0_0_n66), .ZN(
        aes_sbox_mult_msb_gf4_mul_0_0_n63) );
  XNOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U2 ( .A(aes_sbox_Y0_4xDP[0]), .B(
        aes_sbox_Y0_4xDP[2]), .ZN(aes_sbox_mult_msb_gf4_mul_0_0_n69) );
  XOR2_X1 aes_sbox_mult_msb_gf4_mul_0_0_U1 ( .A(aes_sbox_Y0_4xDP[1]), .B(
        aes_sbox_Y0_4xDP[3]), .Z(aes_sbox_mult_msb_gf4_mul_0_0_n64) );
  XOR2_X1 aes_sbox_mult_lsb_U18 ( .A(aes_sbox_mult_lsb_n2), .B(
        aes_sbox_mult_lsb_n1), .Z(aes_sbox_InvUnmappedxD[11]) );
  XOR2_X1 aes_sbox_mult_lsb_U17 ( .A(aes_sbox_mult_lsb_n6), .B(
        aes_sbox_mult_lsb_n5), .Z(aes_sbox_InvUnmappedxD[9]) );
  XOR2_X1 aes_sbox_mult_lsb_U16 ( .A(aes_sbox_mult_lsb_n10), .B(
        aes_sbox_mult_lsb_n9), .Z(aes_sbox_InvUnmappedxD[3]) );
  XOR2_X1 aes_sbox_mult_lsb_U15 ( .A(aes_sbox_mult_lsb_n14), .B(
        aes_sbox_mult_lsb_n13), .Z(aes_sbox_InvUnmappedxD[1]) );
  XOR2_X1 aes_sbox_mult_lsb_U14 ( .A(aes_sbox_mult_lsb_n8), .B(
        aes_sbox_mult_lsb_n7), .Z(aes_sbox_InvUnmappedxD[8]) );
  XOR2_X1 aes_sbox_mult_lsb_U13 ( .A(Zmul3xDI[0]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__0_), .Z(aes_sbox_mult_lsb_FFxDN[4]) );
  XOR2_X1 aes_sbox_mult_lsb_U12 ( .A(aes_sbox_mult_lsb_n4), .B(
        aes_sbox_mult_lsb_n3), .Z(aes_sbox_InvUnmappedxD[10]) );
  XOR2_X1 aes_sbox_mult_lsb_U11 ( .A(aes_sbox_mult_lsb_n12), .B(
        aes_sbox_mult_lsb_n11), .Z(aes_sbox_InvUnmappedxD[2]) );
  XOR2_X1 aes_sbox_mult_lsb_U10 ( .A(Zmul3xDI[1]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__1_), .Z(aes_sbox_mult_lsb_FFxDN[5]) );
  XOR2_X1 aes_sbox_mult_lsb_U9 ( .A(aes_sbox_mult_lsb_n16), .B(
        aes_sbox_mult_lsb_n15), .Z(aes_sbox_InvUnmappedxD[0]) );
  XOR2_X1 aes_sbox_mult_lsb_U8 ( .A(Zmul3xDI[3]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__3_), .Z(aes_sbox_mult_lsb_FFxDN[11]) );
  XOR2_X1 aes_sbox_mult_lsb_U7 ( .A(Zmul3xDI[3]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__3_), .Z(aes_sbox_mult_lsb_FFxDN[7]) );
  XOR2_X1 aes_sbox_mult_lsb_U6 ( .A(Zmul3xDI[2]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__2_), .Z(aes_sbox_mult_lsb_FFxDN[10]) );
  XOR2_X1 aes_sbox_mult_lsb_U5 ( .A(Zmul3xDI[1]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__1_), .Z(aes_sbox_mult_lsb_FFxDN[9]) );
  XOR2_X1 aes_sbox_mult_lsb_U4 ( .A(Zmul3xDI[2]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__2_), .Z(aes_sbox_mult_lsb_FFxDN[6]) );
  XOR2_X1 aes_sbox_mult_lsb_U3 ( .A(Zmul3xDI[0]), .B(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__0_), .Z(aes_sbox_mult_lsb_FFxDN[8]) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_0__0_ ( .D(aes_sbox_mult_lsb_FFxDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n15) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_0__1_ ( .D(aes_sbox_mult_lsb_FFxDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n13) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_0__2_ ( .D(aes_sbox_mult_lsb_FFxDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n11) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_0__3_ ( .D(aes_sbox_mult_lsb_FFxDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n9) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_1__0_ ( .D(aes_sbox_mult_lsb_FFxDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n16) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_1__1_ ( .D(aes_sbox_mult_lsb_FFxDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n14) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_1__2_ ( .D(aes_sbox_mult_lsb_FFxDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n12) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_1__3_ ( .D(aes_sbox_mult_lsb_FFxDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n10) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_2__0_ ( .D(aes_sbox_mult_lsb_FFxDN[8]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n7) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_2__1_ ( .D(aes_sbox_mult_lsb_FFxDN[9]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n5) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_2__2_ ( .D(aes_sbox_mult_lsb_FFxDN[10]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n3) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_2__3_ ( .D(aes_sbox_mult_lsb_FFxDN[11]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n1) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_3__0_ ( .D(aes_sbox_mult_lsb_FFxDN[12]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n8) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_3__1_ ( .D(aes_sbox_mult_lsb_FFxDN[13]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n6) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_3__2_ ( .D(aes_sbox_mult_lsb_FFxDN[14]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n4) );
  DFFR_X1 aes_sbox_mult_lsb_FFxDP_reg_3__3_ ( .D(aes_sbox_mult_lsb_FFxDN[15]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(), .QN(aes_sbox_mult_lsb_n2) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U28 ( .B1(aes_sbox_Y1_4xDP[6]), .B2(
        aes_sbox_Y1_4xDP[7]), .C1(aes_sbox_InverterOutxD_1__2_), .C2(
        aes_sbox_InverterOutxD_1__3_), .A(aes_sbox_mult_lsb_gf4_mul_1_1_n73), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n75) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U27 ( .A1(aes_sbox_Y1_4xDP[6]), .A2(
        aes_sbox_Y1_4xDP[7]), .B1(aes_sbox_InverterOutxD_1__3_), .B2(
        aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n73)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U26 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n63), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n62), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n74) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U25 ( .A(aes_sbox_InverterOutxD_1__1_), 
        .B(aes_sbox_InverterOutxD_1__3_), .Z(aes_sbox_mult_lsb_gf4_mul_1_1_n67) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U24 ( .A(aes_sbox_InverterOutxD_1__0_), .B(aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n66) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U23 ( .B1(aes_sbox_Y1_4xDP[4]), .B2(
        aes_sbox_Y1_4xDP[5]), .C1(aes_sbox_InverterOutxD_1__0_), .C2(
        aes_sbox_InverterOutxD_1__1_), .A(aes_sbox_mult_lsb_gf4_mul_1_1_n61), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n72) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U22 ( .A1(aes_sbox_Y1_4xDP[4]), .A2(
        aes_sbox_Y1_4xDP[5]), .B1(aes_sbox_InverterOutxD_1__1_), .B2(
        aes_sbox_InverterOutxD_1__0_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n61)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U21 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n59), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n60), .ZN(aes_sbox_mult_lsb_FFxDN[15])
         );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U20 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n75), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_1_n60) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U19 ( .A1(aes_sbox_Y1_4xDP[7]), .A2(
        aes_sbox_InverterOutxD_1__3_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n59)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U18 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n57), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n58), .ZN(aes_sbox_mult_lsb_FFxDN[14])
         );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U17 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n75), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n74), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_1_n58) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U16 ( .A1(
        aes_sbox_InverterOutxD_1__2_), .A2(aes_sbox_Y1_4xDP[6]), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n57) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U15 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n55), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n56), .ZN(aes_sbox_mult_lsb_FFxDN[13])
         );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U14 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n72), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_1_n56) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U13 ( .A1(aes_sbox_Y1_4xDP[5]), .A2(
        aes_sbox_InverterOutxD_1__1_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n55)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U12 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n53), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n54), .ZN(aes_sbox_mult_lsb_FFxDN[12])
         );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U11 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n72), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n74), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_1_n54) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U10 ( .A1(
        aes_sbox_InverterOutxD_1__0_), .A2(aes_sbox_Y1_4xDP[4]), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n53) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U9 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_1_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_1_n69), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n65) );
  INV_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U8 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n71) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U7 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_1_n66), .B(
        aes_sbox_mult_lsb_gf4_mul_1_1_n65), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n70) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U6 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_1_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_1_n71), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n68) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U5 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_1_n71), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_1_n70), .B1(
        aes_sbox_mult_lsb_gf4_mul_1_1_n69), .B2(
        aes_sbox_mult_lsb_gf4_mul_1_1_n68), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n76) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U4 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_1_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_1_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n62) );
  NOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U3 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_1_n69), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_1_n66), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_1_n63) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U2 ( .A(aes_sbox_Y1_4xDP[4]), .B(
        aes_sbox_Y1_4xDP[6]), .ZN(aes_sbox_mult_lsb_gf4_mul_1_1_n69) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_1_U1 ( .A(aes_sbox_Y1_4xDP[5]), .B(
        aes_sbox_Y1_4xDP[7]), .Z(aes_sbox_mult_lsb_gf4_mul_1_1_n64) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U28 ( .B1(aes_sbox_Y1_4xDP[2]), .B2(
        aes_sbox_Y1_4xDP[3]), .C1(aes_sbox_InverterOutxD_1__2_), .C2(
        aes_sbox_InverterOutxD_1__3_), .A(aes_sbox_mult_lsb_gf4_mul_1_0_n73), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n75) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U27 ( .A1(aes_sbox_Y1_4xDP[2]), .A2(
        aes_sbox_Y1_4xDP[3]), .B1(aes_sbox_InverterOutxD_1__3_), .B2(
        aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n73)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U26 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n63), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n62), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n74) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U25 ( .A(aes_sbox_InverterOutxD_1__1_), 
        .B(aes_sbox_InverterOutxD_1__3_), .Z(aes_sbox_mult_lsb_gf4_mul_1_0_n67) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U24 ( .A(aes_sbox_InverterOutxD_1__0_), .B(aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n66) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U23 ( .B1(aes_sbox_Y1_4xDP[0]), .B2(
        aes_sbox_Y1_4xDP[1]), .C1(aes_sbox_InverterOutxD_1__0_), .C2(
        aes_sbox_InverterOutxD_1__1_), .A(aes_sbox_mult_lsb_gf4_mul_1_0_n61), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n72) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U22 ( .A1(aes_sbox_Y1_4xDP[0]), .A2(
        aes_sbox_Y1_4xDP[1]), .B1(aes_sbox_InverterOutxD_1__1_), .B2(
        aes_sbox_InverterOutxD_1__0_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n61)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U21 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n59), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n60), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__3_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U20 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n75), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_0_n60) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U19 ( .A1(aes_sbox_Y1_4xDP[3]), .A2(
        aes_sbox_InverterOutxD_1__3_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n59)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U18 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n57), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n58), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__2_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U17 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n74), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n75), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_0_n58) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U16 ( .A1(aes_sbox_Y1_4xDP[2]), .A2(
        aes_sbox_InverterOutxD_1__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n57)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U15 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n55), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n56), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__1_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U14 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n72), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_0_n56) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U13 ( .A1(aes_sbox_Y1_4xDP[1]), .A2(
        aes_sbox_InverterOutxD_1__1_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n55)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U12 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n53), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n54), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_2__0_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U11 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n72), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n74), .Z(
        aes_sbox_mult_lsb_gf4_mul_1_0_n54) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U10 ( .A1(aes_sbox_Y1_4xDP[0]), .A2(
        aes_sbox_InverterOutxD_1__0_), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n53)
         );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U9 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_0_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_0_n69), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n65) );
  INV_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U8 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n71) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U7 ( .A(
        aes_sbox_mult_lsb_gf4_mul_1_0_n66), .B(
        aes_sbox_mult_lsb_gf4_mul_1_0_n65), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n70) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U6 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_0_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_0_n71), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n68) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U5 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_0_n71), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_0_n70), .B1(
        aes_sbox_mult_lsb_gf4_mul_1_0_n69), .B2(
        aes_sbox_mult_lsb_gf4_mul_1_0_n68), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n76) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U4 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_0_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_0_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n62) );
  NOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U3 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_1_0_n69), .A2(
        aes_sbox_mult_lsb_gf4_mul_1_0_n66), .ZN(
        aes_sbox_mult_lsb_gf4_mul_1_0_n63) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U2 ( .A(aes_sbox_Y1_4xDP[0]), .B(
        aes_sbox_Y1_4xDP[2]), .ZN(aes_sbox_mult_lsb_gf4_mul_1_0_n69) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_1_0_U1 ( .A(aes_sbox_Y1_4xDP[1]), .B(
        aes_sbox_Y1_4xDP[3]), .Z(aes_sbox_mult_lsb_gf4_mul_1_0_n64) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U28 ( .B1(aes_sbox_Y1_4xDP[6]), .B2(
        aes_sbox_Y1_4xDP[7]), .C1(aes_sbox_InverterOutxD_0__2_), .C2(
        aes_sbox_InverterOutxD_0__3_), .A(aes_sbox_mult_lsb_gf4_mul_0_1_n73), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n75) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U27 ( .A1(aes_sbox_Y1_4xDP[6]), .A2(
        aes_sbox_Y1_4xDP[7]), .B1(aes_sbox_InverterOutxD_0__3_), .B2(
        aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n73)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U26 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n63), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n62), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n74) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U25 ( .A(aes_sbox_InverterOutxD_0__1_), 
        .B(aes_sbox_InverterOutxD_0__3_), .Z(aes_sbox_mult_lsb_gf4_mul_0_1_n67) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U24 ( .A(aes_sbox_InverterOutxD_0__0_), .B(aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n66) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U23 ( .B1(aes_sbox_Y1_4xDP[4]), .B2(
        aes_sbox_Y1_4xDP[5]), .C1(aes_sbox_InverterOutxD_0__0_), .C2(
        aes_sbox_InverterOutxD_0__1_), .A(aes_sbox_mult_lsb_gf4_mul_0_1_n61), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n72) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U22 ( .A1(aes_sbox_Y1_4xDP[4]), .A2(
        aes_sbox_Y1_4xDP[5]), .B1(aes_sbox_InverterOutxD_0__1_), .B2(
        aes_sbox_InverterOutxD_0__0_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n61)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U21 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n59), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n60), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__0_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U20 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n74), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n72), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_1_n60) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U19 ( .A1(aes_sbox_Y1_4xDP[4]), .A2(
        aes_sbox_InverterOutxD_0__0_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n59)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U18 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n57), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n58), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__1_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U17 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n72), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_1_n58) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U16 ( .A1(aes_sbox_Y1_4xDP[5]), .A2(
        aes_sbox_InverterOutxD_0__1_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n57)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U15 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n55), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n56), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__3_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U14 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n75), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_1_n56) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U13 ( .A1(aes_sbox_Y1_4xDP[7]), .A2(
        aes_sbox_InverterOutxD_0__3_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n55)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U12 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n53), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n54), .ZN(
        aes_sbox_mult_lsb_Xi_mul_Yj_1__2_) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U11 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n75), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n74), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_1_n54) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U10 ( .A1(aes_sbox_Y1_4xDP[6]), .A2(
        aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n53)
         );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U9 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_1_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_1_n69), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n65) );
  INV_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U8 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n71) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U7 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_1_n66), .B(
        aes_sbox_mult_lsb_gf4_mul_0_1_n65), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n70) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U6 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_1_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_1_n71), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n68) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U5 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_1_n71), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_1_n70), .B1(
        aes_sbox_mult_lsb_gf4_mul_0_1_n69), .B2(
        aes_sbox_mult_lsb_gf4_mul_0_1_n68), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n76) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U4 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_1_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_1_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n62) );
  NOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U3 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_1_n69), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_1_n66), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_1_n63) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U2 ( .A(aes_sbox_Y1_4xDP[4]), .B(
        aes_sbox_Y1_4xDP[6]), .ZN(aes_sbox_mult_lsb_gf4_mul_0_1_n69) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_1_U1 ( .A(aes_sbox_Y1_4xDP[5]), .B(
        aes_sbox_Y1_4xDP[7]), .Z(aes_sbox_mult_lsb_gf4_mul_0_1_n64) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U28 ( .B1(aes_sbox_Y1_4xDP[2]), .B2(
        aes_sbox_Y1_4xDP[3]), .C1(aes_sbox_InverterOutxD_0__2_), .C2(
        aes_sbox_InverterOutxD_0__3_), .A(aes_sbox_mult_lsb_gf4_mul_0_0_n73), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n75) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U27 ( .A1(aes_sbox_Y1_4xDP[2]), .A2(
        aes_sbox_Y1_4xDP[3]), .B1(aes_sbox_InverterOutxD_0__3_), .B2(
        aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n73)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U26 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n63), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n62), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n74) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U25 ( .A(aes_sbox_InverterOutxD_0__1_), 
        .B(aes_sbox_InverterOutxD_0__3_), .Z(aes_sbox_mult_lsb_gf4_mul_0_0_n67) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U24 ( .A(aes_sbox_InverterOutxD_0__0_), .B(aes_sbox_InverterOutxD_0__2_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n66) );
  AOI221_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U23 ( .B1(aes_sbox_Y1_4xDP[0]), .B2(
        aes_sbox_Y1_4xDP[1]), .C1(aes_sbox_InverterOutxD_0__0_), .C2(
        aes_sbox_InverterOutxD_0__1_), .A(aes_sbox_mult_lsb_gf4_mul_0_0_n61), 
        .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n72) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U22 ( .A1(aes_sbox_Y1_4xDP[0]), .A2(
        aes_sbox_Y1_4xDP[1]), .B1(aes_sbox_InverterOutxD_0__1_), .B2(
        aes_sbox_InverterOutxD_0__0_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n61)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U21 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n59), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n60), .ZN(aes_sbox_mult_lsb_FFxDN[3]) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U20 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n75), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_0_n60) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U19 ( .A1(aes_sbox_Y1_4xDP[3]), .A2(
        aes_sbox_InverterOutxD_0__3_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n59)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U18 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n57), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n58), .ZN(aes_sbox_mult_lsb_FFxDN[2]) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U17 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n75), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n74), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_0_n58) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U16 ( .A1(
        aes_sbox_InverterOutxD_0__2_), .A2(aes_sbox_Y1_4xDP[2]), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n57) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U15 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n55), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n56), .ZN(aes_sbox_mult_lsb_FFxDN[1]) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U14 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n76), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n72), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_0_n56) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U13 ( .A1(aes_sbox_Y1_4xDP[1]), .A2(
        aes_sbox_InverterOutxD_0__1_), .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n55)
         );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U12 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n53), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n54), .ZN(aes_sbox_mult_lsb_FFxDN[0]) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U11 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n72), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n74), .Z(
        aes_sbox_mult_lsb_gf4_mul_0_0_n54) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U10 ( .A1(
        aes_sbox_InverterOutxD_0__0_), .A2(aes_sbox_Y1_4xDP[0]), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n53) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U9 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_0_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_0_n69), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n65) );
  INV_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U8 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n71) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U7 ( .A(
        aes_sbox_mult_lsb_gf4_mul_0_0_n66), .B(
        aes_sbox_mult_lsb_gf4_mul_0_0_n65), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n70) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U6 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_0_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_0_n71), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n68) );
  OAI22_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U5 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_0_n71), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_0_n70), .B1(
        aes_sbox_mult_lsb_gf4_mul_0_0_n69), .B2(
        aes_sbox_mult_lsb_gf4_mul_0_0_n68), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n76) );
  NAND2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U4 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_0_n67), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_0_n64), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n62) );
  NOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U3 ( .A1(
        aes_sbox_mult_lsb_gf4_mul_0_0_n69), .A2(
        aes_sbox_mult_lsb_gf4_mul_0_0_n66), .ZN(
        aes_sbox_mult_lsb_gf4_mul_0_0_n63) );
  XNOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U2 ( .A(aes_sbox_Y1_4xDP[0]), .B(
        aes_sbox_Y1_4xDP[2]), .ZN(aes_sbox_mult_lsb_gf4_mul_0_0_n69) );
  XOR2_X1 aes_sbox_mult_lsb_gf4_mul_0_0_U1 ( .A(aes_sbox_Y1_4xDP[1]), .B(
        aes_sbox_Y1_4xDP[3]), .Z(aes_sbox_mult_lsb_gf4_mul_0_0_n64) );
  BUF_X1 aes_key_regs_1_U3 ( .A(n114), .Z(aes_key_regs_1_n4) );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_0_ ( .D(aes_key_regs_1_K00xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_0_ ( .D(aes_key_regs_1_K10xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_0_ ( .D(aes_key_regs_1_K20xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_0_ ( .D(aes_key_regs_1_K01xDP_0_), .SI(
        KeyOutxD[8]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_0_ ( .D(aes_key_regs_1_K01xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_0_ ( .D(aes_key_regs_1_K11xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_0_ ( .D(aes_key_regs_1_K21xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_0_ ( .D(aes_key_regs_1_K02xDP_0_), .SI(
        aes_key_regs_1_K01xDP_0_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_0_ ( .D(aes_key_regs_1_K02xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_0_ ( .D(aes_key_regs_1_K12xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_0_ ( .D(aes_key_regs_1_K22xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_0_ ( .D(K03xD[8]), .SI(
        aes_key_regs_1_K02xDP_0_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_1_ ( .D(aes_key_regs_1_K00xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_1_ ( .D(aes_key_regs_1_K10xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_1_ ( .D(aes_key_regs_1_K20xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_1_ ( .D(aes_key_regs_1_K01xDP_1_), .SI(
        KeyOutxD[9]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_1_ ( .D(aes_key_regs_1_K01xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_1_ ( .D(aes_key_regs_1_K11xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_1_ ( .D(aes_key_regs_1_K21xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_1_ ( .D(aes_key_regs_1_K02xDP_1_), .SI(
        aes_key_regs_1_K01xDP_1_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_1_ ( .D(aes_key_regs_1_K02xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_1_ ( .D(aes_key_regs_1_K12xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_1_ ( .D(aes_key_regs_1_K22xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_1_ ( .D(K03xD[9]), .SI(
        aes_key_regs_1_K02xDP_1_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_2_ ( .D(aes_key_regs_1_K00xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_2_ ( .D(aes_key_regs_1_K10xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_2_ ( .D(aes_key_regs_1_K20xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_2_ ( .D(aes_key_regs_1_K01xDP_2_), .SI(
        KeyOutxD[10]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_2_ ( .D(aes_key_regs_1_K01xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_2_ ( .D(aes_key_regs_1_K11xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_2_ ( .D(aes_key_regs_1_K21xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_2_ ( .D(aes_key_regs_1_K02xDP_2_), .SI(
        aes_key_regs_1_K01xDP_2_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_2_ ( .D(aes_key_regs_1_K02xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_2_ ( .D(aes_key_regs_1_K12xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_2_ ( .D(aes_key_regs_1_K22xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_2_ ( .D(K03xD[10]), .SI(
        aes_key_regs_1_K02xDP_2_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_3_ ( .D(aes_key_regs_1_K00xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_3_ ( .D(aes_key_regs_1_K10xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_3_ ( .D(aes_key_regs_1_K20xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_3_ ( .D(aes_key_regs_1_K01xDP_3_), .SI(
        KeyOutxD[11]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_3_ ( .D(aes_key_regs_1_K01xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_3_ ( .D(aes_key_regs_1_K11xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_3_ ( .D(aes_key_regs_1_K21xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_3_ ( .D(aes_key_regs_1_K02xDP_3_), .SI(
        aes_key_regs_1_K01xDP_3_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_3_ ( .D(aes_key_regs_1_K02xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_3_ ( .D(aes_key_regs_1_K12xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_3_ ( .D(aes_key_regs_1_K22xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_3_ ( .D(K03xD[11]), .SI(
        aes_key_regs_1_K02xDP_3_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_4_ ( .D(aes_key_regs_1_K00xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_4_ ( .D(aes_key_regs_1_K10xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_4_ ( .D(aes_key_regs_1_K20xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_4_ ( .D(aes_key_regs_1_K01xDP_4_), .SI(
        KeyOutxD[12]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_4_ ( .D(aes_key_regs_1_K01xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_4_ ( .D(aes_key_regs_1_K11xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_4_ ( .D(aes_key_regs_1_K21xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_4_ ( .D(aes_key_regs_1_K02xDP_4_), .SI(
        aes_key_regs_1_K01xDP_4_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_4_ ( .D(aes_key_regs_1_K02xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_4_ ( .D(aes_key_regs_1_K12xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_4_ ( .D(aes_key_regs_1_K22xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_4_ ( .D(K03xD[12]), .SI(
        aes_key_regs_1_K02xDP_4_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_5_ ( .D(aes_key_regs_1_K00xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_5_ ( .D(aes_key_regs_1_K10xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_5_ ( .D(aes_key_regs_1_K20xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_5_ ( .D(aes_key_regs_1_K01xDP_5_), .SI(
        KeyOutxD[13]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_5_ ( .D(aes_key_regs_1_K01xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_5_ ( .D(aes_key_regs_1_K11xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_5_ ( .D(aes_key_regs_1_K21xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_5_ ( .D(aes_key_regs_1_K02xDP_5_), .SI(
        aes_key_regs_1_K01xDP_5_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_5_ ( .D(aes_key_regs_1_K02xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_5_ ( .D(aes_key_regs_1_K12xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_5_ ( .D(aes_key_regs_1_K22xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_5_ ( .D(K03xD[13]), .SI(
        aes_key_regs_1_K02xDP_5_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K22xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_6_ ( .D(aes_key_regs_1_K00xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_6_ ( .D(aes_key_regs_1_K10xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_6_ ( .D(aes_key_regs_1_K20xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_6_ ( .D(aes_key_regs_1_K01xDP_6_), .SI(
        KeyOutxD[14]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K20xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_6_ ( .D(aes_key_regs_1_K01xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_6_ ( .D(aes_key_regs_1_K11xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_6_ ( .D(aes_key_regs_1_K21xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_6_ ( .D(aes_key_regs_1_K02xDP_6_), .SI(
        aes_key_regs_1_K01xDP_6_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K21xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_6_ ( .D(aes_key_regs_1_K02xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_6_ ( .D(aes_key_regs_1_K12xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_6_ ( .D(aes_key_regs_1_K22xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_6_ ( .D(K03xD[14]), .SI(
        aes_key_regs_1_K02xDP_6_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K00xDP_reg_7_ ( .D(aes_key_regs_1_K00xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K10xDP_reg_7_ ( .D(aes_key_regs_1_K10xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K00xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K20xDP_reg_7_ ( .D(aes_key_regs_1_K20xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K10xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K30xDP_reg_7_ ( .D(aes_key_regs_1_K01xDP_7_), .SI(
        KeyOutxD[15]), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K20xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K01xDP_reg_7_ ( .D(aes_key_regs_1_K01xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_1_K11xDP_reg_7_ ( .D(aes_key_regs_1_K11xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K01xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K21xDP_reg_7_ ( .D(aes_key_regs_1_K21xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K11xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K31xDP_reg_7_ ( .D(aes_key_regs_1_K02xDP_7_), .SI(
        aes_key_regs_1_K01xDP_7_), .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_1_K21xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K02xDP_reg_7_ ( .D(aes_key_regs_1_K02xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_1_K12xDP_reg_7_ ( .D(aes_key_regs_1_K12xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K02xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K22xDP_reg_7_ ( .D(aes_key_regs_1_K22xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K12xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K32xDP_reg_7_ ( .D(K03xD[15]), .SI(
        aes_key_regs_1_K02xDP_7_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_1_K22xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_0_ ( .D(KeyInxD[8]), .SI(K03xD[8]), .SE(
        aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_0_ ( .D(KeyToSboxOutxD[8]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_0_ ( .D(aes_key_regs_1_K13xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[8]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_0_ ( .D(aes_key_regs_1_K23xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_1_ ( .D(KeyInxD[9]), .SI(K03xD[9]), .SE(
        aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_1_ ( .D(KeyToSboxOutxD[9]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_1_ ( .D(aes_key_regs_1_K13xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[9]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_1_ ( .D(aes_key_regs_1_K23xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_2_ ( .D(KeyInxD[10]), .SI(K03xD[10]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_2_ ( .D(KeyToSboxOutxD[10]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_2_ ( .D(aes_key_regs_1_K13xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[10]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_2_ ( .D(aes_key_regs_1_K23xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_3_ ( .D(KeyInxD[11]), .SI(K03xD[11]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_3_ ( .D(KeyToSboxOutxD[11]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_3_ ( .D(aes_key_regs_1_K13xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[11]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_3_ ( .D(aes_key_regs_1_K23xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_4_ ( .D(KeyInxD[12]), .SI(K03xD[12]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_4_ ( .D(KeyToSboxOutxD[12]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_4_ ( .D(aes_key_regs_1_K13xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[12]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_4_ ( .D(aes_key_regs_1_K23xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_5_ ( .D(KeyInxD[13]), .SI(K03xD[13]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_5_ ( .D(KeyToSboxOutxD[13]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_5_ ( .D(aes_key_regs_1_K13xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[13]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_5_ ( .D(aes_key_regs_1_K23xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_6_ ( .D(KeyInxD[14]), .SI(K03xD[14]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_6_ ( .D(KeyToSboxOutxD[14]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_6_ ( .D(aes_key_regs_1_K13xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[14]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_6_ ( .D(aes_key_regs_1_K23xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_1_K33xDP_reg_7_ ( .D(KeyInxD[15]), .SI(K03xD[15]), 
        .SE(aes_key_regs_1_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_1_K23xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_1_K03xDP_reg_7_ ( .D(KeyToSboxOutxD[15]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K13xDP_reg_7_ ( .D(aes_key_regs_1_K13xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[15]), .QN() );
  DFFR_X1 aes_key_regs_1_K23xDP_reg_7_ ( .D(aes_key_regs_1_K23xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_1_K13xDN[7]), .QN() );
  INV_X1 aes_state_regs_1_U56 ( .A(aes_state_regs_1_MixColumnsS2xD[7]), .ZN(
        aes_state_regs_1_n80) );
  INV_X1 aes_state_regs_1_U55 ( .A(aes_state_regs_1_MixColumnsS2xD[6]), .ZN(
        aes_state_regs_1_n79) );
  INV_X1 aes_state_regs_1_U54 ( .A(aes_state_regs_1_MixColumnsS2xD[5]), .ZN(
        aes_state_regs_1_n78) );
  INV_X1 aes_state_regs_1_U53 ( .A(aes_state_regs_1_MixColumnsS2xD[4]), .ZN(
        aes_state_regs_1_n77) );
  INV_X1 aes_state_regs_1_U52 ( .A(aes_state_regs_1_MixColumnsS2xD[3]), .ZN(
        aes_state_regs_1_n76) );
  INV_X1 aes_state_regs_1_U51 ( .A(aes_state_regs_1_MixColumnsS2xD[2]), .ZN(
        aes_state_regs_1_n75) );
  INV_X2 aes_state_regs_1_U50 ( .A(aes_state_regs_1_n74), .ZN(
        aes_state_regs_1_n73) );
  INV_X2 aes_state_regs_1_U49 ( .A(aes_state_regs_1_n74), .ZN(
        aes_state_regs_1_n72) );
  OAI222_X1 aes_state_regs_1_U48 ( .A1(aes_state_regs_1_n69), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n62), .C1(aes_state_regs_1_n81), .C2(
        aes_state_regs_1_n97), .ZN(aes_state_regs_1_S20xDN[0]) );
  INV_X1 aes_state_regs_1_U47 ( .A(aes_state_regs_1_MixColumnsS3xD[0]), .ZN(
        aes_state_regs_1_n69) );
  OAI222_X1 aes_state_regs_1_U46 ( .A1(aes_state_regs_1_n68), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n60), .C1(aes_state_regs_1_n81), .C2(
        aes_state_regs_1_n95), .ZN(aes_state_regs_1_S20xDN[2]) );
  INV_X1 aes_state_regs_1_U45 ( .A(aes_state_regs_1_MixColumnsS3xD[2]), .ZN(
        aes_state_regs_1_n68) );
  OAI222_X1 aes_state_regs_1_U44 ( .A1(aes_state_regs_1_n67), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n54), .C1(aes_state_regs_1_n105), .C2(
        aes_state_regs_1_n81), .ZN(aes_state_regs_1_S10xDN[0]) );
  INV_X1 aes_state_regs_1_U43 ( .A(aes_state_regs_1_MixColumnsS2xD[0]), .ZN(
        aes_state_regs_1_n67) );
  OAI21_X1 aes_state_regs_1_U42 ( .B1(aes_state_regs_1_n91), .B2(
        aes_state_regs_1_n81), .A(aes_state_regs_1_n66), .ZN(
        aes_state_regs_1_S20xDN[6]) );
  AOI22_X1 aes_state_regs_1_U41 ( .A1(aes_state_regs_1_MixColumnsS3xD[6]), 
        .A2(aes_state_regs_1_n70), .B1(aes_state_regs_1_n8), .B2(
        aes_state_regs_1_n73), .ZN(aes_state_regs_1_n66) );
  OAI222_X1 aes_state_regs_1_U40 ( .A1(aes_state_regs_1_n65), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n61), .C1(aes_state_regs_1_n81), .C2(
        aes_state_regs_1_n96), .ZN(aes_state_regs_1_S20xDN[1]) );
  INV_X1 aes_state_regs_1_U39 ( .A(aes_state_regs_1_MixColumnsS3xD[1]), .ZN(
        aes_state_regs_1_n65) );
  OAI222_X1 aes_state_regs_1_U38 ( .A1(aes_state_regs_1_n64), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n59), .C1(aes_state_regs_1_n81), .C2(
        aes_state_regs_1_n94), .ZN(aes_state_regs_1_S20xDN[3]) );
  INV_X1 aes_state_regs_1_U37 ( .A(aes_state_regs_1_MixColumnsS3xD[3]), .ZN(
        aes_state_regs_1_n64) );
  OAI222_X1 aes_state_regs_1_U36 ( .A1(aes_state_regs_1_n63), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n53), .C1(aes_state_regs_1_n104), .C2(
        aes_state_regs_1_n81), .ZN(aes_state_regs_1_S10xDN[1]) );
  INV_X1 aes_state_regs_1_U35 ( .A(aes_state_regs_1_MixColumnsS2xD[1]), .ZN(
        aes_state_regs_1_n63) );
  OAI222_X1 aes_state_regs_1_U34 ( .A1(aes_state_regs_1_n56), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n55), .C1(aes_state_regs_1_n81), .C2(
        aes_state_regs_1_n90), .ZN(aes_state_regs_1_S20xDN[7]) );
  INV_X1 aes_state_regs_1_U33 ( .A(aes_state_regs_1_MixColumnsS3xD[7]), .ZN(
        aes_state_regs_1_n56) );
  OAI222_X1 aes_state_regs_1_U32 ( .A1(aes_state_regs_1_n46), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n58), .C1(aes_state_regs_1_n81), .C2(
        aes_state_regs_1_n93), .ZN(aes_state_regs_1_S20xDN[4]) );
  INV_X1 aes_state_regs_1_U31 ( .A(aes_state_regs_1_MixColumnsS3xD[4]), .ZN(
        aes_state_regs_1_n46) );
  OAI222_X1 aes_state_regs_1_U30 ( .A1(aes_state_regs_1_n45), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n74), .B2(
        aes_state_regs_1_n57), .C1(aes_state_regs_1_n81), .C2(
        aes_state_regs_1_n92), .ZN(aes_state_regs_1_S20xDN[5]) );
  INV_X1 aes_state_regs_1_U29 ( .A(aes_state_regs_1_MixColumnsS3xD[5]), .ZN(
        aes_state_regs_1_n45) );
  INV_X2 aes_state_regs_1_U28 ( .A(aes_state_regs_1_n70), .ZN(
        aes_state_regs_1_n71) );
  OAI222_X1 aes_state_regs_1_U27 ( .A1(aes_state_regs_1_n75), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n81), .B2(
        aes_state_regs_1_n103), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n52), .ZN(aes_state_regs_1_S10xDN[2]) );
  OAI222_X1 aes_state_regs_1_U26 ( .A1(aes_state_regs_1_n76), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n81), .B2(
        aes_state_regs_1_n102), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n51), .ZN(aes_state_regs_1_S10xDN[3]) );
  OAI222_X1 aes_state_regs_1_U25 ( .A1(aes_state_regs_1_n77), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n81), .B2(
        aes_state_regs_1_n101), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n50), .ZN(aes_state_regs_1_S10xDN[4]) );
  OAI222_X1 aes_state_regs_1_U24 ( .A1(aes_state_regs_1_n78), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n81), .B2(
        aes_state_regs_1_n100), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n49), .ZN(aes_state_regs_1_S10xDN[5]) );
  OAI222_X1 aes_state_regs_1_U23 ( .A1(aes_state_regs_1_n79), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n81), .B2(
        aes_state_regs_1_n99), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n48), .ZN(aes_state_regs_1_S10xDN[6]) );
  OAI222_X1 aes_state_regs_1_U22 ( .A1(aes_state_regs_1_n80), .A2(
        aes_state_regs_1_n71), .B1(aes_state_regs_1_n81), .B2(
        aes_state_regs_1_n98), .C1(aes_state_regs_1_n74), .C2(
        aes_state_regs_1_n47), .ZN(aes_state_regs_1_S10xDN[7]) );
  NAND2_X1 aes_state_regs_1_U21 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[7]), .ZN(aes_state_regs_1_n106) );
  OAI21_X1 aes_state_regs_1_U20 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n82), .A(aes_state_regs_1_n106), .ZN(StateOutxD[15])
         );
  NAND2_X1 aes_state_regs_1_U19 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[4]), .ZN(aes_state_regs_1_n109) );
  OAI21_X1 aes_state_regs_1_U18 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n86), .A(aes_state_regs_1_n109), .ZN(StateOutxD[12])
         );
  NAND2_X1 aes_state_regs_1_U17 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[3]), .ZN(aes_state_regs_1_n110) );
  OAI21_X1 aes_state_regs_1_U16 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n85), .A(aes_state_regs_1_n110), .ZN(StateOutxD[11])
         );
  NAND2_X1 aes_state_regs_1_U15 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[2]), .ZN(aes_state_regs_1_n111) );
  OAI21_X1 aes_state_regs_1_U14 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n84), .A(aes_state_regs_1_n111), .ZN(StateOutxD[10])
         );
  OAI21_X1 aes_state_regs_1_U13 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n83), .A(aes_state_regs_1_n112), .ZN(StateOutxD[9])
         );
  NAND2_X1 aes_state_regs_1_U12 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[0]), .ZN(aes_state_regs_1_n113) );
  OAI21_X1 aes_state_regs_1_U11 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n89), .A(aes_state_regs_1_n113), .ZN(StateOutxD[8])
         );
  INV_X1 aes_state_regs_1_U10 ( .A(nextRCONxS), .ZN(aes_state_regs_1_n74) );
  OR2_X1 aes_state_regs_1_U9 ( .A1(aes_state_regs_1_n73), .A2(doMixColumnsxS), 
        .ZN(aes_state_regs_1_n81) );
  AND2_X2 aes_state_regs_1_U8 ( .A1(doMixColumnsxS), .A2(aes_state_regs_1_n74), 
        .ZN(aes_state_regs_1_n70) );
  NAND2_X1 aes_state_regs_1_U7 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[6]), .ZN(aes_state_regs_1_n107) );
  OAI21_X1 aes_state_regs_1_U6 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n88), .A(aes_state_regs_1_n107), .ZN(StateOutxD[14])
         );
  NAND2_X1 aes_state_regs_1_U5 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[5]), .ZN(aes_state_regs_1_n108) );
  OAI21_X1 aes_state_regs_1_U4 ( .B1(aes_state_regs_1_n70), .B2(
        aes_state_regs_1_n87), .A(aes_state_regs_1_n108), .ZN(StateOutxD[13])
         );
  NAND2_X1 aes_state_regs_1_U3 ( .A1(aes_state_regs_1_n70), .A2(
        aes_state_regs_1_MixColumnsS0xD[1]), .ZN(aes_state_regs_1_n112) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_7_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[7]), .SI(aes_state_regs_1_S10xDP_7_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[7]), .QN(aes_state_regs_1_n82) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_6_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[6]), .SI(aes_state_regs_1_S10xDP_6_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[6]), .QN(aes_state_regs_1_n88) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_5_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[5]), .SI(aes_state_regs_1_S10xDP_5_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[5]), .QN(aes_state_regs_1_n87) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_4_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[4]), .SI(aes_state_regs_1_S10xDP_4_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[4]), .QN(aes_state_regs_1_n86) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_3_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[3]), .SI(aes_state_regs_1_S10xDP_3_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[3]), .QN(aes_state_regs_1_n85) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_2_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[2]), .SI(aes_state_regs_1_S10xDP_2_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[2]), .QN(aes_state_regs_1_n84) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_1_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[1]), .SI(aes_state_regs_1_S10xDP_1_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[1]), .QN(aes_state_regs_1_n83) );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_7_ ( .D(aes_state_regs_1_S10xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_7_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_6_ ( .D(aes_state_regs_1_S10xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_6_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_5_ ( .D(aes_state_regs_1_S10xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_5_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_4_ ( .D(aes_state_regs_1_S10xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_4_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_3_ ( .D(aes_state_regs_1_S10xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_3_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_2_ ( .D(aes_state_regs_1_S10xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_2_), .QN() );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_1_ ( .D(aes_state_regs_1_S10xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_7_ ( .D(aes_state_regs_1_S01xDO_7_), 
        .SI(StateInxD[15]), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_7_), .QN(aes_state_regs_1_n90) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_7_ ( .D(aes_state_regs_1_n1), .SI(
        aes_state_regs_1_n4), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[7]), .QN(aes_state_regs_1_n47) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_7_ ( .D(aes_state_regs_1_S02xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_7_ ( .D(aes_state_regs_1_n2), .SI(
        aes_state_regs_1_S23xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_7_ ( .D(aes_state_regs_1_n4), .SI(
        aes_state_regs_1_n1), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_7_ ( .D(aes_state_regs_1_S02xDP_7_), 
        .SI(aes_state_regs_1_S01xDO_7_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n1), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_7_ ( .D(aes_state_regs_1_S01xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_7_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_7_ ( .D(aes_state_regs_1_S21xDP[7]), 
        .SI(aes_state_regs_1_n2), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S01xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_7_ ( .D(aes_state_regs_1_n3), .SI(
        aes_state_regs_1_S30xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n2), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_7_ ( .D(aes_state_regs_1_n5), .SI(
        aes_state_regs_1_S02xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n3), .QN(aes_state_regs_1_n55) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_7_ ( .D(StateInxD[15]), .SI(
        aes_state_regs_1_n5), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n4), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_7_ ( .D(aes_state_regs_1_S03xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n5), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_7_ ( .D(aes_state_regs_1_S23xDP_7_), 
        .SI(aes_state_regs_1_S20xDP_7_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[7]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_7_ ( .D(aes_state_regs_1_S20xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_7_), .QN(
        aes_state_regs_1_n98) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_6_ ( .D(aes_state_regs_1_S01xDO_6_), 
        .SI(StateInxD[14]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_6_), .QN(aes_state_regs_1_n91) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_6_ ( .D(aes_state_regs_1_n6), .SI(
        aes_state_regs_1_n9), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[6]), .QN(aes_state_regs_1_n48) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_6_ ( .D(aes_state_regs_1_S02xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_6_ ( .D(aes_state_regs_1_n7), .SI(
        aes_state_regs_1_S23xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_6_ ( .D(aes_state_regs_1_n9), .SI(
        aes_state_regs_1_n6), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_6_ ( .D(aes_state_regs_1_S02xDP_6_), 
        .SI(aes_state_regs_1_S01xDO_6_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n6), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_6_ ( .D(aes_state_regs_1_S01xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_6_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_6_ ( .D(aes_state_regs_1_S21xDP[6]), 
        .SI(aes_state_regs_1_n7), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S01xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_6_ ( .D(aes_state_regs_1_n8), .SI(
        aes_state_regs_1_S30xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n7), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_6_ ( .D(aes_state_regs_1_n10), .SI(
        aes_state_regs_1_S02xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n8), .QN() );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_6_ ( .D(StateInxD[14]), .SI(
        aes_state_regs_1_n10), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n9), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_6_ ( .D(aes_state_regs_1_S03xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n10), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_6_ ( .D(aes_state_regs_1_S23xDP_6_), 
        .SI(aes_state_regs_1_S20xDP_6_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[6]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_6_ ( .D(aes_state_regs_1_S20xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_6_), .QN(
        aes_state_regs_1_n99) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_5_ ( .D(aes_state_regs_1_S01xDO_5_), 
        .SI(StateInxD[13]), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_5_), .QN(aes_state_regs_1_n92) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_5_ ( .D(aes_state_regs_1_n11), .SI(
        aes_state_regs_1_n14), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[5]), .QN(aes_state_regs_1_n49) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_5_ ( .D(aes_state_regs_1_S02xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_5_ ( .D(aes_state_regs_1_n12), .SI(
        aes_state_regs_1_S23xDP_5_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_5_ ( .D(aes_state_regs_1_n14), .SI(
        aes_state_regs_1_n11), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_5_ ( .D(aes_state_regs_1_S02xDP_5_), 
        .SI(aes_state_regs_1_S01xDO_5_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n11), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_5_ ( .D(aes_state_regs_1_S01xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_5_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_5_ ( .D(aes_state_regs_1_S21xDP[5]), 
        .SI(aes_state_regs_1_n12), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_5_ ( .D(aes_state_regs_1_n13), .SI(
        aes_state_regs_1_S30xDP_5_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n12), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_5_ ( .D(aes_state_regs_1_n15), .SI(
        aes_state_regs_1_S02xDP_5_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n13), .QN(aes_state_regs_1_n57) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_5_ ( .D(StateInxD[13]), .SI(
        aes_state_regs_1_n15), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n14), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_5_ ( .D(aes_state_regs_1_S03xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n15), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_5_ ( .D(aes_state_regs_1_S23xDP_5_), 
        .SI(aes_state_regs_1_S20xDP_5_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[5]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_5_ ( .D(aes_state_regs_1_S20xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_5_), .QN(
        aes_state_regs_1_n100) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_4_ ( .D(aes_state_regs_1_S01xDO_4_), 
        .SI(StateInxD[12]), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_4_), .QN(aes_state_regs_1_n93) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_4_ ( .D(aes_state_regs_1_n16), .SI(
        aes_state_regs_1_n19), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[4]), .QN(aes_state_regs_1_n50) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_4_ ( .D(aes_state_regs_1_S02xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_4_ ( .D(aes_state_regs_1_n17), .SI(
        aes_state_regs_1_S23xDP_4_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_4_ ( .D(aes_state_regs_1_n19), .SI(
        aes_state_regs_1_n16), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_4_ ( .D(aes_state_regs_1_S02xDP_4_), 
        .SI(aes_state_regs_1_S01xDO_4_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n16), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_4_ ( .D(aes_state_regs_1_S01xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_4_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_4_ ( .D(aes_state_regs_1_S21xDP[4]), 
        .SI(aes_state_regs_1_n17), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_4_ ( .D(aes_state_regs_1_n18), .SI(
        aes_state_regs_1_S30xDP_4_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n17), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_4_ ( .D(aes_state_regs_1_n20), .SI(
        aes_state_regs_1_S02xDP_4_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n18), .QN(aes_state_regs_1_n58) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_4_ ( .D(StateInxD[12]), .SI(
        aes_state_regs_1_n20), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n19), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_4_ ( .D(aes_state_regs_1_S03xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n20), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_4_ ( .D(aes_state_regs_1_S23xDP_4_), 
        .SI(aes_state_regs_1_S20xDP_4_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[4]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_4_ ( .D(aes_state_regs_1_S20xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_4_), .QN(
        aes_state_regs_1_n101) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_3_ ( .D(aes_state_regs_1_S01xDO_3_), 
        .SI(StateInxD[11]), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_3_), .QN(aes_state_regs_1_n94) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_3_ ( .D(aes_state_regs_1_n21), .SI(
        aes_state_regs_1_n24), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[3]), .QN(aes_state_regs_1_n51) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_3_ ( .D(aes_state_regs_1_S02xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_3_ ( .D(aes_state_regs_1_n22), .SI(
        aes_state_regs_1_S23xDP_3_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_3_ ( .D(aes_state_regs_1_n24), .SI(
        aes_state_regs_1_n21), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_3_ ( .D(aes_state_regs_1_S02xDP_3_), 
        .SI(aes_state_regs_1_S01xDO_3_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n21), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_3_ ( .D(aes_state_regs_1_S01xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_3_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_3_ ( .D(aes_state_regs_1_S21xDP[3]), 
        .SI(aes_state_regs_1_n22), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_3_ ( .D(aes_state_regs_1_n23), .SI(
        aes_state_regs_1_S30xDP_3_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n22), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_3_ ( .D(aes_state_regs_1_n25), .SI(
        aes_state_regs_1_S02xDP_3_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n23), .QN(aes_state_regs_1_n59) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_3_ ( .D(StateInxD[11]), .SI(
        aes_state_regs_1_n25), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n24), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_3_ ( .D(aes_state_regs_1_S03xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n25), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_3_ ( .D(aes_state_regs_1_S23xDP_3_), 
        .SI(aes_state_regs_1_S20xDP_3_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[3]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_3_ ( .D(aes_state_regs_1_S20xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_3_), .QN(
        aes_state_regs_1_n102) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_2_ ( .D(aes_state_regs_1_S01xDO_2_), 
        .SI(StateInxD[10]), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S30xDP_2_), .QN(aes_state_regs_1_n95) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_2_ ( .D(aes_state_regs_1_n26), .SI(
        aes_state_regs_1_n29), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[2]), .QN(aes_state_regs_1_n52) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_2_ ( .D(aes_state_regs_1_S02xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_2_ ( .D(aes_state_regs_1_n27), .SI(
        aes_state_regs_1_S23xDP_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_2_ ( .D(aes_state_regs_1_n29), .SI(
        aes_state_regs_1_n26), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_2_ ( .D(aes_state_regs_1_S02xDP_2_), 
        .SI(aes_state_regs_1_S01xDO_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n26), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_2_ ( .D(aes_state_regs_1_S01xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_2_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_2_ ( .D(aes_state_regs_1_S21xDP[2]), 
        .SI(aes_state_regs_1_n27), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_2_ ( .D(aes_state_regs_1_n28), .SI(
        aes_state_regs_1_S30xDP_2_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n27), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_2_ ( .D(aes_state_regs_1_n30), .SI(
        aes_state_regs_1_S02xDP_2_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n28), .QN(aes_state_regs_1_n60) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_2_ ( .D(StateInxD[10]), .SI(
        aes_state_regs_1_n30), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n29), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_2_ ( .D(aes_state_regs_1_S03xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n30), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_2_ ( .D(aes_state_regs_1_S23xDP_2_), 
        .SI(aes_state_regs_1_S20xDP_2_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[2]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_2_ ( .D(aes_state_regs_1_S20xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_2_), .QN(
        aes_state_regs_1_n103) );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_1_ ( .D(aes_state_regs_1_S01xDO_1_), 
        .SI(StateInxD[9]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), 
        .Q(aes_state_regs_1_S30xDP_1_), .QN(aes_state_regs_1_n96) );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_1_ ( .D(aes_state_regs_1_n31), .SI(
        aes_state_regs_1_n34), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S21xDP[1]), .QN(aes_state_regs_1_n53) );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_1_ ( .D(aes_state_regs_1_S02xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_1_ ( .D(aes_state_regs_1_n32), .SI(
        aes_state_regs_1_S23xDP_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_1_ ( .D(aes_state_regs_1_n34), .SI(
        aes_state_regs_1_n31), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_S23xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_1_ ( .D(aes_state_regs_1_S02xDP_1_), 
        .SI(aes_state_regs_1_S01xDO_1_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n31), .QN() );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_1_ ( .D(aes_state_regs_1_S01xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_1_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_1_ ( .D(aes_state_regs_1_S21xDP[1]), 
        .SI(aes_state_regs_1_n32), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_1_ ( .D(aes_state_regs_1_n33), .SI(
        aes_state_regs_1_S30xDP_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n32), .QN() );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_1_ ( .D(aes_state_regs_1_n35), .SI(
        aes_state_regs_1_S02xDP_1_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n33), .QN(aes_state_regs_1_n61) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_1_ ( .D(StateInxD[9]), .SI(
        aes_state_regs_1_n35), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_1_n34), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_1_ ( .D(aes_state_regs_1_S03xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n35), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_1_ ( .D(aes_state_regs_1_S23xDP_1_), 
        .SI(aes_state_regs_1_S20xDP_1_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[1]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_1_ ( .D(aes_state_regs_1_S20xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_1_), .QN(
        aes_state_regs_1_n104) );
  SDFFR_X1 aes_state_regs_1_S00xDP_reg_0_ ( .D(
        aes_state_regs_1_MixColumnsS1xD[0]), .SI(aes_state_regs_1_S10xDP_0_), 
        .SE(aes_state_regs_1_n71), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_1_S00xDP[0]), .QN(aes_state_regs_1_n89) );
  DFFR_X1 aes_state_regs_1_S10xDP_reg_0_ ( .D(aes_state_regs_1_S10xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S10xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S23xDP_reg_0_ ( .D(aes_state_regs_1_n37), .SI(
        aes_state_regs_1_S31xDP_0_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S23xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S31xDP_reg_0_ ( .D(aes_state_regs_1_S02xDP_0_), 
        .SI(aes_state_regs_1_S01xDO_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S31xDP_0_), .QN() );
  DFFR_X1 aes_state_regs_1_S02xDP_reg_0_ ( .D(aes_state_regs_1_S02xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S12xDP_reg_0_ ( .D(aes_state_regs_1_S22xDP_0_), 
        .SI(aes_state_regs_1_S23xDP_0_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S02xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_1_S22xDP_reg_0_ ( .D(aes_state_regs_1_n38), .SI(
        aes_state_regs_1_S30xDP_0_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S22xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S30xDP_reg_0_ ( .D(aes_state_regs_1_S01xDO_0_), 
        .SI(StateInxD[8]), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), 
        .Q(aes_state_regs_1_S30xDP_0_), .QN(aes_state_regs_1_n97) );
  DFFR_X1 aes_state_regs_1_S01xDP_reg_0_ ( .D(aes_state_regs_1_S01xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S01xDO_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S11xDP_reg_0_ ( .D(aes_state_regs_1_n36), .SI(
        aes_state_regs_1_S22xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_S01xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_1_S21xDP_reg_0_ ( .D(aes_state_regs_1_S31xDP_0_), 
        .SI(aes_state_regs_1_n37), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n36), .QN(aes_state_regs_1_n54) );
  SDFFR_X1 aes_state_regs_1_S33xDP_reg_0_ ( .D(StateInxD[8]), .SI(
        aes_state_regs_1_S03xDP_0_), .SE(aes_state_regs_1_n72), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_1_n37), .QN() );
  DFFR_X1 aes_state_regs_1_S03xDP_reg_0_ ( .D(aes_state_regs_1_S03xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_1_S13xDP_reg_0_ ( .D(aes_state_regs_1_S23xDP_0_), 
        .SI(aes_state_regs_1_S20xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S03xDN[0]), .QN() );
  DFFR_X1 aes_state_regs_1_S20xDP_reg_0_ ( .D(aes_state_regs_1_S20xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_S20xDP_0_), .QN(
        aes_state_regs_1_n105) );
  SDFFR_X1 aes_state_regs_1_S32xDP_reg_0_ ( .D(aes_state_regs_1_S03xDP_0_), 
        .SI(aes_state_regs_1_S02xDP_0_), .SE(aes_state_regs_1_n73), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_1_n38), .QN(aes_state_regs_1_n62) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U119 ( .A(
        aes_state_regs_1_mix_columns_1_n206), .B(
        aes_state_regs_1_mix_columns_1_n205), .ZN(
        aes_state_regs_1_mix_columns_1_n215) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U118 ( .A(
        aes_state_regs_1_mix_columns_1_n191), .B(
        aes_state_regs_1_mix_columns_1_n233), .ZN(
        aes_state_regs_1_MixColumnsS3xD[0]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U117 ( .A1(
        aes_state_regs_1_S20xDP_0_), .A2(aes_state_regs_1_mix_columns_1_n232), 
        .B1(aes_state_regs_1_mix_columns_1_n231), .B2(
        aes_state_regs_1_mix_columns_1_n230), .ZN(
        aes_state_regs_1_mix_columns_1_n191) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U116 ( .A(
        aes_state_regs_1_mix_columns_1_n189), .B(
        aes_state_regs_1_mix_columns_1_n190), .ZN(
        aes_state_regs_1_MixColumnsS1xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U115 ( .A(aes_state_regs_1_S20xDP_1_), .B(aes_state_regs_1_S10xDP_1_), .ZN(aes_state_regs_1_mix_columns_1_n190) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U114 ( .A(
        aes_state_regs_1_mix_columns_1_n212), .B(aes_state_regs_1_S20xDP_2_), 
        .Z(aes_state_regs_1_mix_columns_1_n189) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U113 ( .A(
        aes_state_regs_1_mix_columns_1_n188), .B(
        aes_state_regs_1_mix_columns_1_n215), .ZN(
        aes_state_regs_1_MixColumnsS1xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U112 ( .A(aes_state_regs_1_S20xDP_3_), .B(aes_state_regs_1_mix_columns_1_n203), .ZN(
        aes_state_regs_1_mix_columns_1_n188) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U111 ( .A(
        aes_state_regs_1_mix_columns_1_n186), .B(
        aes_state_regs_1_mix_columns_1_n187), .ZN(
        aes_state_regs_1_MixColumnsS1xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U110 ( .A(aes_state_regs_1_S20xDP_5_), .B(aes_state_regs_1_S10xDP_5_), .ZN(aes_state_regs_1_mix_columns_1_n187) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U109 ( .A(aes_state_regs_1_S00xDP[6]), 
        .B(aes_state_regs_1_mix_columns_1_n229), .Z(
        aes_state_regs_1_mix_columns_1_n186) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U108 ( .A(
        aes_state_regs_1_mix_columns_1_n184), .B(
        aes_state_regs_1_mix_columns_1_n185), .ZN(
        aes_state_regs_1_MixColumnsS3xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U107 ( .A(aes_state_regs_1_S00xDP[2]), .B(aes_state_regs_1_S00xDP[1]), .ZN(aes_state_regs_1_mix_columns_1_n185) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U106 ( .A(
        aes_state_regs_1_mix_columns_1_n236), .B(aes_state_regs_1_S30xDP_1_), 
        .Z(aes_state_regs_1_mix_columns_1_n184) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U105 ( .A(
        aes_state_regs_1_mix_columns_1_n183), .B(
        aes_state_regs_1_mix_columns_1_n217), .ZN(
        aes_state_regs_1_MixColumnsS1xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U104 ( .A(
        aes_state_regs_1_mix_columns_1_n207), .B(aes_state_regs_1_S00xDP[4]), 
        .ZN(aes_state_regs_1_mix_columns_1_n183) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U103 ( .A(
        aes_state_regs_1_mix_columns_1_n182), .B(
        aes_state_regs_1_mix_columns_1_n233), .ZN(
        aes_state_regs_1_MixColumnsS2xD[0]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U102 ( .A(aes_state_regs_1_S20xDP_7_), .B(aes_state_regs_1_mix_columns_1_n210), .ZN(
        aes_state_regs_1_mix_columns_1_n182) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U101 ( .A(
        aes_state_regs_1_mix_columns_1_n180), .B(
        aes_state_regs_1_mix_columns_1_n181), .ZN(
        aes_state_regs_1_MixColumnsS1xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U100 ( .A(aes_state_regs_1_S20xDP_4_), .B(aes_state_regs_1_S10xDP_4_), .ZN(aes_state_regs_1_mix_columns_1_n181) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U99 ( .A(aes_state_regs_1_S00xDP[5]), 
        .B(aes_state_regs_1_mix_columns_1_n225), .Z(
        aes_state_regs_1_mix_columns_1_n180) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U98 ( .A(
        aes_state_regs_1_mix_columns_1_n179), .B(
        aes_state_regs_1_mix_columns_1_n244), .ZN(
        aes_state_regs_1_MixColumnsS1xD[0]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U97 ( .A(
        aes_state_regs_1_mix_columns_1_n201), .B(aes_state_regs_1_S00xDP[0]), 
        .ZN(aes_state_regs_1_mix_columns_1_n179) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U96 ( .A(
        aes_state_regs_1_mix_columns_1_n178), .B(
        aes_state_regs_1_mix_columns_1_n177), .ZN(
        aes_state_regs_1_MixColumnsS3xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U95 ( .A(aes_state_regs_1_S30xDP_5_), 
        .B(aes_state_regs_1_S00xDP[5]), .ZN(
        aes_state_regs_1_mix_columns_1_n178) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U94 ( .A1(
        aes_state_regs_1_mix_columns_1_n243), .A2(aes_state_regs_1_S20xDP_6_), 
        .B1(aes_state_regs_1_mix_columns_1_n242), .B2(
        aes_state_regs_1_mix_columns_1_n176), .ZN(
        aes_state_regs_1_mix_columns_1_n177) );
  INV_X1 aes_state_regs_1_mix_columns_1_U93 ( .A(
        aes_state_regs_1_mix_columns_1_n243), .ZN(
        aes_state_regs_1_mix_columns_1_n176) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U92 ( .A1(aes_state_regs_1_S30xDP_2_), .A2(aes_state_regs_1_S30xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n219), 
        .B2(aes_state_regs_1_mix_columns_1_n175), .ZN(
        aes_state_regs_1_mix_columns_1_n238) );
  INV_X1 aes_state_regs_1_mix_columns_1_U91 ( .A(aes_state_regs_1_S30xDP_2_), 
        .ZN(aes_state_regs_1_mix_columns_1_n175) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U90 ( .A(
        aes_state_regs_1_mix_columns_1_n174), .B(
        aes_state_regs_1_mix_columns_1_n235), .ZN(
        aes_state_regs_1_MixColumnsS3xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U89 ( .A(
        aes_state_regs_1_mix_columns_1_n234), .B(aes_state_regs_1_S20xDP_1_), 
        .ZN(aes_state_regs_1_mix_columns_1_n174) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U88 ( .A(
        aes_state_regs_1_mix_columns_1_n173), .B(
        aes_state_regs_1_mix_columns_1_n209), .ZN(
        aes_state_regs_1_MixColumnsS1xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U87 ( .A(
        aes_state_regs_1_mix_columns_1_n202), .B(aes_state_regs_1_S00xDP[1]), 
        .ZN(aes_state_regs_1_mix_columns_1_n173) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U86 ( .A(
        aes_state_regs_1_mix_columns_1_n172), .B(
        aes_state_regs_1_mix_columns_1_n223), .ZN(
        aes_state_regs_1_mix_columns_1_n207) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U85 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_3_), .ZN(
        aes_state_regs_1_mix_columns_1_n172) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U84 ( .A(
        aes_state_regs_1_mix_columns_1_n171), .B(
        aes_state_regs_1_mix_columns_1_n238), .ZN(
        aes_state_regs_1_MixColumnsS3xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U83 ( .A(
        aes_state_regs_1_mix_columns_1_n237), .B(aes_state_regs_1_S00xDP[3]), 
        .ZN(aes_state_regs_1_mix_columns_1_n171) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U82 ( .A(
        aes_state_regs_1_mix_columns_1_n170), .B(
        aes_state_regs_1_mix_columns_1_n235), .ZN(
        aes_state_regs_1_MixColumnsS2xD[1]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U81 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_mix_columns_1_n209), .ZN(
        aes_state_regs_1_mix_columns_1_n170) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U80 ( .A(
        aes_state_regs_1_mix_columns_1_n168), .B(
        aes_state_regs_1_mix_columns_1_n169), .ZN(
        aes_state_regs_1_mix_columns_1_n237) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U79 ( .A(aes_state_regs_1_S20xDP_3_), 
        .B(aes_state_regs_1_S00xDP[7]), .ZN(
        aes_state_regs_1_mix_columns_1_n169) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U78 ( .A(aes_state_regs_1_S00xDP[2]), 
        .B(aes_state_regs_1_S10xDP_3_), .Z(aes_state_regs_1_mix_columns_1_n168) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U77 ( .A(
        aes_state_regs_1_mix_columns_1_n167), .B(
        aes_state_regs_1_mix_columns_1_n166), .ZN(
        aes_state_regs_1_MixColumnsS3xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U76 ( .A(
        aes_state_regs_1_mix_columns_1_n244), .B(aes_state_regs_1_S30xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n167) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U75 ( .A1(aes_state_regs_1_S00xDP[6]), .A2(aes_state_regs_1_S00xDP[7]), .B1(aes_state_regs_1_mix_columns_1_n245), 
        .B2(aes_state_regs_1_mix_columns_1_n165), .ZN(
        aes_state_regs_1_mix_columns_1_n166) );
  INV_X1 aes_state_regs_1_mix_columns_1_U74 ( .A(aes_state_regs_1_S00xDP[6]), 
        .ZN(aes_state_regs_1_mix_columns_1_n165) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U73 ( .A(
        aes_state_regs_1_mix_columns_1_n164), .B(
        aes_state_regs_1_mix_columns_1_n240), .ZN(
        aes_state_regs_1_MixColumnsS3xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U72 ( .A(
        aes_state_regs_1_mix_columns_1_n239), .B(aes_state_regs_1_S20xDP_4_), 
        .ZN(aes_state_regs_1_mix_columns_1_n164) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U71 ( .A1(aes_state_regs_1_S20xDP_3_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n208), 
        .B2(aes_state_regs_1_mix_columns_1_n163), .ZN(
        aes_state_regs_1_mix_columns_1_n217) );
  INV_X1 aes_state_regs_1_mix_columns_1_U70 ( .A(aes_state_regs_1_S20xDP_3_), 
        .ZN(aes_state_regs_1_mix_columns_1_n163) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U69 ( .A(
        aes_state_regs_1_mix_columns_1_n161), .B(
        aes_state_regs_1_mix_columns_1_n162), .ZN(
        aes_state_regs_1_MixColumnsS3xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U68 ( .A(
        aes_state_regs_1_mix_columns_1_n241), .B(aes_state_regs_1_S20xDP_5_), 
        .ZN(aes_state_regs_1_mix_columns_1_n162) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U67 ( .A(aes_state_regs_1_S00xDP[4]), 
        .B(aes_state_regs_1_S30xDP_4_), .Z(aes_state_regs_1_mix_columns_1_n161) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U66 ( .A(
        aes_state_regs_1_mix_columns_1_n159), .B(
        aes_state_regs_1_mix_columns_1_n160), .ZN(
        aes_state_regs_1_MixColumnsS1xD[7]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U65 ( .A1(aes_state_regs_1_S20xDP_6_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n208), 
        .B2(aes_state_regs_1_mix_columns_1_n242), .ZN(
        aes_state_regs_1_mix_columns_1_n160) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U64 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_mix_columns_1_n231), .ZN(
        aes_state_regs_1_mix_columns_1_n159) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U63 ( .A(aes_state_regs_1_S10xDP_2_), 
        .B(aes_state_regs_1_mix_columns_1_n212), .Z(
        aes_state_regs_1_mix_columns_1_n213) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U62 ( .A(
        aes_state_regs_1_mix_columns_1_n214), .B(
        aes_state_regs_1_mix_columns_1_n213), .ZN(
        aes_state_regs_1_MixColumnsS2xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U61 ( .A(aes_state_regs_1_S10xDP_3_), 
        .B(aes_state_regs_1_mix_columns_1_n215), .ZN(
        aes_state_regs_1_mix_columns_1_n216) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U60 ( .A(
        aes_state_regs_1_mix_columns_1_n216), .B(
        aes_state_regs_1_mix_columns_1_n238), .ZN(
        aes_state_regs_1_MixColumnsS2xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U59 ( .A(aes_state_regs_1_S30xDP_4_), 
        .B(aes_state_regs_1_mix_columns_1_n217), .ZN(
        aes_state_regs_1_mix_columns_1_n222) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U58 ( .A(
        aes_state_regs_1_mix_columns_1_n222), .B(
        aes_state_regs_1_mix_columns_1_n240), .ZN(
        aes_state_regs_1_MixColumnsS2xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U57 ( .A(
        aes_state_regs_1_mix_columns_1_n223), .B(aes_state_regs_1_S30xDP_5_), 
        .ZN(aes_state_regs_1_mix_columns_1_n224) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U56 ( .A(
        aes_state_regs_1_mix_columns_1_n224), .B(
        aes_state_regs_1_mix_columns_1_n241), .ZN(
        aes_state_regs_1_MixColumnsS2xD[5]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U55 ( .A(
        aes_state_regs_1_mix_columns_1_n225), .B(aes_state_regs_1_S30xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n226) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U54 ( .A(
        aes_state_regs_1_mix_columns_1_n226), .B(
        aes_state_regs_1_mix_columns_1_n243), .ZN(
        aes_state_regs_1_MixColumnsS2xD[6]) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U53 ( .A1(aes_state_regs_1_S10xDP_7_), .A2(aes_state_regs_1_mix_columns_1_n232), .B1(
        aes_state_regs_1_mix_columns_1_n231), .B2(
        aes_state_regs_1_mix_columns_1_n227), .ZN(
        aes_state_regs_1_mix_columns_1_n228) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U52 ( .A(
        aes_state_regs_1_mix_columns_1_n229), .B(
        aes_state_regs_1_mix_columns_1_n228), .ZN(
        aes_state_regs_1_MixColumnsS2xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U51 ( .A(
        aes_state_regs_1_mix_columns_1_n244), .B(
        aes_state_regs_1_mix_columns_1_n243), .ZN(
        aes_state_regs_1_mix_columns_1_n200) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U50 ( .A(
        aes_state_regs_1_mix_columns_1_n200), .B(aes_state_regs_1_S30xDP_7_), 
        .ZN(aes_state_regs_1_MixColumnsS0xD[7]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U49 ( .A(aes_state_regs_1_S10xDP_4_), 
        .B(aes_state_regs_1_mix_columns_1_n239), .ZN(
        aes_state_regs_1_mix_columns_1_n197) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U48 ( .A(
        aes_state_regs_1_mix_columns_1_n197), .B(
        aes_state_regs_1_mix_columns_1_n207), .ZN(
        aes_state_regs_1_MixColumnsS0xD[4]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U47 ( .A(aes_state_regs_1_S30xDP_3_), 
        .B(aes_state_regs_1_mix_columns_1_n237), .ZN(
        aes_state_regs_1_mix_columns_1_n196) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U46 ( .A(
        aes_state_regs_1_mix_columns_1_n196), .B(
        aes_state_regs_1_mix_columns_1_n203), .ZN(
        aes_state_regs_1_MixColumnsS0xD[3]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U45 ( .A(aes_state_regs_1_S30xDP_2_), 
        .B(aes_state_regs_1_mix_columns_1_n236), .ZN(
        aes_state_regs_1_mix_columns_1_n195) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U44 ( .A(
        aes_state_regs_1_mix_columns_1_n195), .B(
        aes_state_regs_1_mix_columns_1_n211), .ZN(
        aes_state_regs_1_MixColumnsS0xD[2]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U43 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_mix_columns_1_n193), .ZN(
        aes_state_regs_1_mix_columns_1_n192) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U42 ( .A(
        aes_state_regs_1_mix_columns_1_n192), .B(
        aes_state_regs_1_mix_columns_1_n201), .ZN(
        aes_state_regs_1_MixColumnsS0xD[0]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U41 ( .A(aes_state_regs_1_S10xDP_0_), 
        .B(aes_state_regs_1_S00xDP[0]), .Z(aes_state_regs_1_mix_columns_1_n233) );
  INV_X1 aes_state_regs_1_mix_columns_1_U40 ( .A(
        aes_state_regs_1_mix_columns_1_n231), .ZN(
        aes_state_regs_1_mix_columns_1_n232) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U39 ( .A1(aes_state_regs_1_S00xDP[7]), .A2(aes_state_regs_1_S30xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n219), 
        .B2(aes_state_regs_1_mix_columns_1_n245), .ZN(
        aes_state_regs_1_mix_columns_1_n231) );
  INV_X1 aes_state_regs_1_mix_columns_1_U38 ( .A(aes_state_regs_1_S20xDP_0_), 
        .ZN(aes_state_regs_1_mix_columns_1_n230) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U37 ( .A(aes_state_regs_1_S30xDP_0_), 
        .B(aes_state_regs_1_mix_columns_1_n219), .ZN(
        aes_state_regs_1_mix_columns_1_n210) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U36 ( .A(aes_state_regs_1_S30xDP_0_), 
        .B(aes_state_regs_1_S20xDP_0_), .Z(aes_state_regs_1_mix_columns_1_n201) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U35 ( .A1(aes_state_regs_1_S10xDP_7_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n208), 
        .B2(aes_state_regs_1_mix_columns_1_n227), .ZN(
        aes_state_regs_1_mix_columns_1_n244) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U34 ( .A(
        aes_state_regs_1_mix_columns_1_n211), .B(
        aes_state_regs_1_mix_columns_1_n210), .Z(
        aes_state_regs_1_mix_columns_1_n235) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U33 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_S00xDP[0]), .Z(aes_state_regs_1_mix_columns_1_n234) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U32 ( .A(aes_state_regs_1_S10xDP_2_), 
        .B(aes_state_regs_1_S20xDP_2_), .Z(aes_state_regs_1_mix_columns_1_n236) );
  INV_X1 aes_state_regs_1_mix_columns_1_U31 ( .A(aes_state_regs_1_S30xDP_3_), 
        .ZN(aes_state_regs_1_mix_columns_1_n218) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U30 ( .A1(aes_state_regs_1_S30xDP_3_), .A2(aes_state_regs_1_mix_columns_1_n219), .B1(aes_state_regs_1_S30xDP_7_), 
        .B2(aes_state_regs_1_mix_columns_1_n218), .ZN(
        aes_state_regs_1_mix_columns_1_n220) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U29 ( .A(
        aes_state_regs_1_mix_columns_1_n221), .B(
        aes_state_regs_1_mix_columns_1_n220), .ZN(
        aes_state_regs_1_mix_columns_1_n240) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U28 ( .A(aes_state_regs_1_S00xDP[7]), 
        .B(aes_state_regs_1_S00xDP[3]), .Z(aes_state_regs_1_mix_columns_1_n239) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U27 ( .A(aes_state_regs_1_S10xDP_5_), 
        .B(aes_state_regs_1_S00xDP[5]), .Z(aes_state_regs_1_mix_columns_1_n241) );
  INV_X1 aes_state_regs_1_mix_columns_1_U26 ( .A(aes_state_regs_1_S20xDP_6_), 
        .ZN(aes_state_regs_1_mix_columns_1_n242) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U25 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_S00xDP[6]), .Z(aes_state_regs_1_mix_columns_1_n243) );
  INV_X1 aes_state_regs_1_mix_columns_1_U24 ( .A(aes_state_regs_1_S00xDP[7]), 
        .ZN(aes_state_regs_1_mix_columns_1_n245) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U23 ( .A1(aes_state_regs_1_S20xDP_0_), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n208), 
        .B2(aes_state_regs_1_mix_columns_1_n230), .ZN(
        aes_state_regs_1_mix_columns_1_n209) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U22 ( .A(aes_state_regs_1_S30xDP_2_), 
        .B(aes_state_regs_1_S00xDP[2]), .Z(aes_state_regs_1_mix_columns_1_n212) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U21 ( .A(aes_state_regs_1_S30xDP_1_), 
        .B(aes_state_regs_1_S20xDP_1_), .ZN(
        aes_state_regs_1_mix_columns_1_n214) );
  INV_X1 aes_state_regs_1_mix_columns_1_U20 ( .A(aes_state_regs_1_S00xDP[3]), 
        .ZN(aes_state_regs_1_mix_columns_1_n204) );
  AOI22_X1 aes_state_regs_1_mix_columns_1_U19 ( .A1(aes_state_regs_1_S00xDP[3]), .A2(aes_state_regs_1_S20xDP_7_), .B1(aes_state_regs_1_mix_columns_1_n208), 
        .B2(aes_state_regs_1_mix_columns_1_n204), .ZN(
        aes_state_regs_1_mix_columns_1_n205) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U18 ( .A(aes_state_regs_1_S20xDP_2_), 
        .B(aes_state_regs_1_S30xDP_3_), .ZN(
        aes_state_regs_1_mix_columns_1_n206) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U17 ( .A(aes_state_regs_1_S30xDP_4_), 
        .B(aes_state_regs_1_S20xDP_4_), .Z(aes_state_regs_1_mix_columns_1_n223) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U16 ( .A(aes_state_regs_1_S30xDP_5_), 
        .B(aes_state_regs_1_S20xDP_5_), .Z(aes_state_regs_1_mix_columns_1_n225) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U15 ( .A(aes_state_regs_1_S30xDP_6_), 
        .B(aes_state_regs_1_S20xDP_6_), .Z(aes_state_regs_1_mix_columns_1_n229) );
  INV_X1 aes_state_regs_1_mix_columns_1_U14 ( .A(aes_state_regs_1_S10xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n227) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U13 ( .A(
        aes_state_regs_1_mix_columns_1_n193), .B(
        aes_state_regs_1_mix_columns_1_n214), .ZN(
        aes_state_regs_1_mix_columns_1_n202) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U12 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_2_), .Z(aes_state_regs_1_mix_columns_1_n203) );
  INV_X1 aes_state_regs_1_mix_columns_1_U11 ( .A(aes_state_regs_1_S20xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n208) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U10 ( .A(aes_state_regs_1_S10xDP_6_), 
        .B(aes_state_regs_1_mix_columns_1_n241), .ZN(
        aes_state_regs_1_mix_columns_1_n199) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U9 ( .A(
        aes_state_regs_1_mix_columns_1_n199), .B(
        aes_state_regs_1_mix_columns_1_n229), .ZN(
        aes_state_regs_1_MixColumnsS0xD[6]) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U8 ( .A(aes_state_regs_1_S10xDP_5_), 
        .B(aes_state_regs_1_mix_columns_1_n221), .ZN(
        aes_state_regs_1_mix_columns_1_n198) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U7 ( .A(
        aes_state_regs_1_mix_columns_1_n198), .B(
        aes_state_regs_1_mix_columns_1_n225), .ZN(
        aes_state_regs_1_MixColumnsS0xD[5]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U6 ( .A(aes_state_regs_1_S10xDP_1_), 
        .B(aes_state_regs_1_S00xDP[1]), .Z(aes_state_regs_1_mix_columns_1_n211) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U5 ( .A(aes_state_regs_1_S10xDP_1_), 
        .B(aes_state_regs_1_mix_columns_1_n234), .ZN(
        aes_state_regs_1_mix_columns_1_n194) );
  XNOR2_X1 aes_state_regs_1_mix_columns_1_U4 ( .A(
        aes_state_regs_1_mix_columns_1_n194), .B(
        aes_state_regs_1_mix_columns_1_n202), .ZN(
        aes_state_regs_1_MixColumnsS0xD[1]) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U3 ( .A(aes_state_regs_1_S10xDP_7_), 
        .B(aes_state_regs_1_S10xDP_0_), .Z(aes_state_regs_1_mix_columns_1_n193) );
  INV_X1 aes_state_regs_1_mix_columns_1_U2 ( .A(aes_state_regs_1_S30xDP_7_), 
        .ZN(aes_state_regs_1_mix_columns_1_n219) );
  XOR2_X1 aes_state_regs_1_mix_columns_1_U1 ( .A(aes_state_regs_1_S10xDP_4_), 
        .B(aes_state_regs_1_S00xDP[4]), .Z(aes_state_regs_1_mix_columns_1_n221) );
  BUF_X1 aes_key_regs_0_U3 ( .A(n114), .Z(aes_key_regs_0_n4) );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_0_ ( .D(aes_key_regs_0_K00xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_0_ ( .D(aes_key_regs_0_K10xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_0_ ( .D(aes_key_regs_0_K20xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_0_ ( .D(aes_key_regs_0_K01xDP_0_), .SI(
        KeyOutxD[0]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_0_ ( .D(aes_key_regs_0_K01xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_0_ ( .D(aes_key_regs_0_K11xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_0_ ( .D(aes_key_regs_0_K21xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_0_ ( .D(aes_key_regs_0_K02xDP_0_), .SI(
        aes_key_regs_0_K01xDP_0_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_0_ ( .D(aes_key_regs_0_K02xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_0_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_0_ ( .D(aes_key_regs_0_K12xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_0_ ( .D(aes_key_regs_0_K22xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_0_ ( .D(K03xD[0]), .SI(
        aes_key_regs_0_K02xDP_0_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_1_ ( .D(aes_key_regs_0_K00xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_1_ ( .D(aes_key_regs_0_K10xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_1_ ( .D(aes_key_regs_0_K20xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_1_ ( .D(aes_key_regs_0_K01xDP_1_), .SI(
        KeyOutxD[1]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_1_ ( .D(aes_key_regs_0_K01xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_1_ ( .D(aes_key_regs_0_K11xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_1_ ( .D(aes_key_regs_0_K21xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_1_ ( .D(aes_key_regs_0_K02xDP_1_), .SI(
        aes_key_regs_0_K01xDP_1_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_1_ ( .D(aes_key_regs_0_K02xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_1_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_1_ ( .D(aes_key_regs_0_K12xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_1_ ( .D(aes_key_regs_0_K22xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_1_ ( .D(K03xD[1]), .SI(
        aes_key_regs_0_K02xDP_1_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_2_ ( .D(aes_key_regs_0_K00xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_2_ ( .D(aes_key_regs_0_K10xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_2_ ( .D(aes_key_regs_0_K20xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_2_ ( .D(aes_key_regs_0_K01xDP_2_), .SI(
        KeyOutxD[2]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_2_ ( .D(aes_key_regs_0_K01xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_2_ ( .D(aes_key_regs_0_K11xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_2_ ( .D(aes_key_regs_0_K21xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_2_ ( .D(aes_key_regs_0_K02xDP_2_), .SI(
        aes_key_regs_0_K01xDP_2_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K21xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_2_ ( .D(aes_key_regs_0_K02xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_2_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_2_ ( .D(aes_key_regs_0_K12xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_2_ ( .D(aes_key_regs_0_K22xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_2_ ( .D(K03xD[2]), .SI(
        aes_key_regs_0_K02xDP_2_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_3_ ( .D(aes_key_regs_0_K00xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_3_ ( .D(aes_key_regs_0_K10xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_3_ ( .D(aes_key_regs_0_K20xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_3_ ( .D(aes_key_regs_0_K01xDP_3_), .SI(
        KeyOutxD[3]), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K20xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_3_ ( .D(aes_key_regs_0_K01xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_3_ ( .D(aes_key_regs_0_K11xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_3_ ( .D(aes_key_regs_0_K21xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_3_ ( .D(aes_key_regs_0_K02xDP_3_), .SI(
        aes_key_regs_0_K01xDP_3_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_3_ ( .D(aes_key_regs_0_K02xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_3_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_3_ ( .D(aes_key_regs_0_K12xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_3_ ( .D(aes_key_regs_0_K22xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_3_ ( .D(K03xD[3]), .SI(
        aes_key_regs_0_K02xDP_3_), .SE(aes_key_regs_0_n4), .CK(ClkKeyRegxC), 
        .RN(RstxBI), .Q(aes_key_regs_0_K22xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_4_ ( .D(aes_key_regs_0_K00xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_4_ ( .D(aes_key_regs_0_K10xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_4_ ( .D(aes_key_regs_0_K20xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_4_ ( .D(aes_key_regs_0_K01xDP_4_), .SI(
        KeyOutxD[4]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_4_ ( .D(aes_key_regs_0_K01xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_4_ ( .D(aes_key_regs_0_K11xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_4_ ( .D(aes_key_regs_0_K21xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_4_ ( .D(aes_key_regs_0_K02xDP_4_), .SI(
        aes_key_regs_0_K01xDP_4_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_4_ ( .D(aes_key_regs_0_K02xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_4_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_4_ ( .D(aes_key_regs_0_K12xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_4_ ( .D(aes_key_regs_0_K22xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_4_ ( .D(K03xD[4]), .SI(
        aes_key_regs_0_K02xDP_4_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_5_ ( .D(aes_key_regs_0_K00xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_5_ ( .D(aes_key_regs_0_K10xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_5_ ( .D(aes_key_regs_0_K20xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_5_ ( .D(aes_key_regs_0_K01xDP_5_), .SI(
        KeyOutxD[5]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_5_ ( .D(aes_key_regs_0_K01xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_5_ ( .D(aes_key_regs_0_K11xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_5_ ( .D(aes_key_regs_0_K21xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_5_ ( .D(aes_key_regs_0_K02xDP_5_), .SI(
        aes_key_regs_0_K01xDP_5_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_5_ ( .D(aes_key_regs_0_K02xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_5_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_5_ ( .D(aes_key_regs_0_K12xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_5_ ( .D(aes_key_regs_0_K22xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_5_ ( .D(K03xD[5]), .SI(
        aes_key_regs_0_K02xDP_5_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_6_ ( .D(aes_key_regs_0_K00xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_6_ ( .D(aes_key_regs_0_K10xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_6_ ( .D(aes_key_regs_0_K20xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_6_ ( .D(aes_key_regs_0_K01xDP_6_), .SI(
        KeyOutxD[6]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_6_ ( .D(aes_key_regs_0_K01xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_6_ ( .D(aes_key_regs_0_K11xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_6_ ( .D(aes_key_regs_0_K21xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_6_ ( .D(aes_key_regs_0_K02xDP_6_), .SI(
        aes_key_regs_0_K01xDP_6_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_6_ ( .D(aes_key_regs_0_K02xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_6_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_6_ ( .D(aes_key_regs_0_K12xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_6_ ( .D(aes_key_regs_0_K22xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_6_ ( .D(K03xD[6]), .SI(
        aes_key_regs_0_K02xDP_6_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K00xDP_reg_7_ ( .D(aes_key_regs_0_K00xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyOutxD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K10xDP_reg_7_ ( .D(aes_key_regs_0_K10xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K00xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K20xDP_reg_7_ ( .D(aes_key_regs_0_K20xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K10xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K30xDP_reg_7_ ( .D(aes_key_regs_0_K01xDP_7_), .SI(
        KeyOutxD[7]), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K20xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K01xDP_reg_7_ ( .D(aes_key_regs_0_K01xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_0_K11xDP_reg_7_ ( .D(aes_key_regs_0_K11xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K01xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K21xDP_reg_7_ ( .D(aes_key_regs_0_K21xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K11xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K31xDP_reg_7_ ( .D(aes_key_regs_0_K02xDP_7_), .SI(
        aes_key_regs_0_K01xDP_7_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K21xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K02xDP_reg_7_ ( .D(aes_key_regs_0_K02xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDP_7_), .QN() );
  DFFR_X1 aes_key_regs_0_K12xDP_reg_7_ ( .D(aes_key_regs_0_K12xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K02xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K22xDP_reg_7_ ( .D(aes_key_regs_0_K22xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K12xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K32xDP_reg_7_ ( .D(K03xD[7]), .SI(
        aes_key_regs_0_K02xDP_7_), .SE(n114), .CK(ClkKeyRegxC), .RN(RstxBI), 
        .Q(aes_key_regs_0_K22xDN[7]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_0_ ( .D(KeyInxD[0]), .SI(K03xD[0]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_0_ ( .D(KeyToSboxOutxD[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_0_ ( .D(aes_key_regs_0_K13xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[0]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_0_ ( .D(aes_key_regs_0_K23xDN[0]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[0]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_1_ ( .D(KeyInxD[1]), .SI(K03xD[1]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_1_ ( .D(KeyToSboxOutxD[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_1_ ( .D(aes_key_regs_0_K13xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[1]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_1_ ( .D(aes_key_regs_0_K23xDN[1]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[1]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_2_ ( .D(KeyInxD[2]), .SI(K03xD[2]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_2_ ( .D(KeyToSboxOutxD[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_2_ ( .D(aes_key_regs_0_K13xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[2]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_2_ ( .D(aes_key_regs_0_K23xDN[2]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[2]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_3_ ( .D(KeyInxD[3]), .SI(K03xD[3]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_3_ ( .D(KeyToSboxOutxD[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_3_ ( .D(aes_key_regs_0_K13xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[3]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_3_ ( .D(aes_key_regs_0_K23xDN[3]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[3]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_4_ ( .D(KeyInxD[4]), .SI(K03xD[4]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_4_ ( .D(KeyToSboxOutxD[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_4_ ( .D(aes_key_regs_0_K13xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[4]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_4_ ( .D(aes_key_regs_0_K23xDN[4]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[4]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_5_ ( .D(KeyInxD[5]), .SI(K03xD[5]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_5_ ( .D(KeyToSboxOutxD[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_5_ ( .D(aes_key_regs_0_K13xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[5]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_5_ ( .D(aes_key_regs_0_K23xDN[5]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[5]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_6_ ( .D(KeyInxD[6]), .SI(K03xD[6]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_6_ ( .D(KeyToSboxOutxD[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_6_ ( .D(aes_key_regs_0_K13xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[6]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_6_ ( .D(aes_key_regs_0_K23xDN[6]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[6]), .QN() );
  SDFFR_X1 aes_key_regs_0_K33xDP_reg_7_ ( .D(KeyInxD[7]), .SI(K03xD[7]), .SE(
        aes_key_regs_0_n4), .CK(ClkKeyRegxC), .RN(RstxBI), .Q(
        aes_key_regs_0_K23xDN[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K03xDP_reg_7_ ( .D(KeyToSboxOutxD[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(K03xD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K13xDP_reg_7_ ( .D(aes_key_regs_0_K13xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(KeyToSboxOutxD[7]), .QN() );
  DFFR_X1 aes_key_regs_0_K23xDP_reg_7_ ( .D(aes_key_regs_0_K23xDN[7]), .CK(
        ClkKeyRegxC), .RN(RstxBI), .Q(aes_key_regs_0_K13xDN[7]), .QN() );
  AOI22_X1 aes_state_regs_0_U56 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n151), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[3]), .ZN(aes_state_regs_0_n190) );
  AOI22_X1 aes_state_regs_0_U55 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n146), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[2]), .ZN(aes_state_regs_0_n189) );
  AOI22_X1 aes_state_regs_0_U54 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n141), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[1]), .ZN(aes_state_regs_0_n188) );
  AOI22_X1 aes_state_regs_0_U53 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n136), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[0]), .ZN(aes_state_regs_0_n187) );
  OAI222_X1 aes_state_regs_0_U52 ( .A1(aes_state_regs_0_n186), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n44), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n127), .ZN(aes_state_regs_0_S10xDN[7]) );
  INV_X1 aes_state_regs_0_U51 ( .A(aes_state_regs_0_MixColumnsS2xD[7]), .ZN(
        aes_state_regs_0_n186) );
  OAI222_X1 aes_state_regs_0_U50 ( .A1(aes_state_regs_0_n185), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n45), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n126), .ZN(aes_state_regs_0_S10xDN[6]) );
  INV_X1 aes_state_regs_0_U49 ( .A(aes_state_regs_0_MixColumnsS2xD[6]), .ZN(
        aes_state_regs_0_n185) );
  OAI222_X1 aes_state_regs_0_U48 ( .A1(aes_state_regs_0_n184), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n46), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n125), .ZN(aes_state_regs_0_S10xDN[5]) );
  INV_X1 aes_state_regs_0_U47 ( .A(aes_state_regs_0_MixColumnsS2xD[5]), .ZN(
        aes_state_regs_0_n184) );
  OAI222_X1 aes_state_regs_0_U46 ( .A1(aes_state_regs_0_n183), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n47), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n124), .ZN(aes_state_regs_0_S10xDN[4]) );
  INV_X1 aes_state_regs_0_U45 ( .A(aes_state_regs_0_MixColumnsS2xD[4]), .ZN(
        aes_state_regs_0_n183) );
  OAI222_X1 aes_state_regs_0_U44 ( .A1(aes_state_regs_0_n182), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n48), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n123), .ZN(aes_state_regs_0_S10xDN[3]) );
  INV_X1 aes_state_regs_0_U43 ( .A(aes_state_regs_0_MixColumnsS2xD[3]), .ZN(
        aes_state_regs_0_n182) );
  OAI222_X1 aes_state_regs_0_U42 ( .A1(aes_state_regs_0_n181), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n49), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n122), .ZN(aes_state_regs_0_S10xDN[2]) );
  INV_X1 aes_state_regs_0_U41 ( .A(aes_state_regs_0_MixColumnsS2xD[2]), .ZN(
        aes_state_regs_0_n181) );
  OAI222_X1 aes_state_regs_0_U40 ( .A1(aes_state_regs_0_n180), .A2(
        aes_state_regs_0_n109), .B1(aes_state_regs_0_n195), .B2(
        aes_state_regs_0_n50), .C1(aes_state_regs_0_n178), .C2(
        aes_state_regs_0_n121), .ZN(aes_state_regs_0_S10xDN[1]) );
  INV_X1 aes_state_regs_0_U39 ( .A(aes_state_regs_0_MixColumnsS2xD[1]), .ZN(
        aes_state_regs_0_n180) );
  AOI22_X1 aes_state_regs_0_U38 ( .A1(aes_state_regs_0_n177), .A2(
        aes_state_regs_0_n138), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS2xD[0]), .ZN(aes_state_regs_0_n179) );
  NAND2_X1 aes_state_regs_0_U37 ( .A1(doMixColumnsxS), .A2(
        aes_state_regs_0_n178), .ZN(aes_state_regs_0_n109) );
  INV_X1 aes_state_regs_0_U36 ( .A(nextRCONxS), .ZN(aes_state_regs_0_n178) );
  INV_X1 aes_state_regs_0_U35 ( .A(aes_state_regs_0_n178), .ZN(
        aes_state_regs_0_n177) );
  INV_X4 aes_state_regs_0_U34 ( .A(aes_state_regs_0_n178), .ZN(
        aes_state_regs_0_n176) );
  OAI21_X1 aes_state_regs_0_U33 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n35), .A(aes_state_regs_0_n175), .ZN(StateOutxD[0])
         );
  NAND2_X1 aes_state_regs_0_U32 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[0]), .ZN(aes_state_regs_0_n175) );
  OAI21_X1 aes_state_regs_0_U31 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n33), .A(aes_state_regs_0_n174), .ZN(StateOutxD[5])
         );
  NAND2_X1 aes_state_regs_0_U30 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[5]), .ZN(aes_state_regs_0_n174) );
  OAI21_X1 aes_state_regs_0_U29 ( .B1(aes_state_regs_0_n43), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n187), .ZN(
        aes_state_regs_0_S20xDN[0]) );
  OAI21_X1 aes_state_regs_0_U28 ( .B1(aes_state_regs_0_n51), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n179), .ZN(
        aes_state_regs_0_S10xDN[0]) );
  OAI21_X1 aes_state_regs_0_U27 ( .B1(aes_state_regs_0_n42), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n188), .ZN(
        aes_state_regs_0_S20xDN[1]) );
  OAI21_X1 aes_state_regs_0_U26 ( .B1(aes_state_regs_0_n41), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n189), .ZN(
        aes_state_regs_0_S20xDN[2]) );
  OAI21_X1 aes_state_regs_0_U25 ( .B1(aes_state_regs_0_n40), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n190), .ZN(
        aes_state_regs_0_S20xDN[3]) );
  AOI22_X1 aes_state_regs_0_U24 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n156), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[4]), .ZN(aes_state_regs_0_n191) );
  OAI21_X1 aes_state_regs_0_U23 ( .B1(aes_state_regs_0_n39), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n191), .ZN(
        aes_state_regs_0_S20xDN[4]) );
  AOI22_X1 aes_state_regs_0_U22 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n161), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[5]), .ZN(aes_state_regs_0_n192) );
  OAI21_X1 aes_state_regs_0_U21 ( .B1(aes_state_regs_0_n38), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n192), .ZN(
        aes_state_regs_0_S20xDN[5]) );
  AOI22_X1 aes_state_regs_0_U20 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n166), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[6]), .ZN(aes_state_regs_0_n193) );
  OAI21_X1 aes_state_regs_0_U19 ( .B1(aes_state_regs_0_n37), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n193), .ZN(
        aes_state_regs_0_S20xDN[6]) );
  AOI22_X1 aes_state_regs_0_U18 ( .A1(aes_state_regs_0_n176), .A2(
        aes_state_regs_0_n171), .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_MixColumnsS3xD[7]), .ZN(aes_state_regs_0_n194) );
  OAI21_X1 aes_state_regs_0_U17 ( .B1(aes_state_regs_0_n36), .B2(
        aes_state_regs_0_n195), .A(aes_state_regs_0_n194), .ZN(
        aes_state_regs_0_S20xDN[7]) );
  NAND2_X1 aes_state_regs_0_U16 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[7]), .ZN(aes_state_regs_0_n196) );
  OAI21_X1 aes_state_regs_0_U15 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n28), .A(aes_state_regs_0_n196), .ZN(StateOutxD[7])
         );
  NAND2_X1 aes_state_regs_0_U14 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[6]), .ZN(aes_state_regs_0_n197) );
  OAI21_X1 aes_state_regs_0_U13 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n34), .A(aes_state_regs_0_n197), .ZN(StateOutxD[6])
         );
  NAND2_X1 aes_state_regs_0_U12 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[4]), .ZN(aes_state_regs_0_n198) );
  OAI21_X1 aes_state_regs_0_U11 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n32), .A(aes_state_regs_0_n198), .ZN(StateOutxD[4])
         );
  NAND2_X1 aes_state_regs_0_U10 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[3]), .ZN(aes_state_regs_0_n199) );
  OAI21_X1 aes_state_regs_0_U9 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n31), .A(aes_state_regs_0_n199), .ZN(StateOutxD[3])
         );
  NAND2_X1 aes_state_regs_0_U8 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[2]), .ZN(aes_state_regs_0_n200) );
  OAI21_X1 aes_state_regs_0_U7 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n30), .A(aes_state_regs_0_n200), .ZN(StateOutxD[2])
         );
  NAND2_X1 aes_state_regs_0_U6 ( .A1(aes_state_regs_0_n202), .A2(
        aes_state_regs_0_MixColumnsS0xD[1]), .ZN(aes_state_regs_0_n201) );
  OAI21_X1 aes_state_regs_0_U5 ( .B1(aes_state_regs_0_n202), .B2(
        aes_state_regs_0_n29), .A(aes_state_regs_0_n201), .ZN(StateOutxD[1])
         );
  OR2_X1 aes_state_regs_0_U4 ( .A1(aes_state_regs_0_n177), .A2(doMixColumnsxS), 
        .ZN(aes_state_regs_0_n195) );
  INV_X2 aes_state_regs_0_U3 ( .A(aes_state_regs_0_n109), .ZN(
        aes_state_regs_0_n202) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_7_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[7]), .SI(aes_state_regs_0_S10xDP_7_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[7]), .QN(aes_state_regs_0_n28) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_6_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[6]), .SI(aes_state_regs_0_S10xDP_6_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[6]), .QN(aes_state_regs_0_n34) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_5_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[5]), .SI(aes_state_regs_0_S10xDP_5_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[5]), .QN(aes_state_regs_0_n33) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_4_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[4]), .SI(aes_state_regs_0_S10xDP_4_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[4]), .QN(aes_state_regs_0_n32) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_3_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[3]), .SI(aes_state_regs_0_S10xDP_3_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[3]), .QN(aes_state_regs_0_n31) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_2_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[2]), .SI(aes_state_regs_0_S10xDP_2_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[2]), .QN(aes_state_regs_0_n30) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_1_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[1]), .SI(aes_state_regs_0_S10xDP_1_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[1]), .QN(aes_state_regs_0_n29) );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_7_ ( .D(aes_state_regs_0_S10xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_7_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_6_ ( .D(aes_state_regs_0_S10xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_6_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_5_ ( .D(aes_state_regs_0_S10xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_5_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_4_ ( .D(aes_state_regs_0_S10xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_4_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_3_ ( .D(aes_state_regs_0_S10xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_3_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_2_ ( .D(aes_state_regs_0_S10xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_2_), .QN() );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_1_ ( .D(aes_state_regs_0_S10xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_7_ ( .D(aes_state_regs_0_S01xDO_7_), 
        .SI(StateInxD[7]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_7_), .QN(aes_state_regs_0_n36) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_7_ ( .D(aes_state_regs_0_n173), .SI(
        aes_state_regs_0_n170), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[7]), .QN(aes_state_regs_0_n127) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_7_ ( .D(aes_state_regs_0_S02xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_7_ ( .D(aes_state_regs_0_n172), .SI(
        aes_state_regs_0_S23xDP_7_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_7_ ( .D(aes_state_regs_0_n170), .SI(
        aes_state_regs_0_n173), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_7_ ( .D(aes_state_regs_0_S02xDP_7_), 
        .SI(aes_state_regs_0_S01xDO_7_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n173), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_7_ ( .D(aes_state_regs_0_S01xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_7_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_7_ ( .D(aes_state_regs_0_S21xDP[7]), 
        .SI(aes_state_regs_0_n172), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[7]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_7_ ( .D(aes_state_regs_0_n171), .SI(
        aes_state_regs_0_S30xDP_7_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n172), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_7_ ( .D(aes_state_regs_0_n169), .SI(
        aes_state_regs_0_S02xDP_7_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n171), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_7_ ( .D(StateInxD[7]), .SI(
        aes_state_regs_0_n169), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n170), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_7_ ( .D(aes_state_regs_0_S03xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n169), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_7_ ( .D(aes_state_regs_0_S23xDP_7_), 
        .SI(aes_state_regs_0_S20xDP_7_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[7]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_7_ ( .D(aes_state_regs_0_S20xDN[7]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_7_), .QN(
        aes_state_regs_0_n44) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_6_ ( .D(aes_state_regs_0_S01xDO_6_), 
        .SI(StateInxD[6]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_6_), .QN(aes_state_regs_0_n37) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_6_ ( .D(aes_state_regs_0_n168), .SI(
        aes_state_regs_0_n165), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[6]), .QN(aes_state_regs_0_n126) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_6_ ( .D(aes_state_regs_0_S02xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_6_ ( .D(aes_state_regs_0_n167), .SI(
        aes_state_regs_0_S23xDP_6_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_6_ ( .D(aes_state_regs_0_n165), .SI(
        aes_state_regs_0_n168), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_6_ ( .D(aes_state_regs_0_S02xDP_6_), 
        .SI(aes_state_regs_0_S01xDO_6_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n168), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_6_ ( .D(aes_state_regs_0_S01xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_6_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_6_ ( .D(aes_state_regs_0_S21xDP[6]), 
        .SI(aes_state_regs_0_n167), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[6]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_6_ ( .D(aes_state_regs_0_n166), .SI(
        aes_state_regs_0_S30xDP_6_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n167), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_6_ ( .D(aes_state_regs_0_n164), .SI(
        aes_state_regs_0_S02xDP_6_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n166), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_6_ ( .D(StateInxD[6]), .SI(
        aes_state_regs_0_n164), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n165), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_6_ ( .D(aes_state_regs_0_S03xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n164), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_6_ ( .D(aes_state_regs_0_S23xDP_6_), 
        .SI(aes_state_regs_0_S20xDP_6_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[6]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_6_ ( .D(aes_state_regs_0_S20xDN[6]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_6_), .QN(
        aes_state_regs_0_n45) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_5_ ( .D(aes_state_regs_0_S01xDO_5_), 
        .SI(StateInxD[5]), .SE(nextRCONxS), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S30xDP_5_), .QN(aes_state_regs_0_n38) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_5_ ( .D(aes_state_regs_0_n163), .SI(
        aes_state_regs_0_n160), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[5]), .QN(aes_state_regs_0_n125) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_5_ ( .D(aes_state_regs_0_S02xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_5_ ( .D(aes_state_regs_0_n162), .SI(
        aes_state_regs_0_S23xDP_5_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_5_ ( .D(aes_state_regs_0_n160), .SI(
        aes_state_regs_0_n163), .SE(nextRCONxS), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S23xDP_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_5_ ( .D(aes_state_regs_0_S02xDP_5_), 
        .SI(aes_state_regs_0_S01xDO_5_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n163), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_5_ ( .D(aes_state_regs_0_S01xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_5_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_5_ ( .D(aes_state_regs_0_S21xDP[5]), 
        .SI(aes_state_regs_0_n162), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[5]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_5_ ( .D(aes_state_regs_0_n161), .SI(
        aes_state_regs_0_S30xDP_5_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n162), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_5_ ( .D(aes_state_regs_0_n159), .SI(
        aes_state_regs_0_S02xDP_5_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n161), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_5_ ( .D(StateInxD[5]), .SI(
        aes_state_regs_0_n159), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n160), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_5_ ( .D(aes_state_regs_0_S03xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n159), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_5_ ( .D(aes_state_regs_0_S23xDP_5_), 
        .SI(aes_state_regs_0_S20xDP_5_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[5]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_5_ ( .D(aes_state_regs_0_S20xDN[5]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_5_), .QN(
        aes_state_regs_0_n46) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_4_ ( .D(aes_state_regs_0_S01xDO_4_), 
        .SI(StateInxD[4]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_4_), .QN(aes_state_regs_0_n39) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_4_ ( .D(aes_state_regs_0_n158), .SI(
        aes_state_regs_0_n155), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[4]), .QN(aes_state_regs_0_n124) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_4_ ( .D(aes_state_regs_0_S02xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_4_ ( .D(aes_state_regs_0_n157), .SI(
        aes_state_regs_0_S23xDP_4_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_4_ ( .D(aes_state_regs_0_n155), .SI(
        aes_state_regs_0_n158), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_4_ ( .D(aes_state_regs_0_S02xDP_4_), 
        .SI(aes_state_regs_0_S01xDO_4_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n158), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_4_ ( .D(aes_state_regs_0_S01xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_4_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_4_ ( .D(aes_state_regs_0_S21xDP[4]), 
        .SI(aes_state_regs_0_n157), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[4]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_4_ ( .D(aes_state_regs_0_n156), .SI(
        aes_state_regs_0_S30xDP_4_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n157), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_4_ ( .D(aes_state_regs_0_n154), .SI(
        aes_state_regs_0_S02xDP_4_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n156), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_4_ ( .D(StateInxD[4]), .SI(
        aes_state_regs_0_n154), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n155), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_4_ ( .D(aes_state_regs_0_S03xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n154), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_4_ ( .D(aes_state_regs_0_S23xDP_4_), 
        .SI(aes_state_regs_0_S20xDP_4_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[4]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_4_ ( .D(aes_state_regs_0_S20xDN[4]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_4_), .QN(
        aes_state_regs_0_n47) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_3_ ( .D(aes_state_regs_0_S01xDO_3_), 
        .SI(StateInxD[3]), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_3_), .QN(aes_state_regs_0_n40) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_3_ ( .D(aes_state_regs_0_n153), .SI(
        aes_state_regs_0_n150), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[3]), .QN(aes_state_regs_0_n123) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_3_ ( .D(aes_state_regs_0_S02xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_3_ ( .D(aes_state_regs_0_n152), .SI(
        aes_state_regs_0_S23xDP_3_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_3_ ( .D(aes_state_regs_0_n150), .SI(
        aes_state_regs_0_n153), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_3_ ( .D(aes_state_regs_0_S02xDP_3_), 
        .SI(aes_state_regs_0_S01xDO_3_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n153), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_3_ ( .D(aes_state_regs_0_S01xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_3_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_3_ ( .D(aes_state_regs_0_S21xDP[3]), 
        .SI(aes_state_regs_0_n152), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[3]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_3_ ( .D(aes_state_regs_0_n151), .SI(
        aes_state_regs_0_S30xDP_3_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n152), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_3_ ( .D(aes_state_regs_0_n149), .SI(
        aes_state_regs_0_S02xDP_3_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n151), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_3_ ( .D(StateInxD[3]), .SI(
        aes_state_regs_0_n149), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n150), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_3_ ( .D(aes_state_regs_0_S03xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n149), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_3_ ( .D(aes_state_regs_0_S23xDP_3_), 
        .SI(aes_state_regs_0_S20xDP_3_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[3]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_3_ ( .D(aes_state_regs_0_S20xDN[3]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_3_), .QN(
        aes_state_regs_0_n48) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_2_ ( .D(aes_state_regs_0_S01xDO_2_), 
        .SI(StateInxD[2]), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_2_), .QN(aes_state_regs_0_n41) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_2_ ( .D(aes_state_regs_0_n148), .SI(
        aes_state_regs_0_n145), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[2]), .QN(aes_state_regs_0_n122) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_2_ ( .D(aes_state_regs_0_S02xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_2_ ( .D(aes_state_regs_0_n147), .SI(
        aes_state_regs_0_S23xDP_2_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_2_ ( .D(aes_state_regs_0_n145), .SI(
        aes_state_regs_0_n148), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_2_ ( .D(aes_state_regs_0_S02xDP_2_), 
        .SI(aes_state_regs_0_S01xDO_2_), .SE(aes_state_regs_0_n177), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n148), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_2_ ( .D(aes_state_regs_0_S01xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_2_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_2_ ( .D(aes_state_regs_0_S21xDP[2]), 
        .SI(aes_state_regs_0_n147), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[2]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_2_ ( .D(aes_state_regs_0_n146), .SI(
        aes_state_regs_0_S30xDP_2_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n147), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_2_ ( .D(aes_state_regs_0_n144), .SI(
        aes_state_regs_0_S02xDP_2_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n146), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_2_ ( .D(StateInxD[2]), .SI(
        aes_state_regs_0_n144), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n145), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_2_ ( .D(aes_state_regs_0_S03xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n144), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_2_ ( .D(aes_state_regs_0_S23xDP_2_), 
        .SI(aes_state_regs_0_S20xDP_2_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[2]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_2_ ( .D(aes_state_regs_0_S20xDN[2]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_2_), .QN(
        aes_state_regs_0_n49) );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_1_ ( .D(aes_state_regs_0_S01xDO_1_), 
        .SI(StateInxD[1]), .SE(aes_state_regs_0_n177), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_1_), .QN(aes_state_regs_0_n42) );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_1_ ( .D(aes_state_regs_0_n143), .SI(
        aes_state_regs_0_n140), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S21xDP[1]), .QN(aes_state_regs_0_n121) );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_1_ ( .D(aes_state_regs_0_S02xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_1_ ( .D(aes_state_regs_0_n142), .SI(
        aes_state_regs_0_S23xDP_1_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_1_ ( .D(aes_state_regs_0_n140), .SI(
        aes_state_regs_0_n143), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_S23xDP_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_1_ ( .D(aes_state_regs_0_S02xDP_1_), 
        .SI(aes_state_regs_0_S01xDO_1_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n143), .QN() );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_1_ ( .D(aes_state_regs_0_S01xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_1_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_1_ ( .D(aes_state_regs_0_S21xDP[1]), 
        .SI(aes_state_regs_0_n142), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[1]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_1_ ( .D(aes_state_regs_0_n141), .SI(
        aes_state_regs_0_S30xDP_1_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n142), .QN() );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_1_ ( .D(aes_state_regs_0_n139), .SI(
        aes_state_regs_0_S02xDP_1_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n141), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_1_ ( .D(StateInxD[1]), .SI(
        aes_state_regs_0_n139), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(
        RstxBI), .Q(aes_state_regs_0_n140), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_1_ ( .D(aes_state_regs_0_S03xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n139), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_1_ ( .D(aes_state_regs_0_S23xDP_1_), 
        .SI(aes_state_regs_0_S20xDP_1_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[1]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_1_ ( .D(aes_state_regs_0_S20xDN[1]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_1_), .QN(
        aes_state_regs_0_n50) );
  SDFFR_X1 aes_state_regs_0_S00xDP_reg_0_ ( .D(
        aes_state_regs_0_MixColumnsS1xD[0]), .SI(aes_state_regs_0_S10xDP_0_), 
        .SE(aes_state_regs_0_n109), .CK(ClkxCI), .RN(RstxBI), .Q(
        aes_state_regs_0_S00xDP[0]), .QN(aes_state_regs_0_n35) );
  DFFR_X1 aes_state_regs_0_S10xDP_reg_0_ ( .D(aes_state_regs_0_S10xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S10xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S23xDP_reg_0_ ( .D(aes_state_regs_0_n137), .SI(
        aes_state_regs_0_S31xDP_0_), .SE(aes_state_regs_0_n177), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S23xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S31xDP_reg_0_ ( .D(aes_state_regs_0_S02xDP_0_), 
        .SI(aes_state_regs_0_S01xDO_0_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S31xDP_0_), .QN() );
  DFFR_X1 aes_state_regs_0_S02xDP_reg_0_ ( .D(aes_state_regs_0_S02xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S12xDP_reg_0_ ( .D(aes_state_regs_0_S22xDP_0_), 
        .SI(aes_state_regs_0_S23xDP_0_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S02xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_0_S22xDP_reg_0_ ( .D(aes_state_regs_0_n136), .SI(
        aes_state_regs_0_S30xDP_0_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S22xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S30xDP_reg_0_ ( .D(aes_state_regs_0_S01xDO_0_), 
        .SI(StateInxD[0]), .SE(aes_state_regs_0_n176), .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S30xDP_0_), .QN(aes_state_regs_0_n43) );
  DFFR_X1 aes_state_regs_0_S01xDP_reg_0_ ( .D(aes_state_regs_0_S01xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S01xDO_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S11xDP_reg_0_ ( .D(aes_state_regs_0_n138), .SI(
        aes_state_regs_0_S22xDP_0_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_S01xDN[0]), .QN() );
  SDFFR_X1 aes_state_regs_0_S21xDP_reg_0_ ( .D(aes_state_regs_0_S31xDP_0_), 
        .SI(aes_state_regs_0_n137), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n138), .QN() );
  SDFFR_X1 aes_state_regs_0_S33xDP_reg_0_ ( .D(StateInxD[0]), .SI(
        aes_state_regs_0_S03xDP_0_), .SE(aes_state_regs_0_n176), .CK(ClkxCI), 
        .RN(RstxBI), .Q(aes_state_regs_0_n137), .QN() );
  DFFR_X1 aes_state_regs_0_S03xDP_reg_0_ ( .D(aes_state_regs_0_S03xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDP_0_), .QN() );
  SDFFR_X1 aes_state_regs_0_S13xDP_reg_0_ ( .D(aes_state_regs_0_S23xDP_0_), 
        .SI(aes_state_regs_0_S20xDP_0_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S03xDN[0]), .QN() );
  DFFR_X1 aes_state_regs_0_S20xDP_reg_0_ ( .D(aes_state_regs_0_S20xDN[0]), 
        .CK(ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_S20xDP_0_), .QN(
        aes_state_regs_0_n51) );
  SDFFR_X1 aes_state_regs_0_S32xDP_reg_0_ ( .D(aes_state_regs_0_S03xDP_0_), 
        .SI(aes_state_regs_0_S02xDP_0_), .SE(aes_state_regs_0_n176), .CK(
        ClkxCI), .RN(RstxBI), .Q(aes_state_regs_0_n136), .QN() );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U119 ( .A(
        aes_state_regs_0_mix_columns_1_n245), .B(
        aes_state_regs_0_mix_columns_1_n244), .ZN(
        aes_state_regs_0_MixColumnsS3xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U118 ( .A(
        aes_state_regs_0_mix_columns_1_n240), .B(
        aes_state_regs_0_mix_columns_1_n239), .ZN(
        aes_state_regs_0_MixColumnsS3xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U117 ( .A(
        aes_state_regs_0_mix_columns_1_n235), .B(
        aes_state_regs_0_mix_columns_1_n234), .ZN(
        aes_state_regs_0_MixColumnsS3xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U116 ( .A(
        aes_state_regs_0_mix_columns_1_n226), .B(
        aes_state_regs_0_mix_columns_1_n225), .ZN(
        aes_state_regs_0_MixColumnsS3xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U115 ( .A(
        aes_state_regs_0_mix_columns_1_n183), .B(
        aes_state_regs_0_mix_columns_1_n196), .ZN(
        aes_state_regs_0_MixColumnsS1xD[1]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U114 ( .A(
        aes_state_regs_0_mix_columns_1_n191), .B(aes_state_regs_0_S00xDP[1]), 
        .ZN(aes_state_regs_0_mix_columns_1_n183) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U113 ( .A(
        aes_state_regs_0_mix_columns_1_n182), .B(
        aes_state_regs_0_mix_columns_1_n203), .ZN(
        aes_state_regs_0_MixColumnsS1xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U112 ( .A(aes_state_regs_0_S20xDP_3_), .B(aes_state_regs_0_mix_columns_1_n192), .ZN(
        aes_state_regs_0_mix_columns_1_n182) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U111 ( .A(
        aes_state_regs_0_mix_columns_1_n207), .B(
        aes_state_regs_0_mix_columns_1_n181), .ZN(
        aes_state_regs_0_mix_columns_1_n231) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U110 ( .A1(
        aes_state_regs_0_S30xDP_3_), .A2(aes_state_regs_0_mix_columns_1_n206), 
        .B1(aes_state_regs_0_S30xDP_7_), .B2(
        aes_state_regs_0_mix_columns_1_n180), .ZN(
        aes_state_regs_0_mix_columns_1_n181) );
  INV_X1 aes_state_regs_0_mix_columns_1_U109 ( .A(aes_state_regs_0_S30xDP_3_), 
        .ZN(aes_state_regs_0_mix_columns_1_n180) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U108 ( .A(
        aes_state_regs_0_mix_columns_1_n179), .B(
        aes_state_regs_0_mix_columns_1_n241), .ZN(
        aes_state_regs_0_MixColumnsS1xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U107 ( .A(
        aes_state_regs_0_mix_columns_1_n190), .B(aes_state_regs_0_S00xDP[0]), 
        .ZN(aes_state_regs_0_mix_columns_1_n179) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U106 ( .A(
        aes_state_regs_0_mix_columns_1_n177), .B(
        aes_state_regs_0_mix_columns_1_n178), .ZN(
        aes_state_regs_0_MixColumnsS1xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U105 ( .A(aes_state_regs_0_S20xDP_1_), .B(aes_state_regs_0_S10xDP_1_), .ZN(aes_state_regs_0_mix_columns_1_n178) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U104 ( .A(
        aes_state_regs_0_mix_columns_1_n200), .B(aes_state_regs_0_S20xDP_2_), 
        .Z(aes_state_regs_0_mix_columns_1_n177) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U103 ( .A(
        aes_state_regs_0_mix_columns_1_n176), .B(
        aes_state_regs_0_mix_columns_1_n205), .ZN(
        aes_state_regs_0_MixColumnsS1xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U102 ( .A(
        aes_state_regs_0_mix_columns_1_n193), .B(aes_state_regs_0_S00xDP[4]), 
        .ZN(aes_state_regs_0_mix_columns_1_n176) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U101 ( .A(
        aes_state_regs_0_mix_columns_1_n175), .B(
        aes_state_regs_0_mix_columns_1_n215), .ZN(
        aes_state_regs_0_MixColumnsS0xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U100 ( .A(aes_state_regs_0_S10xDP_6_), .B(aes_state_regs_0_mix_columns_1_n233), .ZN(
        aes_state_regs_0_mix_columns_1_n175) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U99 ( .A(
        aes_state_regs_0_mix_columns_1_n173), .B(
        aes_state_regs_0_mix_columns_1_n174), .ZN(
        aes_state_regs_0_MixColumnsS1xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U98 ( .A(aes_state_regs_0_S20xDP_4_), 
        .B(aes_state_regs_0_S10xDP_4_), .ZN(
        aes_state_regs_0_mix_columns_1_n174) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U97 ( .A(aes_state_regs_0_S00xDP[5]), 
        .B(aes_state_regs_0_mix_columns_1_n211), .Z(
        aes_state_regs_0_mix_columns_1_n173) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U96 ( .A(
        aes_state_regs_0_mix_columns_1_n172), .B(
        aes_state_regs_0_mix_columns_1_n171), .ZN(
        aes_state_regs_0_MixColumnsS1xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U95 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n217), .ZN(
        aes_state_regs_0_mix_columns_1_n172) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U94 ( .A1(aes_state_regs_0_S20xDP_6_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n236), .ZN(
        aes_state_regs_0_mix_columns_1_n171) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U93 ( .A(
        aes_state_regs_0_mix_columns_1_n169), .B(
        aes_state_regs_0_mix_columns_1_n170), .ZN(
        aes_state_regs_0_MixColumnsS1xD[6]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U92 ( .A(aes_state_regs_0_S20xDP_5_), 
        .B(aes_state_regs_0_S10xDP_5_), .ZN(
        aes_state_regs_0_mix_columns_1_n170) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U91 ( .A(aes_state_regs_0_S00xDP[6]), 
        .B(aes_state_regs_0_mix_columns_1_n215), .Z(
        aes_state_regs_0_mix_columns_1_n169) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U90 ( .A1(aes_state_regs_0_S20xDP_3_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n168), .ZN(
        aes_state_regs_0_mix_columns_1_n205) );
  INV_X1 aes_state_regs_0_mix_columns_1_U89 ( .A(aes_state_regs_0_S20xDP_3_), 
        .ZN(aes_state_regs_0_mix_columns_1_n168) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U88 ( .A(
        aes_state_regs_0_mix_columns_1_n167), .B(
        aes_state_regs_0_mix_columns_1_n190), .ZN(
        aes_state_regs_0_MixColumnsS0xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U87 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_mix_columns_1_n184), .ZN(
        aes_state_regs_0_mix_columns_1_n167) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U86 ( .A1(aes_state_regs_0_S30xDP_2_), .A2(aes_state_regs_0_S30xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n206), 
        .B2(aes_state_regs_0_mix_columns_1_n166), .ZN(
        aes_state_regs_0_mix_columns_1_n228) );
  INV_X1 aes_state_regs_0_mix_columns_1_U85 ( .A(aes_state_regs_0_S30xDP_2_), 
        .ZN(aes_state_regs_0_mix_columns_1_n166) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U84 ( .A(
        aes_state_regs_0_mix_columns_1_n164), .B(
        aes_state_regs_0_mix_columns_1_n165), .ZN(
        aes_state_regs_0_mix_columns_1_n227) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U83 ( .A(aes_state_regs_0_S20xDP_3_), 
        .B(aes_state_regs_0_S00xDP[7]), .ZN(
        aes_state_regs_0_mix_columns_1_n165) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U82 ( .A(aes_state_regs_0_S00xDP[2]), 
        .B(aes_state_regs_0_S10xDP_3_), .Z(aes_state_regs_0_mix_columns_1_n164) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U81 ( .A(
        aes_state_regs_0_mix_columns_1_n163), .B(
        aes_state_regs_0_mix_columns_1_n162), .ZN(
        aes_state_regs_0_mix_columns_1_n203) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U80 ( .A(aes_state_regs_0_S20xDP_2_), 
        .B(aes_state_regs_0_S30xDP_3_), .ZN(
        aes_state_regs_0_mix_columns_1_n163) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U79 ( .A1(aes_state_regs_0_S00xDP[3]), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n161), .ZN(
        aes_state_regs_0_mix_columns_1_n162) );
  INV_X1 aes_state_regs_0_mix_columns_1_U78 ( .A(aes_state_regs_0_S00xDP[3]), 
        .ZN(aes_state_regs_0_mix_columns_1_n161) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U77 ( .A(
        aes_state_regs_0_mix_columns_1_n160), .B(
        aes_state_regs_0_mix_columns_1_n209), .ZN(
        aes_state_regs_0_mix_columns_1_n193) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U76 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_3_), .ZN(
        aes_state_regs_0_mix_columns_1_n160) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U75 ( .A(
        aes_state_regs_0_mix_columns_1_n159), .B(
        aes_state_regs_0_mix_columns_1_n211), .ZN(
        aes_state_regs_0_MixColumnsS0xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U74 ( .A(aes_state_regs_0_S10xDP_5_), 
        .B(aes_state_regs_0_mix_columns_1_n207), .ZN(
        aes_state_regs_0_mix_columns_1_n159) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U73 ( .A1(aes_state_regs_0_S20xDP_0_), .A2(aes_state_regs_0_mix_columns_1_n218), .B1(
        aes_state_regs_0_mix_columns_1_n217), .B2(
        aes_state_regs_0_mix_columns_1_n216), .ZN(
        aes_state_regs_0_mix_columns_1_n219) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U72 ( .A(
        aes_state_regs_0_mix_columns_1_n220), .B(
        aes_state_regs_0_mix_columns_1_n219), .ZN(
        aes_state_regs_0_MixColumnsS3xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U71 ( .A(aes_state_regs_0_S20xDP_7_), 
        .B(aes_state_regs_0_mix_columns_1_n197), .ZN(
        aes_state_regs_0_mix_columns_1_n195) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U70 ( .A(
        aes_state_regs_0_mix_columns_1_n195), .B(
        aes_state_regs_0_mix_columns_1_n220), .ZN(
        aes_state_regs_0_MixColumnsS2xD[0]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U69 ( .A(
        aes_state_regs_0_mix_columns_1_n221), .B(aes_state_regs_0_S20xDP_1_), 
        .ZN(aes_state_regs_0_mix_columns_1_n223) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U68 ( .A(
        aes_state_regs_0_mix_columns_1_n223), .B(
        aes_state_regs_0_mix_columns_1_n222), .ZN(
        aes_state_regs_0_MixColumnsS3xD[1]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U67 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n224), .ZN(
        aes_state_regs_0_mix_columns_1_n225) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U66 ( .A(aes_state_regs_0_S00xDP[2]), 
        .B(aes_state_regs_0_S00xDP[1]), .Z(aes_state_regs_0_mix_columns_1_n226) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U65 ( .A(
        aes_state_regs_0_mix_columns_1_n227), .B(aes_state_regs_0_S00xDP[3]), 
        .ZN(aes_state_regs_0_mix_columns_1_n229) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U64 ( .A(
        aes_state_regs_0_mix_columns_1_n229), .B(
        aes_state_regs_0_mix_columns_1_n228), .ZN(
        aes_state_regs_0_MixColumnsS3xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U63 ( .A(
        aes_state_regs_0_mix_columns_1_n230), .B(aes_state_regs_0_S20xDP_4_), 
        .ZN(aes_state_regs_0_mix_columns_1_n232) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U62 ( .A(
        aes_state_regs_0_mix_columns_1_n232), .B(
        aes_state_regs_0_mix_columns_1_n231), .ZN(
        aes_state_regs_0_MixColumnsS3xD[4]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U61 ( .A(
        aes_state_regs_0_mix_columns_1_n233), .B(aes_state_regs_0_S20xDP_5_), 
        .Z(aes_state_regs_0_mix_columns_1_n235) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U60 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_S00xDP[4]), .ZN(
        aes_state_regs_0_mix_columns_1_n234) );
  INV_X1 aes_state_regs_0_mix_columns_1_U59 ( .A(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_mix_columns_1_n237) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U58 ( .A1(aes_state_regs_0_S20xDP_6_), .A2(aes_state_regs_0_mix_columns_1_n238), .B1(
        aes_state_regs_0_mix_columns_1_n237), .B2(
        aes_state_regs_0_mix_columns_1_n236), .ZN(
        aes_state_regs_0_mix_columns_1_n239) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U57 ( .A(aes_state_regs_0_S30xDP_5_), 
        .B(aes_state_regs_0_S00xDP[5]), .ZN(
        aes_state_regs_0_mix_columns_1_n240) );
  INV_X1 aes_state_regs_0_mix_columns_1_U56 ( .A(aes_state_regs_0_S00xDP[6]), 
        .ZN(aes_state_regs_0_mix_columns_1_n243) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U55 ( .A(aes_state_regs_0_S30xDP_6_), 
        .B(aes_state_regs_0_mix_columns_1_n241), .ZN(
        aes_state_regs_0_mix_columns_1_n245) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U54 ( .A1(aes_state_regs_0_S00xDP[7]), .A2(aes_state_regs_0_S00xDP[6]), .B1(aes_state_regs_0_mix_columns_1_n243), 
        .B2(aes_state_regs_0_mix_columns_1_n242), .ZN(
        aes_state_regs_0_mix_columns_1_n244) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U53 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n196), .ZN(
        aes_state_regs_0_mix_columns_1_n199) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U52 ( .A(
        aes_state_regs_0_mix_columns_1_n199), .B(
        aes_state_regs_0_mix_columns_1_n222), .ZN(
        aes_state_regs_0_MixColumnsS2xD[1]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U51 ( .A(aes_state_regs_0_S10xDP_2_), 
        .B(aes_state_regs_0_mix_columns_1_n200), .Z(
        aes_state_regs_0_mix_columns_1_n201) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U50 ( .A(
        aes_state_regs_0_mix_columns_1_n202), .B(
        aes_state_regs_0_mix_columns_1_n201), .ZN(
        aes_state_regs_0_MixColumnsS2xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U49 ( .A(aes_state_regs_0_S10xDP_3_), 
        .B(aes_state_regs_0_mix_columns_1_n203), .ZN(
        aes_state_regs_0_mix_columns_1_n204) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U48 ( .A(
        aes_state_regs_0_mix_columns_1_n204), .B(
        aes_state_regs_0_mix_columns_1_n228), .ZN(
        aes_state_regs_0_MixColumnsS2xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U47 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_mix_columns_1_n205), .ZN(
        aes_state_regs_0_mix_columns_1_n208) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U46 ( .A(
        aes_state_regs_0_mix_columns_1_n208), .B(
        aes_state_regs_0_mix_columns_1_n231), .ZN(
        aes_state_regs_0_MixColumnsS2xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U45 ( .A(
        aes_state_regs_0_mix_columns_1_n209), .B(aes_state_regs_0_S30xDP_5_), 
        .ZN(aes_state_regs_0_mix_columns_1_n210) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U44 ( .A(
        aes_state_regs_0_mix_columns_1_n210), .B(
        aes_state_regs_0_mix_columns_1_n233), .ZN(
        aes_state_regs_0_MixColumnsS2xD[5]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U43 ( .A(
        aes_state_regs_0_mix_columns_1_n211), .B(aes_state_regs_0_S30xDP_6_), 
        .ZN(aes_state_regs_0_mix_columns_1_n212) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U42 ( .A(
        aes_state_regs_0_mix_columns_1_n212), .B(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_MixColumnsS2xD[6]) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U41 ( .A1(aes_state_regs_0_S10xDP_7_), .A2(aes_state_regs_0_mix_columns_1_n218), .B1(
        aes_state_regs_0_mix_columns_1_n217), .B2(
        aes_state_regs_0_mix_columns_1_n213), .ZN(
        aes_state_regs_0_mix_columns_1_n214) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U40 ( .A(
        aes_state_regs_0_mix_columns_1_n215), .B(
        aes_state_regs_0_mix_columns_1_n214), .ZN(
        aes_state_regs_0_MixColumnsS2xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U39 ( .A(
        aes_state_regs_0_mix_columns_1_n241), .B(
        aes_state_regs_0_mix_columns_1_n238), .ZN(
        aes_state_regs_0_mix_columns_1_n189) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U38 ( .A(
        aes_state_regs_0_mix_columns_1_n189), .B(aes_state_regs_0_S30xDP_7_), 
        .ZN(aes_state_regs_0_MixColumnsS0xD[7]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U37 ( .A(aes_state_regs_0_S10xDP_4_), 
        .B(aes_state_regs_0_mix_columns_1_n230), .ZN(
        aes_state_regs_0_mix_columns_1_n188) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U36 ( .A(
        aes_state_regs_0_mix_columns_1_n188), .B(
        aes_state_regs_0_mix_columns_1_n193), .ZN(
        aes_state_regs_0_MixColumnsS0xD[4]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U35 ( .A(aes_state_regs_0_S30xDP_3_), 
        .B(aes_state_regs_0_mix_columns_1_n227), .ZN(
        aes_state_regs_0_mix_columns_1_n187) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U34 ( .A(
        aes_state_regs_0_mix_columns_1_n187), .B(
        aes_state_regs_0_mix_columns_1_n192), .ZN(
        aes_state_regs_0_MixColumnsS0xD[3]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U33 ( .A(aes_state_regs_0_S30xDP_2_), 
        .B(aes_state_regs_0_mix_columns_1_n224), .ZN(
        aes_state_regs_0_mix_columns_1_n186) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U32 ( .A(
        aes_state_regs_0_mix_columns_1_n186), .B(
        aes_state_regs_0_mix_columns_1_n198), .ZN(
        aes_state_regs_0_MixColumnsS0xD[2]) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U31 ( .A(aes_state_regs_0_S10xDP_1_), 
        .B(aes_state_regs_0_mix_columns_1_n221), .ZN(
        aes_state_regs_0_mix_columns_1_n185) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U30 ( .A(
        aes_state_regs_0_mix_columns_1_n185), .B(
        aes_state_regs_0_mix_columns_1_n191), .ZN(
        aes_state_regs_0_MixColumnsS0xD[1]) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U29 ( .A(aes_state_regs_0_S10xDP_0_), 
        .B(aes_state_regs_0_S00xDP[0]), .Z(aes_state_regs_0_mix_columns_1_n220) );
  INV_X1 aes_state_regs_0_mix_columns_1_U28 ( .A(
        aes_state_regs_0_mix_columns_1_n217), .ZN(
        aes_state_regs_0_mix_columns_1_n218) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U27 ( .A1(aes_state_regs_0_S00xDP[7]), .A2(aes_state_regs_0_S30xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n206), 
        .B2(aes_state_regs_0_mix_columns_1_n242), .ZN(
        aes_state_regs_0_mix_columns_1_n217) );
  INV_X1 aes_state_regs_0_mix_columns_1_U26 ( .A(aes_state_regs_0_S20xDP_0_), 
        .ZN(aes_state_regs_0_mix_columns_1_n216) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U25 ( .A(aes_state_regs_0_S30xDP_0_), 
        .B(aes_state_regs_0_mix_columns_1_n206), .ZN(
        aes_state_regs_0_mix_columns_1_n197) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U24 ( .A1(aes_state_regs_0_S10xDP_7_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n213), .ZN(
        aes_state_regs_0_mix_columns_1_n241) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U23 ( .A(aes_state_regs_0_S30xDP_0_), 
        .B(aes_state_regs_0_S20xDP_0_), .Z(aes_state_regs_0_mix_columns_1_n190) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U22 ( .A(
        aes_state_regs_0_mix_columns_1_n198), .B(
        aes_state_regs_0_mix_columns_1_n197), .Z(
        aes_state_regs_0_mix_columns_1_n222) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U21 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_S00xDP[0]), .Z(aes_state_regs_0_mix_columns_1_n221) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U20 ( .A(aes_state_regs_0_S10xDP_2_), 
        .B(aes_state_regs_0_S20xDP_2_), .Z(aes_state_regs_0_mix_columns_1_n224) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U19 ( .A(aes_state_regs_0_S00xDP[7]), 
        .B(aes_state_regs_0_S00xDP[3]), .Z(aes_state_regs_0_mix_columns_1_n230) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U18 ( .A(aes_state_regs_0_S10xDP_5_), 
        .B(aes_state_regs_0_S00xDP[5]), .Z(aes_state_regs_0_mix_columns_1_n233) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U17 ( .A(aes_state_regs_0_S10xDP_6_), 
        .B(aes_state_regs_0_S00xDP[6]), .Z(aes_state_regs_0_mix_columns_1_n238) );
  INV_X1 aes_state_regs_0_mix_columns_1_U16 ( .A(aes_state_regs_0_S20xDP_6_), 
        .ZN(aes_state_regs_0_mix_columns_1_n236) );
  INV_X1 aes_state_regs_0_mix_columns_1_U15 ( .A(aes_state_regs_0_S00xDP[7]), 
        .ZN(aes_state_regs_0_mix_columns_1_n242) );
  AOI22_X1 aes_state_regs_0_mix_columns_1_U14 ( .A1(aes_state_regs_0_S20xDP_0_), .A2(aes_state_regs_0_S20xDP_7_), .B1(aes_state_regs_0_mix_columns_1_n194), 
        .B2(aes_state_regs_0_mix_columns_1_n216), .ZN(
        aes_state_regs_0_mix_columns_1_n196) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U13 ( .A(aes_state_regs_0_S30xDP_2_), 
        .B(aes_state_regs_0_S00xDP[2]), .Z(aes_state_regs_0_mix_columns_1_n200) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U12 ( .A(aes_state_regs_0_S30xDP_1_), 
        .B(aes_state_regs_0_S20xDP_1_), .ZN(
        aes_state_regs_0_mix_columns_1_n202) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U11 ( .A(aes_state_regs_0_S30xDP_4_), 
        .B(aes_state_regs_0_S20xDP_4_), .Z(aes_state_regs_0_mix_columns_1_n209) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U10 ( .A(aes_state_regs_0_S30xDP_5_), 
        .B(aes_state_regs_0_S20xDP_5_), .Z(aes_state_regs_0_mix_columns_1_n211) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U9 ( .A(aes_state_regs_0_S30xDP_6_), 
        .B(aes_state_regs_0_S20xDP_6_), .Z(aes_state_regs_0_mix_columns_1_n215) );
  INV_X1 aes_state_regs_0_mix_columns_1_U8 ( .A(aes_state_regs_0_S10xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n213) );
  XNOR2_X1 aes_state_regs_0_mix_columns_1_U7 ( .A(
        aes_state_regs_0_mix_columns_1_n184), .B(
        aes_state_regs_0_mix_columns_1_n202), .ZN(
        aes_state_regs_0_mix_columns_1_n191) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U6 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_2_), .Z(aes_state_regs_0_mix_columns_1_n192) );
  INV_X1 aes_state_regs_0_mix_columns_1_U5 ( .A(aes_state_regs_0_S20xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n194) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U4 ( .A(aes_state_regs_0_S10xDP_1_), 
        .B(aes_state_regs_0_S00xDP[1]), .Z(aes_state_regs_0_mix_columns_1_n198) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U3 ( .A(aes_state_regs_0_S10xDP_7_), 
        .B(aes_state_regs_0_S10xDP_0_), .Z(aes_state_regs_0_mix_columns_1_n184) );
  INV_X1 aes_state_regs_0_mix_columns_1_U2 ( .A(aes_state_regs_0_S30xDP_7_), 
        .ZN(aes_state_regs_0_mix_columns_1_n206) );
  XOR2_X1 aes_state_regs_0_mix_columns_1_U1 ( .A(aes_state_regs_0_S10xDP_4_), 
        .B(aes_state_regs_0_S00xDP[4]), .Z(aes_state_regs_0_mix_columns_1_n207) );
endmodule

