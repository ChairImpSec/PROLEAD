
module circuit ( clk, nReset, dataIn1, dataIn2, key, dataOut1, dataOut2, done
 );
  input [3:0] dataIn1;
  input [3:0] dataIn2;
  input [3:0] key;
  output [3:0] dataOut1;
  output [3:0] dataOut2;
  input clk, nReset;
  output done;
  wire   selInit, selP, enKey, fsm_n21, fsm_n20, fsm_n19, fsm_n18, fsm_n15,
         fsm_n14, fsm_n12, fsm_n11, fsm_n10, fsm_n9, fsm_n7, fsm_n13, fsm_n17,
         fsm_n16, fsm_ps_state_0_, fsm_ps_state_1_, fsm_ps_state_2_,
         fsm_rst_countSerial, fsm_en_countRound, fsm_cnt_rnd_n40,
         fsm_cnt_rnd_n39, fsm_cnt_rnd_n38, fsm_cnt_rnd_n37, fsm_cnt_rnd_n36,
         fsm_cnt_rnd_n35, fsm_cnt_rnd_n34, fsm_cnt_rnd_n33, fsm_cnt_rnd_n32,
         fsm_cnt_rnd_n31, fsm_cnt_rnd_n30, fsm_cnt_rnd_n29, fsm_cnt_rnd_n28,
         fsm_cnt_rnd_n27, fsm_cnt_rnd_n26, fsm_cnt_rnd_n24, fsm_cnt_rnd_n19,
         fsm_cnt_rnd_n18, fsm_cnt_rnd_n23, fsm_cnt_rnd_n22, fsm_cnt_rnd_n21,
         fsm_cnt_rnd_n20, fsm_cnt_rnd_n5, fsm_cnt_ser_n21, fsm_cnt_ser_n16,
         fsm_cnt_ser_n15, fsm_cnt_ser_n14, fsm_cnt_ser_n13, fsm_cnt_ser_n12,
         fsm_cnt_ser_n11, fsm_cnt_ser_n10, fsm_cnt_ser_n9, fsm_cnt_ser_n20,
         fsm_cnt_ser_n19, fsm_cnt_ser_n18, fsm_cnt_ser_n17, stateFF_n1,
         stateFF_state_n11, stateFF_state_n10, stateFF_state_n9,
         stateFF_state_n8, stateFF_state_n7, stateFF_state_n6,
         stateFF_state_gff_1_n2, stateFF_state_gff_1_SFF_0_n9,
         stateFF_state_gff_1_SFF_0_n7, stateFF_state_gff_1_SFF_0_n6,
         stateFF_state_gff_1_SFF_1_n11, stateFF_state_gff_1_SFF_1_n10,
         stateFF_state_gff_1_SFF_1_n8, stateFF_state_gff_1_SFF_1_n7,
         stateFF_state_gff_1_SFF_2_n11, stateFF_state_gff_1_SFF_2_n10,
         stateFF_state_gff_1_SFF_2_n8, stateFF_state_gff_1_SFF_2_n7,
         stateFF_state_gff_1_SFF_3_n11, stateFF_state_gff_1_SFF_3_n10,
         stateFF_state_gff_1_SFF_3_n8, stateFF_state_gff_1_SFF_3_n7,
         stateFF_state_gff_2_SFF_0_n12, stateFF_state_gff_2_SFF_0_n11,
         stateFF_state_gff_2_SFF_0_n10, stateFF_state_gff_2_SFF_0_n8,
         stateFF_state_gff_2_SFF_0_n7, stateFF_state_gff_2_SFF_1_n12,
         stateFF_state_gff_2_SFF_1_n11, stateFF_state_gff_2_SFF_1_n10,
         stateFF_state_gff_2_SFF_1_n8, stateFF_state_gff_2_SFF_1_n7,
         stateFF_state_gff_2_SFF_2_n12, stateFF_state_gff_2_SFF_2_n11,
         stateFF_state_gff_2_SFF_2_n10, stateFF_state_gff_2_SFF_2_n8,
         stateFF_state_gff_2_SFF_2_n7, stateFF_state_gff_2_SFF_3_n12,
         stateFF_state_gff_2_SFF_3_n11, stateFF_state_gff_2_SFF_3_n10,
         stateFF_state_gff_2_SFF_3_n8, stateFF_state_gff_2_SFF_3_n7,
         stateFF_state_gff_3_SFF_0_n11, stateFF_state_gff_3_SFF_0_n10,
         stateFF_state_gff_3_SFF_0_n8, stateFF_state_gff_3_SFF_0_n7,
         stateFF_state_gff_3_SFF_1_n11, stateFF_state_gff_3_SFF_1_n10,
         stateFF_state_gff_3_SFF_1_n8, stateFF_state_gff_3_SFF_1_n7,
         stateFF_state_gff_3_SFF_2_n11, stateFF_state_gff_3_SFF_2_n10,
         stateFF_state_gff_3_SFF_2_n8, stateFF_state_gff_3_SFF_2_n7,
         stateFF_state_gff_3_SFF_3_n11, stateFF_state_gff_3_SFF_3_n10,
         stateFF_state_gff_3_SFF_3_n8, stateFF_state_gff_3_SFF_3_n7,
         stateFF_state_gff_4_SFF_0_n11, stateFF_state_gff_4_SFF_0_n10,
         stateFF_state_gff_4_SFF_0_n8, stateFF_state_gff_4_SFF_0_n7,
         stateFF_state_gff_4_SFF_1_n11, stateFF_state_gff_4_SFF_1_n10,
         stateFF_state_gff_4_SFF_1_n8, stateFF_state_gff_4_SFF_1_n7,
         stateFF_state_gff_4_SFF_2_n11, stateFF_state_gff_4_SFF_2_n10,
         stateFF_state_gff_4_SFF_2_n9, stateFF_state_gff_4_SFF_2_n7,
         stateFF_state_gff_4_SFF_2_n6, stateFF_state_gff_4_SFF_3_n11,
         stateFF_state_gff_4_SFF_3_n10, stateFF_state_gff_4_SFF_3_n9,
         stateFF_state_gff_4_SFF_3_n7, stateFF_state_gff_4_SFF_3_n6,
         stateFF_state_gff_5_SFF_0_n11, stateFF_state_gff_5_SFF_0_n10,
         stateFF_state_gff_5_SFF_0_n9, stateFF_state_gff_5_SFF_0_n7,
         stateFF_state_gff_5_SFF_0_n6, stateFF_state_gff_5_SFF_1_n11,
         stateFF_state_gff_5_SFF_1_n10, stateFF_state_gff_5_SFF_1_n9,
         stateFF_state_gff_5_SFF_1_n7, stateFF_state_gff_5_SFF_1_n6,
         stateFF_state_gff_5_SFF_2_n11, stateFF_state_gff_5_SFF_2_n10,
         stateFF_state_gff_5_SFF_2_n9, stateFF_state_gff_5_SFF_2_n7,
         stateFF_state_gff_5_SFF_2_n6, stateFF_state_gff_5_SFF_3_n11,
         stateFF_state_gff_5_SFF_3_n10, stateFF_state_gff_5_SFF_3_n9,
         stateFF_state_gff_5_SFF_3_n7, stateFF_state_gff_5_SFF_3_n6,
         stateFF_state_gff_6_n2, stateFF_state_gff_6_SFF_0_n11,
         stateFF_state_gff_6_SFF_0_n10, stateFF_state_gff_6_SFF_0_n8,
         stateFF_state_gff_6_SFF_0_n7, stateFF_state_gff_6_SFF_1_n10,
         stateFF_state_gff_6_SFF_1_n8, stateFF_state_gff_6_SFF_1_n7,
         stateFF_state_gff_6_SFF_2_n11, stateFF_state_gff_6_SFF_2_n10,
         stateFF_state_gff_6_SFF_2_n8, stateFF_state_gff_6_SFF_2_n7,
         stateFF_state_gff_6_SFF_3_n11, stateFF_state_gff_6_SFF_3_n10,
         stateFF_state_gff_6_SFF_3_n8, stateFF_state_gff_6_SFF_3_n7,
         stateFF_state_gff_7_SFF_0_n12, stateFF_state_gff_7_SFF_0_n11,
         stateFF_state_gff_7_SFF_0_n10, stateFF_state_gff_7_SFF_0_n8,
         stateFF_state_gff_7_SFF_0_n7, stateFF_state_gff_7_SFF_1_n12,
         stateFF_state_gff_7_SFF_1_n11, stateFF_state_gff_7_SFF_1_n10,
         stateFF_state_gff_7_SFF_1_n8, stateFF_state_gff_7_SFF_1_n7,
         stateFF_state_gff_7_SFF_2_n12, stateFF_state_gff_7_SFF_2_n11,
         stateFF_state_gff_7_SFF_2_n10, stateFF_state_gff_7_SFF_2_n8,
         stateFF_state_gff_7_SFF_2_n7, stateFF_state_gff_7_SFF_3_n12,
         stateFF_state_gff_7_SFF_3_n11, stateFF_state_gff_7_SFF_3_n10,
         stateFF_state_gff_7_SFF_3_n8, stateFF_state_gff_7_SFF_3_n7,
         stateFF_state_gff_8_SFF_0_n12, stateFF_state_gff_8_SFF_0_n11,
         stateFF_state_gff_8_SFF_0_n10, stateFF_state_gff_8_SFF_0_n8,
         stateFF_state_gff_8_SFF_0_n7, stateFF_state_gff_8_SFF_1_n12,
         stateFF_state_gff_8_SFF_1_n11, stateFF_state_gff_8_SFF_1_n10,
         stateFF_state_gff_8_SFF_1_n8, stateFF_state_gff_8_SFF_1_n7,
         stateFF_state_gff_8_SFF_2_n11, stateFF_state_gff_8_SFF_2_n10,
         stateFF_state_gff_8_SFF_2_n9, stateFF_state_gff_8_SFF_2_n7,
         stateFF_state_gff_8_SFF_2_n6, stateFF_state_gff_8_SFF_3_n11,
         stateFF_state_gff_8_SFF_3_n10, stateFF_state_gff_8_SFF_3_n9,
         stateFF_state_gff_8_SFF_3_n7, stateFF_state_gff_8_SFF_3_n6,
         stateFF_state_gff_9_SFF_0_n11, stateFF_state_gff_9_SFF_0_n10,
         stateFF_state_gff_9_SFF_0_n9, stateFF_state_gff_9_SFF_0_n7,
         stateFF_state_gff_9_SFF_0_n6, stateFF_state_gff_9_SFF_1_n11,
         stateFF_state_gff_9_SFF_1_n10, stateFF_state_gff_9_SFF_1_n9,
         stateFF_state_gff_9_SFF_1_n7, stateFF_state_gff_9_SFF_1_n6,
         stateFF_state_gff_9_SFF_2_n11, stateFF_state_gff_9_SFF_2_n10,
         stateFF_state_gff_9_SFF_2_n9, stateFF_state_gff_9_SFF_2_n7,
         stateFF_state_gff_9_SFF_2_n6, stateFF_state_gff_9_SFF_3_n11,
         stateFF_state_gff_9_SFF_3_n10, stateFF_state_gff_9_SFF_3_n9,
         stateFF_state_gff_9_SFF_3_n7, stateFF_state_gff_9_SFF_3_n6,
         stateFF_state_gff_10_SFF_0_n12, stateFF_state_gff_10_SFF_0_n11,
         stateFF_state_gff_10_SFF_0_n10, stateFF_state_gff_10_SFF_0_n8,
         stateFF_state_gff_10_SFF_0_n7, stateFF_state_gff_10_SFF_1_n12,
         stateFF_state_gff_10_SFF_1_n11, stateFF_state_gff_10_SFF_1_n10,
         stateFF_state_gff_10_SFF_1_n8, stateFF_state_gff_10_SFF_1_n7,
         stateFF_state_gff_10_SFF_2_n11, stateFF_state_gff_10_SFF_2_n10,
         stateFF_state_gff_10_SFF_2_n8, stateFF_state_gff_10_SFF_2_n7,
         stateFF_state_gff_10_SFF_3_n11, stateFF_state_gff_10_SFF_3_n10,
         stateFF_state_gff_10_SFF_3_n8, stateFF_state_gff_10_SFF_3_n7,
         stateFF_state_gff_11_n2, stateFF_state_gff_11_SFF_0_n11,
         stateFF_state_gff_11_SFF_0_n10, stateFF_state_gff_11_SFF_0_n8,
         stateFF_state_gff_11_SFF_0_n7, stateFF_state_gff_11_SFF_1_n11,
         stateFF_state_gff_11_SFF_1_n10, stateFF_state_gff_11_SFF_1_n8,
         stateFF_state_gff_11_SFF_1_n7, stateFF_state_gff_11_SFF_2_n10,
         stateFF_state_gff_11_SFF_2_n8, stateFF_state_gff_11_SFF_2_n7,
         stateFF_state_gff_11_SFF_3_n11, stateFF_state_gff_11_SFF_3_n10,
         stateFF_state_gff_11_SFF_3_n8, stateFF_state_gff_11_SFF_3_n7,
         stateFF_state_gff_12_SFF_0_n11, stateFF_state_gff_12_SFF_0_n10,
         stateFF_state_gff_12_SFF_0_n8, stateFF_state_gff_12_SFF_0_n7,
         stateFF_state_gff_12_SFF_1_n11, stateFF_state_gff_12_SFF_1_n10,
         stateFF_state_gff_12_SFF_1_n8, stateFF_state_gff_12_SFF_1_n7,
         stateFF_state_gff_12_SFF_2_n11, stateFF_state_gff_12_SFF_2_n10,
         stateFF_state_gff_12_SFF_2_n9, stateFF_state_gff_12_SFF_2_n7,
         stateFF_state_gff_12_SFF_2_n6, stateFF_state_gff_12_SFF_3_n11,
         stateFF_state_gff_12_SFF_3_n10, stateFF_state_gff_12_SFF_3_n9,
         stateFF_state_gff_12_SFF_3_n7, stateFF_state_gff_12_SFF_3_n6,
         stateFF_state_gff_13_SFF_0_n11, stateFF_state_gff_13_SFF_0_n10,
         stateFF_state_gff_13_SFF_0_n9, stateFF_state_gff_13_SFF_0_n7,
         stateFF_state_gff_13_SFF_0_n6, stateFF_state_gff_13_SFF_1_n11,
         stateFF_state_gff_13_SFF_1_n10, stateFF_state_gff_13_SFF_1_n9,
         stateFF_state_gff_13_SFF_1_n7, stateFF_state_gff_13_SFF_1_n6,
         stateFF_state_gff_13_SFF_2_n11, stateFF_state_gff_13_SFF_2_n10,
         stateFF_state_gff_13_SFF_2_n9, stateFF_state_gff_13_SFF_2_n7,
         stateFF_state_gff_13_SFF_2_n6, stateFF_state_gff_13_SFF_3_n11,
         stateFF_state_gff_13_SFF_3_n10, stateFF_state_gff_13_SFF_3_n9,
         stateFF_state_gff_13_SFF_3_n7, stateFF_state_gff_13_SFF_3_n6,
         stateFF_state_gff_14_SFF_0_n11, stateFF_state_gff_14_SFF_0_n10,
         stateFF_state_gff_14_SFF_0_n8, stateFF_state_gff_14_SFF_0_n7,
         stateFF_state_gff_14_SFF_1_n11, stateFF_state_gff_14_SFF_1_n10,
         stateFF_state_gff_14_SFF_1_n8, stateFF_state_gff_14_SFF_1_n7,
         stateFF_state_gff_14_SFF_2_n11, stateFF_state_gff_14_SFF_2_n10,
         stateFF_state_gff_14_SFF_2_n8, stateFF_state_gff_14_SFF_2_n7,
         stateFF_state_gff_14_SFF_3_n11, stateFF_state_gff_14_SFF_3_n10,
         stateFF_state_gff_14_SFF_3_n8, stateFF_state_gff_14_SFF_3_n7,
         stateFF_state_gff_15_SFF_0_n11, stateFF_state_gff_15_SFF_0_n10,
         stateFF_state_gff_15_SFF_0_n8, stateFF_state_gff_15_SFF_0_n7,
         stateFF_state_gff_15_SFF_1_n11, stateFF_state_gff_15_SFF_1_n10,
         stateFF_state_gff_15_SFF_1_n8, stateFF_state_gff_15_SFF_1_n7,
         stateFF_state_gff_15_SFF_2_n11, stateFF_state_gff_15_SFF_2_n10,
         stateFF_state_gff_15_SFF_2_n8, stateFF_state_gff_15_SFF_2_n7,
         stateFF_state_gff_15_SFF_3_n10, stateFF_state_gff_15_SFF_3_n9,
         stateFF_state_gff_15_SFF_3_n7, stateFF_state_gff_15_SFF_3_n6,
         stateFF_state_gff_16_n2, stateFF_state_gff_16_SFF_0_n10,
         stateFF_state_gff_16_SFF_0_n9, stateFF_state_gff_16_SFF_0_n7,
         stateFF_state_gff_16_SFF_0_n6, stateFF_state_gff_16_SFF_1_n10,
         stateFF_state_gff_16_SFF_1_n9, stateFF_state_gff_16_SFF_1_n7,
         stateFF_state_gff_16_SFF_1_n6, stateFF_state_gff_16_SFF_2_n10,
         stateFF_state_gff_16_SFF_2_n9, stateFF_state_gff_16_SFF_2_n7,
         stateFF_state_gff_16_SFF_2_n6, stateFF_state_gff_16_SFF_3_n9,
         stateFF_state_gff_16_SFF_3_n7, stateFF_state_gff_16_SFF_3_n6,
         md1FF_n3, md1FF_state_n12, md1FF_state_n11, md1FF_state_n10,
         md1FF_state_n9, md1FF_state_n8, md1FF_state_n7, md1FF_state_n6,
         md1FF_state_gff_1_n2, md1FF_state_gff_1_SFF_0_n10,
         md1FF_state_gff_1_SFF_0_n8, md1FF_state_gff_1_SFF_0_n7,
         md1FF_state_gff_1_SFF_1_n11, md1FF_state_gff_1_SFF_1_n10,
         md1FF_state_gff_1_SFF_1_n8, md1FF_state_gff_1_SFF_1_n7,
         md1FF_state_gff_1_SFF_2_n11, md1FF_state_gff_1_SFF_2_n10,
         md1FF_state_gff_1_SFF_2_n8, md1FF_state_gff_1_SFF_2_n7,
         md1FF_state_gff_1_SFF_3_n11, md1FF_state_gff_1_SFF_3_n10,
         md1FF_state_gff_1_SFF_3_n8, md1FF_state_gff_1_SFF_3_n7,
         md1FF_state_gff_2_SFF_0_n12, md1FF_state_gff_2_SFF_0_n11,
         md1FF_state_gff_2_SFF_0_n10, md1FF_state_gff_2_SFF_0_n8,
         md1FF_state_gff_2_SFF_0_n7, md1FF_state_gff_2_SFF_1_n12,
         md1FF_state_gff_2_SFF_1_n11, md1FF_state_gff_2_SFF_1_n10,
         md1FF_state_gff_2_SFF_1_n8, md1FF_state_gff_2_SFF_1_n7,
         md1FF_state_gff_2_SFF_2_n12, md1FF_state_gff_2_SFF_2_n11,
         md1FF_state_gff_2_SFF_2_n10, md1FF_state_gff_2_SFF_2_n8,
         md1FF_state_gff_2_SFF_2_n7, md1FF_state_gff_2_SFF_3_n12,
         md1FF_state_gff_2_SFF_3_n11, md1FF_state_gff_2_SFF_3_n10,
         md1FF_state_gff_2_SFF_3_n8, md1FF_state_gff_2_SFF_3_n7,
         md1FF_state_gff_3_SFF_0_n12, md1FF_state_gff_3_SFF_0_n11,
         md1FF_state_gff_3_SFF_0_n10, md1FF_state_gff_3_SFF_0_n8,
         md1FF_state_gff_3_SFF_0_n7, md1FF_state_gff_3_SFF_1_n12,
         md1FF_state_gff_3_SFF_1_n11, md1FF_state_gff_3_SFF_1_n10,
         md1FF_state_gff_3_SFF_1_n8, md1FF_state_gff_3_SFF_1_n7,
         md1FF_state_gff_3_SFF_2_n11, md1FF_state_gff_3_SFF_2_n10,
         md1FF_state_gff_3_SFF_2_n9, md1FF_state_gff_3_SFF_2_n7,
         md1FF_state_gff_3_SFF_2_n6, md1FF_state_gff_3_SFF_3_n11,
         md1FF_state_gff_3_SFF_3_n10, md1FF_state_gff_3_SFF_3_n9,
         md1FF_state_gff_3_SFF_3_n7, md1FF_state_gff_3_SFF_3_n6,
         md1FF_state_gff_4_SFF_0_n11, md1FF_state_gff_4_SFF_0_n10,
         md1FF_state_gff_4_SFF_0_n9, md1FF_state_gff_4_SFF_0_n7,
         md1FF_state_gff_4_SFF_0_n6, md1FF_state_gff_4_SFF_1_n11,
         md1FF_state_gff_4_SFF_1_n10, md1FF_state_gff_4_SFF_1_n9,
         md1FF_state_gff_4_SFF_1_n7, md1FF_state_gff_4_SFF_1_n6,
         md1FF_state_gff_4_SFF_2_n11, md1FF_state_gff_4_SFF_2_n10,
         md1FF_state_gff_4_SFF_2_n9, md1FF_state_gff_4_SFF_2_n7,
         md1FF_state_gff_4_SFF_2_n6, md1FF_state_gff_4_SFF_3_n11,
         md1FF_state_gff_4_SFF_3_n10, md1FF_state_gff_4_SFF_3_n9,
         md1FF_state_gff_4_SFF_3_n7, md1FF_state_gff_4_SFF_3_n6,
         md1FF_state_gff_5_SFF_0_n12, md1FF_state_gff_5_SFF_0_n11,
         md1FF_state_gff_5_SFF_0_n10, md1FF_state_gff_5_SFF_0_n8,
         md1FF_state_gff_5_SFF_0_n7, md1FF_state_gff_5_SFF_1_n12,
         md1FF_state_gff_5_SFF_1_n11, md1FF_state_gff_5_SFF_1_n10,
         md1FF_state_gff_5_SFF_1_n8, md1FF_state_gff_5_SFF_1_n7,
         md1FF_state_gff_5_SFF_2_n12, md1FF_state_gff_5_SFF_2_n11,
         md1FF_state_gff_5_SFF_2_n10, md1FF_state_gff_5_SFF_2_n8,
         md1FF_state_gff_5_SFF_2_n7, md1FF_state_gff_5_SFF_3_n12,
         md1FF_state_gff_5_SFF_3_n11, md1FF_state_gff_5_SFF_3_n10,
         md1FF_state_gff_5_SFF_3_n8, md1FF_state_gff_5_SFF_3_n7,
         md1FF_state_gff_6_n2, md1FF_state_gff_6_SFF_0_n11,
         md1FF_state_gff_6_SFF_0_n10, md1FF_state_gff_6_SFF_0_n8,
         md1FF_state_gff_6_SFF_0_n7, md1FF_state_gff_6_SFF_1_n10,
         md1FF_state_gff_6_SFF_1_n8, md1FF_state_gff_6_SFF_1_n7,
         md1FF_state_gff_6_SFF_2_n11, md1FF_state_gff_6_SFF_2_n10,
         md1FF_state_gff_6_SFF_2_n8, md1FF_state_gff_6_SFF_2_n7,
         md1FF_state_gff_6_SFF_3_n11, md1FF_state_gff_6_SFF_3_n10,
         md1FF_state_gff_6_SFF_3_n8, md1FF_state_gff_6_SFF_3_n7,
         md1FF_state_gff_7_SFF_0_n11, md1FF_state_gff_7_SFF_0_n10,
         md1FF_state_gff_7_SFF_0_n8, md1FF_state_gff_7_SFF_0_n7,
         md1FF_state_gff_7_SFF_1_n11, md1FF_state_gff_7_SFF_1_n10,
         md1FF_state_gff_7_SFF_1_n8, md1FF_state_gff_7_SFF_1_n7,
         md1FF_state_gff_7_SFF_2_n11, md1FF_state_gff_7_SFF_2_n10,
         md1FF_state_gff_7_SFF_2_n9, md1FF_state_gff_7_SFF_2_n7,
         md1FF_state_gff_7_SFF_2_n6, md1FF_state_gff_7_SFF_3_n11,
         md1FF_state_gff_7_SFF_3_n10, md1FF_state_gff_7_SFF_3_n9,
         md1FF_state_gff_7_SFF_3_n7, md1FF_state_gff_7_SFF_3_n6,
         md1FF_state_gff_8_SFF_0_n11, md1FF_state_gff_8_SFF_0_n10,
         md1FF_state_gff_8_SFF_0_n9, md1FF_state_gff_8_SFF_0_n7,
         md1FF_state_gff_8_SFF_0_n6, md1FF_state_gff_8_SFF_1_n11,
         md1FF_state_gff_8_SFF_1_n10, md1FF_state_gff_8_SFF_1_n9,
         md1FF_state_gff_8_SFF_1_n7, md1FF_state_gff_8_SFF_1_n6,
         md1FF_state_gff_8_SFF_2_n11, md1FF_state_gff_8_SFF_2_n10,
         md1FF_state_gff_8_SFF_2_n9, md1FF_state_gff_8_SFF_2_n7,
         md1FF_state_gff_8_SFF_2_n6, md1FF_state_gff_8_SFF_3_n11,
         md1FF_state_gff_8_SFF_3_n10, md1FF_state_gff_8_SFF_3_n9,
         md1FF_state_gff_8_SFF_3_n7, md1FF_state_gff_8_SFF_3_n6,
         md1FF_state_gff_9_SFF_0_n12, md1FF_state_gff_9_SFF_0_n11,
         md1FF_state_gff_9_SFF_0_n10, md1FF_state_gff_9_SFF_0_n8,
         md1FF_state_gff_9_SFF_0_n7, md1FF_state_gff_9_SFF_1_n12,
         md1FF_state_gff_9_SFF_1_n11, md1FF_state_gff_9_SFF_1_n10,
         md1FF_state_gff_9_SFF_1_n8, md1FF_state_gff_9_SFF_1_n7,
         md1FF_state_gff_9_SFF_2_n11, md1FF_state_gff_9_SFF_2_n10,
         md1FF_state_gff_9_SFF_2_n8, md1FF_state_gff_9_SFF_2_n7,
         md1FF_state_gff_9_SFF_3_n11, md1FF_state_gff_9_SFF_3_n10,
         md1FF_state_gff_9_SFF_3_n8, md1FF_state_gff_9_SFF_3_n7,
         md1FF_state_gff_10_SFF_0_n11, md1FF_state_gff_10_SFF_0_n10,
         md1FF_state_gff_10_SFF_0_n8, md1FF_state_gff_10_SFF_0_n7,
         md1FF_state_gff_10_SFF_1_n11, md1FF_state_gff_10_SFF_1_n10,
         md1FF_state_gff_10_SFF_1_n8, md1FF_state_gff_10_SFF_1_n7,
         md1FF_state_gff_10_SFF_2_n11, md1FF_state_gff_10_SFF_2_n10,
         md1FF_state_gff_10_SFF_2_n8, md1FF_state_gff_10_SFF_2_n7,
         md1FF_state_gff_10_SFF_3_n11, md1FF_state_gff_10_SFF_3_n10,
         md1FF_state_gff_10_SFF_3_n8, md1FF_state_gff_10_SFF_3_n7,
         md1FF_state_gff_11_n2, md1FF_state_gff_11_SFF_0_n11,
         md1FF_state_gff_11_SFF_0_n10, md1FF_state_gff_11_SFF_0_n8,
         md1FF_state_gff_11_SFF_0_n7, md1FF_state_gff_11_SFF_1_n11,
         md1FF_state_gff_11_SFF_1_n10, md1FF_state_gff_11_SFF_1_n8,
         md1FF_state_gff_11_SFF_1_n7, md1FF_state_gff_11_SFF_2_n9,
         md1FF_state_gff_11_SFF_2_n7, md1FF_state_gff_11_SFF_2_n6,
         md1FF_state_gff_11_SFF_3_n10, md1FF_state_gff_11_SFF_3_n9,
         md1FF_state_gff_11_SFF_3_n7, md1FF_state_gff_11_SFF_3_n6,
         md1FF_state_gff_12_SFF_0_n10, md1FF_state_gff_12_SFF_0_n9,
         md1FF_state_gff_12_SFF_0_n7, md1FF_state_gff_12_SFF_0_n6,
         md1FF_state_gff_12_SFF_1_n10, md1FF_state_gff_12_SFF_1_n9,
         md1FF_state_gff_12_SFF_1_n7, md1FF_state_gff_12_SFF_1_n6,
         md1FF_state_gff_12_SFF_2_n10, md1FF_state_gff_12_SFF_2_n9,
         md1FF_state_gff_12_SFF_2_n7, md1FF_state_gff_12_SFF_2_n6,
         md1FF_state_gff_12_SFF_3_n10, md1FF_state_gff_12_SFF_3_n9,
         md1FF_state_gff_12_SFF_3_n7, md1FF_state_gff_12_SFF_3_n6,
         md1FF_state_gff_13_SFF_0_n12, md1FF_state_gff_13_SFF_0_n11,
         md1FF_state_gff_13_SFF_0_n10, md1FF_state_gff_13_SFF_0_n8,
         md1FF_state_gff_13_SFF_0_n7, md1FF_state_gff_13_SFF_1_n12,
         md1FF_state_gff_13_SFF_1_n11, md1FF_state_gff_13_SFF_1_n10,
         md1FF_state_gff_13_SFF_1_n8, md1FF_state_gff_13_SFF_1_n7,
         md1FF_state_gff_13_SFF_2_n12, md1FF_state_gff_13_SFF_2_n11,
         md1FF_state_gff_13_SFF_2_n10, md1FF_state_gff_13_SFF_2_n8,
         md1FF_state_gff_13_SFF_2_n7, md1FF_state_gff_13_SFF_3_n12,
         md1FF_state_gff_13_SFF_3_n11, md1FF_state_gff_13_SFF_3_n10,
         md1FF_state_gff_13_SFF_3_n8, md1FF_state_gff_13_SFF_3_n7,
         md1FF_state_gff_14_SFF_0_n11, md1FF_state_gff_14_SFF_0_n10,
         md1FF_state_gff_14_SFF_0_n8, md1FF_state_gff_14_SFF_0_n7,
         md1FF_state_gff_14_SFF_1_n11, md1FF_state_gff_14_SFF_1_n10,
         md1FF_state_gff_14_SFF_1_n8, md1FF_state_gff_14_SFF_1_n7,
         md1FF_state_gff_14_SFF_2_n11, md1FF_state_gff_14_SFF_2_n10,
         md1FF_state_gff_14_SFF_2_n8, md1FF_state_gff_14_SFF_2_n7,
         md1FF_state_gff_14_SFF_3_n11, md1FF_state_gff_14_SFF_3_n10,
         md1FF_state_gff_14_SFF_3_n8, md1FF_state_gff_14_SFF_3_n7,
         md1FF_state_gff_15_SFF_0_n11, md1FF_state_gff_15_SFF_0_n10,
         md1FF_state_gff_15_SFF_0_n8, md1FF_state_gff_15_SFF_0_n7,
         md1FF_state_gff_15_SFF_1_n11, md1FF_state_gff_15_SFF_1_n10,
         md1FF_state_gff_15_SFF_1_n8, md1FF_state_gff_15_SFF_1_n7,
         md1FF_state_gff_15_SFF_2_n11, md1FF_state_gff_15_SFF_2_n10,
         md1FF_state_gff_15_SFF_2_n9, md1FF_state_gff_15_SFF_2_n7,
         md1FF_state_gff_15_SFF_2_n6, md1FF_state_gff_15_SFF_3_n11,
         md1FF_state_gff_15_SFF_3_n10, md1FF_state_gff_15_SFF_3_n9,
         md1FF_state_gff_15_SFF_3_n7, md1FF_state_gff_15_SFF_3_n6,
         md1FF_state_gff_16_n2, md1FF_state_gff_16_SFF_0_n10,
         md1FF_state_gff_16_SFF_0_n9, md1FF_state_gff_16_SFF_0_n7,
         md1FF_state_gff_16_SFF_0_n6, md1FF_state_gff_16_SFF_1_n10,
         md1FF_state_gff_16_SFF_1_n9, md1FF_state_gff_16_SFF_1_n7,
         md1FF_state_gff_16_SFF_1_n6, md1FF_state_gff_16_SFF_2_n10,
         md1FF_state_gff_16_SFF_2_n9, md1FF_state_gff_16_SFF_2_n7,
         md1FF_state_gff_16_SFF_2_n6, md1FF_state_gff_16_SFF_3_n9,
         md1FF_state_gff_16_SFF_3_n7, md1FF_state_gff_16_SFF_3_n6, keyFF_n4,
         keyFF_n3, keyFF_n2, keyFF_n1, keyFF_keystate_n18, keyFF_keystate_n17,
         keyFF_keystate_n16, keyFF_keystate_n15, keyFF_keystate_n14,
         keyFF_keystate_n13, keyFF_keystate_n12, keyFF_keystate_n11,
         keyFF_keystate_n10, keyFF_keystate_gff_1_SFF_0_n12,
         keyFF_keystate_gff_1_SFF_0_n11, keyFF_keystate_gff_1_SFF_0_n10,
         keyFF_keystate_gff_1_SFF_0_n8, keyFF_keystate_gff_1_SFF_0_n7,
         keyFF_keystate_gff_1_SFF_1_n12, keyFF_keystate_gff_1_SFF_1_n11,
         keyFF_keystate_gff_1_SFF_1_n10, keyFF_keystate_gff_1_SFF_1_n8,
         keyFF_keystate_gff_1_SFF_1_n7, keyFF_keystate_gff_1_SFF_2_n12,
         keyFF_keystate_gff_1_SFF_2_n11, keyFF_keystate_gff_1_SFF_2_n10,
         keyFF_keystate_gff_1_SFF_2_n8, keyFF_keystate_gff_1_SFF_2_n7,
         keyFF_keystate_gff_1_SFF_3_n12, keyFF_keystate_gff_1_SFF_3_n11,
         keyFF_keystate_gff_1_SFF_3_n10, keyFF_keystate_gff_1_SFF_3_n8,
         keyFF_keystate_gff_1_SFF_3_n7, keyFF_keystate_gff_2_SFF_0_n12,
         keyFF_keystate_gff_2_SFF_0_n11, keyFF_keystate_gff_2_SFF_0_n10,
         keyFF_keystate_gff_2_SFF_0_n8, keyFF_keystate_gff_2_SFF_0_n7,
         keyFF_keystate_gff_2_SFF_1_n12, keyFF_keystate_gff_2_SFF_1_n11,
         keyFF_keystate_gff_2_SFF_1_n10, keyFF_keystate_gff_2_SFF_1_n8,
         keyFF_keystate_gff_2_SFF_1_n7, keyFF_keystate_gff_2_SFF_2_n12,
         keyFF_keystate_gff_2_SFF_2_n11, keyFF_keystate_gff_2_SFF_2_n10,
         keyFF_keystate_gff_2_SFF_2_n8, keyFF_keystate_gff_2_SFF_2_n7,
         keyFF_keystate_gff_2_SFF_3_n12, keyFF_keystate_gff_2_SFF_3_n11,
         keyFF_keystate_gff_2_SFF_3_n10, keyFF_keystate_gff_2_SFF_3_n8,
         keyFF_keystate_gff_2_SFF_3_n7, keyFF_keystate_gff_3_SFF_0_n12,
         keyFF_keystate_gff_3_SFF_0_n11, keyFF_keystate_gff_3_SFF_0_n10,
         keyFF_keystate_gff_3_SFF_0_n8, keyFF_keystate_gff_3_SFF_0_n7,
         keyFF_keystate_gff_3_SFF_1_n12, keyFF_keystate_gff_3_SFF_1_n11,
         keyFF_keystate_gff_3_SFF_1_n10, keyFF_keystate_gff_3_SFF_1_n8,
         keyFF_keystate_gff_3_SFF_1_n7, keyFF_keystate_gff_3_SFF_2_n11,
         keyFF_keystate_gff_3_SFF_2_n10, keyFF_keystate_gff_3_SFF_2_n9,
         keyFF_keystate_gff_3_SFF_2_n7, keyFF_keystate_gff_3_SFF_2_n6,
         keyFF_keystate_gff_3_SFF_3_n11, keyFF_keystate_gff_3_SFF_3_n10,
         keyFF_keystate_gff_3_SFF_3_n9, keyFF_keystate_gff_3_SFF_3_n7,
         keyFF_keystate_gff_3_SFF_3_n6, keyFF_keystate_gff_4_SFF_0_n11,
         keyFF_keystate_gff_4_SFF_0_n10, keyFF_keystate_gff_4_SFF_0_n9,
         keyFF_keystate_gff_4_SFF_0_n7, keyFF_keystate_gff_4_SFF_0_n6,
         keyFF_keystate_gff_4_SFF_1_n11, keyFF_keystate_gff_4_SFF_1_n10,
         keyFF_keystate_gff_4_SFF_1_n9, keyFF_keystate_gff_4_SFF_1_n7,
         keyFF_keystate_gff_4_SFF_1_n6, keyFF_keystate_gff_4_SFF_2_n11,
         keyFF_keystate_gff_4_SFF_2_n10, keyFF_keystate_gff_4_SFF_2_n9,
         keyFF_keystate_gff_4_SFF_2_n7, keyFF_keystate_gff_4_SFF_2_n6,
         keyFF_keystate_gff_4_SFF_3_n11, keyFF_keystate_gff_4_SFF_3_n10,
         keyFF_keystate_gff_4_SFF_3_n9, keyFF_keystate_gff_4_SFF_3_n7,
         keyFF_keystate_gff_4_SFF_3_n6, keyFF_keystate_gff_5_SFF_0_n12,
         keyFF_keystate_gff_5_SFF_0_n11, keyFF_keystate_gff_5_SFF_0_n10,
         keyFF_keystate_gff_5_SFF_0_n8, keyFF_keystate_gff_5_SFF_0_n7,
         keyFF_keystate_gff_5_SFF_1_n12, keyFF_keystate_gff_5_SFF_1_n11,
         keyFF_keystate_gff_5_SFF_1_n10, keyFF_keystate_gff_5_SFF_1_n8,
         keyFF_keystate_gff_5_SFF_1_n7, keyFF_keystate_gff_5_SFF_2_n11,
         keyFF_keystate_gff_5_SFF_2_n10, keyFF_keystate_gff_5_SFF_2_n8,
         keyFF_keystate_gff_5_SFF_2_n7, keyFF_keystate_gff_5_SFF_3_n11,
         keyFF_keystate_gff_5_SFF_3_n10, keyFF_keystate_gff_5_SFF_3_n8,
         keyFF_keystate_gff_5_SFF_3_n7, keyFF_keystate_gff_6_SFF_0_n11,
         keyFF_keystate_gff_6_SFF_0_n10, keyFF_keystate_gff_6_SFF_0_n8,
         keyFF_keystate_gff_6_SFF_0_n7, keyFF_keystate_gff_6_SFF_1_n11,
         keyFF_keystate_gff_6_SFF_1_n10, keyFF_keystate_gff_6_SFF_1_n8,
         keyFF_keystate_gff_6_SFF_1_n7, keyFF_keystate_gff_6_SFF_2_n11,
         keyFF_keystate_gff_6_SFF_2_n10, keyFF_keystate_gff_6_SFF_2_n8,
         keyFF_keystate_gff_6_SFF_2_n7, keyFF_keystate_gff_6_SFF_3_n11,
         keyFF_keystate_gff_6_SFF_3_n10, keyFF_keystate_gff_6_SFF_3_n8,
         keyFF_keystate_gff_6_SFF_3_n7, keyFF_keystate_gff_7_SFF_0_n12,
         keyFF_keystate_gff_7_SFF_0_n11, keyFF_keystate_gff_7_SFF_0_n10,
         keyFF_keystate_gff_7_SFF_0_n8, keyFF_keystate_gff_7_SFF_0_n7,
         keyFF_keystate_gff_7_SFF_1_n12, keyFF_keystate_gff_7_SFF_1_n11,
         keyFF_keystate_gff_7_SFF_1_n10, keyFF_keystate_gff_7_SFF_1_n8,
         keyFF_keystate_gff_7_SFF_1_n7, keyFF_keystate_gff_7_SFF_2_n11,
         keyFF_keystate_gff_7_SFF_2_n10, keyFF_keystate_gff_7_SFF_2_n9,
         keyFF_keystate_gff_7_SFF_2_n7, keyFF_keystate_gff_7_SFF_2_n6,
         keyFF_keystate_gff_7_SFF_3_n11, keyFF_keystate_gff_7_SFF_3_n10,
         keyFF_keystate_gff_7_SFF_3_n9, keyFF_keystate_gff_7_SFF_3_n7,
         keyFF_keystate_gff_7_SFF_3_n6, keyFF_keystate_gff_8_SFF_0_n11,
         keyFF_keystate_gff_8_SFF_0_n10, keyFF_keystate_gff_8_SFF_0_n9,
         keyFF_keystate_gff_8_SFF_0_n7, keyFF_keystate_gff_8_SFF_0_n6,
         keyFF_keystate_gff_8_SFF_1_n11, keyFF_keystate_gff_8_SFF_1_n10,
         keyFF_keystate_gff_8_SFF_1_n9, keyFF_keystate_gff_8_SFF_1_n7,
         keyFF_keystate_gff_8_SFF_1_n6, keyFF_keystate_gff_8_SFF_2_n11,
         keyFF_keystate_gff_8_SFF_2_n10, keyFF_keystate_gff_8_SFF_2_n9,
         keyFF_keystate_gff_8_SFF_2_n7, keyFF_keystate_gff_8_SFF_2_n6,
         keyFF_keystate_gff_8_SFF_3_n11, keyFF_keystate_gff_8_SFF_3_n10,
         keyFF_keystate_gff_8_SFF_3_n9, keyFF_keystate_gff_8_SFF_3_n7,
         keyFF_keystate_gff_8_SFF_3_n6, keyFF_keystate_gff_9_SFF_0_n12,
         keyFF_keystate_gff_9_SFF_0_n11, keyFF_keystate_gff_9_SFF_0_n10,
         keyFF_keystate_gff_9_SFF_0_n8, keyFF_keystate_gff_9_SFF_0_n7,
         keyFF_keystate_gff_9_SFF_1_n12, keyFF_keystate_gff_9_SFF_1_n11,
         keyFF_keystate_gff_9_SFF_1_n10, keyFF_keystate_gff_9_SFF_1_n8,
         keyFF_keystate_gff_9_SFF_1_n7, keyFF_keystate_gff_9_SFF_2_n12,
         keyFF_keystate_gff_9_SFF_2_n11, keyFF_keystate_gff_9_SFF_2_n10,
         keyFF_keystate_gff_9_SFF_2_n8, keyFF_keystate_gff_9_SFF_2_n7,
         keyFF_keystate_gff_9_SFF_3_n12, keyFF_keystate_gff_9_SFF_3_n11,
         keyFF_keystate_gff_9_SFF_3_n10, keyFF_keystate_gff_9_SFF_3_n8,
         keyFF_keystate_gff_9_SFF_3_n7, keyFF_keystate_gff_10_SFF_0_n12,
         keyFF_keystate_gff_10_SFF_0_n11, keyFF_keystate_gff_10_SFF_0_n10,
         keyFF_keystate_gff_10_SFF_0_n8, keyFF_keystate_gff_10_SFF_0_n7,
         keyFF_keystate_gff_10_SFF_1_n12, keyFF_keystate_gff_10_SFF_1_n11,
         keyFF_keystate_gff_10_SFF_1_n10, keyFF_keystate_gff_10_SFF_1_n8,
         keyFF_keystate_gff_10_SFF_1_n7, keyFF_keystate_gff_10_SFF_2_n12,
         keyFF_keystate_gff_10_SFF_2_n11, keyFF_keystate_gff_10_SFF_2_n10,
         keyFF_keystate_gff_10_SFF_2_n8, keyFF_keystate_gff_10_SFF_2_n7,
         keyFF_keystate_gff_10_SFF_3_n12, keyFF_keystate_gff_10_SFF_3_n11,
         keyFF_keystate_gff_10_SFF_3_n10, keyFF_keystate_gff_10_SFF_3_n8,
         keyFF_keystate_gff_10_SFF_3_n7, keyFF_keystate_gff_11_SFF_0_n11,
         keyFF_keystate_gff_11_SFF_0_n10, keyFF_keystate_gff_11_SFF_0_n8,
         keyFF_keystate_gff_11_SFF_0_n7, keyFF_keystate_gff_11_SFF_1_n11,
         keyFF_keystate_gff_11_SFF_1_n10, keyFF_keystate_gff_11_SFF_1_n8,
         keyFF_keystate_gff_11_SFF_1_n7, keyFF_keystate_gff_11_SFF_2_n11,
         keyFF_keystate_gff_11_SFF_2_n10, keyFF_keystate_gff_11_SFF_2_n9,
         keyFF_keystate_gff_11_SFF_2_n7, keyFF_keystate_gff_11_SFF_2_n6,
         keyFF_keystate_gff_11_SFF_3_n11, keyFF_keystate_gff_11_SFF_3_n10,
         keyFF_keystate_gff_11_SFF_3_n9, keyFF_keystate_gff_11_SFF_3_n7,
         keyFF_keystate_gff_11_SFF_3_n6, keyFF_keystate_gff_12_SFF_0_n11,
         keyFF_keystate_gff_12_SFF_0_n10, keyFF_keystate_gff_12_SFF_0_n9,
         keyFF_keystate_gff_12_SFF_0_n7, keyFF_keystate_gff_12_SFF_0_n6,
         keyFF_keystate_gff_12_SFF_1_n11, keyFF_keystate_gff_12_SFF_1_n10,
         keyFF_keystate_gff_12_SFF_1_n9, keyFF_keystate_gff_12_SFF_1_n7,
         keyFF_keystate_gff_12_SFF_1_n6, keyFF_keystate_gff_12_SFF_2_n11,
         keyFF_keystate_gff_12_SFF_2_n10, keyFF_keystate_gff_12_SFF_2_n9,
         keyFF_keystate_gff_12_SFF_2_n7, keyFF_keystate_gff_12_SFF_2_n6,
         keyFF_keystate_gff_12_SFF_3_n11, keyFF_keystate_gff_12_SFF_3_n10,
         keyFF_keystate_gff_12_SFF_3_n9, keyFF_keystate_gff_12_SFF_3_n7,
         keyFF_keystate_gff_12_SFF_3_n6, keyFF_keystate_gff_13_SFF_0_n12,
         keyFF_keystate_gff_13_SFF_0_n11, keyFF_keystate_gff_13_SFF_0_n10,
         keyFF_keystate_gff_13_SFF_0_n8, keyFF_keystate_gff_13_SFF_0_n7,
         keyFF_keystate_gff_13_SFF_1_n12, keyFF_keystate_gff_13_SFF_1_n11,
         keyFF_keystate_gff_13_SFF_1_n10, keyFF_keystate_gff_13_SFF_1_n8,
         keyFF_keystate_gff_13_SFF_1_n7, keyFF_keystate_gff_13_SFF_2_n11,
         keyFF_keystate_gff_13_SFF_2_n10, keyFF_keystate_gff_13_SFF_2_n8,
         keyFF_keystate_gff_13_SFF_2_n7, keyFF_keystate_gff_13_SFF_3_n11,
         keyFF_keystate_gff_13_SFF_3_n10, keyFF_keystate_gff_13_SFF_3_n8,
         keyFF_keystate_gff_13_SFF_3_n7, keyFF_keystate_gff_14_SFF_0_n11,
         keyFF_keystate_gff_14_SFF_0_n10, keyFF_keystate_gff_14_SFF_0_n8,
         keyFF_keystate_gff_14_SFF_0_n7, keyFF_keystate_gff_14_SFF_1_n11,
         keyFF_keystate_gff_14_SFF_1_n10, keyFF_keystate_gff_14_SFF_1_n8,
         keyFF_keystate_gff_14_SFF_1_n7, keyFF_keystate_gff_14_SFF_2_n11,
         keyFF_keystate_gff_14_SFF_2_n10, keyFF_keystate_gff_14_SFF_2_n8,
         keyFF_keystate_gff_14_SFF_2_n7, keyFF_keystate_gff_14_SFF_3_n11,
         keyFF_keystate_gff_14_SFF_3_n10, keyFF_keystate_gff_14_SFF_3_n8,
         keyFF_keystate_gff_14_SFF_3_n7, keyFF_keystate_gff_15_SFF_0_n11,
         keyFF_keystate_gff_15_SFF_0_n10, keyFF_keystate_gff_15_SFF_0_n8,
         keyFF_keystate_gff_15_SFF_0_n7, keyFF_keystate_gff_15_SFF_1_n11,
         keyFF_keystate_gff_15_SFF_1_n10, keyFF_keystate_gff_15_SFF_1_n8,
         keyFF_keystate_gff_15_SFF_1_n7, keyFF_keystate_gff_15_SFF_2_n11,
         keyFF_keystate_gff_15_SFF_2_n10, keyFF_keystate_gff_15_SFF_2_n9,
         keyFF_keystate_gff_15_SFF_2_n7, keyFF_keystate_gff_15_SFF_2_n6,
         keyFF_keystate_gff_15_SFF_3_n11, keyFF_keystate_gff_15_SFF_3_n10,
         keyFF_keystate_gff_15_SFF_3_n9, keyFF_keystate_gff_15_SFF_3_n7,
         keyFF_keystate_gff_15_SFF_3_n6, keyFF_keystate_gff_16_SFF_0_n11,
         keyFF_keystate_gff_16_SFF_0_n10, keyFF_keystate_gff_16_SFF_0_n9,
         keyFF_keystate_gff_16_SFF_0_n7, keyFF_keystate_gff_16_SFF_0_n6,
         keyFF_keystate_gff_16_SFF_1_n11, keyFF_keystate_gff_16_SFF_1_n10,
         keyFF_keystate_gff_16_SFF_1_n9, keyFF_keystate_gff_16_SFF_1_n7,
         keyFF_keystate_gff_16_SFF_1_n6, keyFF_keystate_gff_16_SFF_2_n10,
         keyFF_keystate_gff_16_SFF_2_n9, keyFF_keystate_gff_16_SFF_2_n7,
         keyFF_keystate_gff_16_SFF_2_n6, keyFF_keystate_gff_16_SFF_3_n10,
         keyFF_keystate_gff_16_SFF_3_n9, keyFF_keystate_gff_16_SFF_3_n7,
         keyFF_keystate_gff_16_SFF_3_n6, keyFF_keystate_gff_17_SFF_0_n12,
         keyFF_keystate_gff_17_SFF_0_n11, keyFF_keystate_gff_17_SFF_0_n10,
         keyFF_keystate_gff_17_SFF_0_n8, keyFF_keystate_gff_17_SFF_0_n7,
         keyFF_keystate_gff_17_SFF_1_n12, keyFF_keystate_gff_17_SFF_1_n11,
         keyFF_keystate_gff_17_SFF_1_n10, keyFF_keystate_gff_17_SFF_1_n8,
         keyFF_keystate_gff_17_SFF_1_n7, keyFF_keystate_gff_17_SFF_2_n11,
         keyFF_keystate_gff_17_SFF_2_n10, keyFF_keystate_gff_17_SFF_2_n8,
         keyFF_keystate_gff_17_SFF_2_n7, keyFF_keystate_gff_17_SFF_3_n11,
         keyFF_keystate_gff_17_SFF_3_n10, keyFF_keystate_gff_17_SFF_3_n8,
         keyFF_keystate_gff_17_SFF_3_n7, keyFF_keystate_gff_18_SFF_0_n11,
         keyFF_keystate_gff_18_SFF_0_n10, keyFF_keystate_gff_18_SFF_0_n8,
         keyFF_keystate_gff_18_SFF_0_n7, keyFF_keystate_gff_18_SFF_1_n11,
         keyFF_keystate_gff_18_SFF_1_n10, keyFF_keystate_gff_18_SFF_1_n8,
         keyFF_keystate_gff_18_SFF_1_n7, keyFF_keystate_gff_18_SFF_2_n11,
         keyFF_keystate_gff_18_SFF_2_n10, keyFF_keystate_gff_18_SFF_2_n8,
         keyFF_keystate_gff_18_SFF_2_n7, keyFF_keystate_gff_18_SFF_3_n11,
         keyFF_keystate_gff_18_SFF_3_n10, keyFF_keystate_gff_18_SFF_3_n8,
         keyFF_keystate_gff_18_SFF_3_n7, keyFF_keystate_gff_19_SFF_0_n11,
         keyFF_keystate_gff_19_SFF_0_n10, keyFF_keystate_gff_19_SFF_0_n8,
         keyFF_keystate_gff_19_SFF_0_n7, keyFF_keystate_gff_19_SFF_1_n11,
         keyFF_keystate_gff_19_SFF_1_n10, keyFF_keystate_gff_19_SFF_1_n8,
         keyFF_keystate_gff_19_SFF_1_n7, keyFF_keystate_gff_19_SFF_2_n11,
         keyFF_keystate_gff_19_SFF_2_n10, keyFF_keystate_gff_19_SFF_2_n9,
         keyFF_keystate_gff_19_SFF_2_n7, keyFF_keystate_gff_19_SFF_2_n6,
         keyFF_keystate_gff_19_SFF_3_n11, keyFF_keystate_gff_19_SFF_3_n10,
         keyFF_keystate_gff_19_SFF_3_n9, keyFF_keystate_gff_19_SFF_3_n7,
         keyFF_keystate_gff_19_SFF_3_n6, keyFF_keystate_gff_20_SFF_0_n10,
         keyFF_keystate_gff_20_SFF_0_n9, keyFF_keystate_gff_20_SFF_0_n7,
         keyFF_keystate_gff_20_SFF_0_n6, keyFF_keystate_gff_20_SFF_1_n10,
         keyFF_keystate_gff_20_SFF_1_n9, keyFF_keystate_gff_20_SFF_1_n7,
         keyFF_keystate_gff_20_SFF_1_n6, keyFF_keystate_gff_20_SFF_2_n10,
         keyFF_keystate_gff_20_SFF_2_n9, keyFF_keystate_gff_20_SFF_2_n7,
         keyFF_keystate_gff_20_SFF_2_n6, keyFF_keystate_gff_20_SFF_3_n10,
         keyFF_keystate_gff_20_SFF_3_n9, keyFF_keystate_gff_20_SFF_3_n7,
         keyFF_keystate_gff_20_SFF_3_n6, sbox_Inst_N_F1_n10, sbox_Inst_N_F1_n9,
         sbox_Inst_N_F1_n8, sbox_Inst_N_F1_n7, sbox_Inst_N_F1_n6,
         sbox_Inst_N_F1_n5, sbox_Inst_N_F2_n9, sbox_Inst_N_F2_n8,
         sbox_Inst_N_F2_n7, sbox_Inst_N_F2_n6, sbox_Inst_N_F2_n5,
         sbox_Inst_N_F3_n10, sbox_Inst_N_F3_n9, sbox_Inst_N_F3_n8,
         sbox_Inst_N_F3_n7, sbox_Inst_N_F3_n6, sbox_Inst_N_F3_n5,
         sbox_Inst_N_F3_n4, sbox_Inst_N_F4_n13, sbox_Inst_N_F4_n12,
         sbox_Inst_N_F4_n11, sbox_Inst_N_F4_n10, sbox_Inst_N_F4_n9,
         sbox_Inst_N_F4_n8, sbox_Inst_N_F4_n7, sbox_Inst_N_F4_n6,
         sbox_Inst_N_F4_n5, sbox_Inst_N_F4_n4, sbox_Inst_N_F5_n11,
         sbox_Inst_N_F5_n10, sbox_Inst_N_F5_n9, sbox_Inst_N_F5_n8,
         sbox_Inst_N_F5_n7, sbox_Inst_N_F5_n6, sbox_Inst_N_F5_n5,
         sbox_Inst_N_F5_n4, sbox_Inst_N_F6_n9, sbox_Inst_N_F6_n8,
         sbox_Inst_N_F6_n7, sbox_Inst_N_F6_n6, sbox_Inst_N_F6_n5,
         sbox_Inst_N_F6_n4, sbox_Inst_N_F6_n3, sbox_Inst_N_F7_n6,
         sbox_Inst_N_F7_n5, sbox_Inst_N_F7_n4, sbox_Inst_N_F7_n3,
         sbox_Inst_N_F7_n2, sbox_Inst_N_F8_n8, sbox_Inst_N_F8_n7,
         sbox_Inst_N_F8_n6, sbox_Inst_N_F8_n5, sbox_Inst_N_F8_n4,
         sbox_Inst_N_F8_n3, sbox_Inst_L_XORInst1_n6, sbox_Inst_L_XORInst1_n5,
         sbox_Inst_L_XORInst2_n6, sbox_Inst_L_XORInst2_n5,
         sbox_Inst_L_XORInst5_n6, sbox_Inst_L_XORInst5_n5,
         sbox_Inst_L_XORInst6_n6, sbox_Inst_L_XORInst6_n5,
         sbox_Inst_L_XORInst7_n6, sbox_Inst_L_XORInst7_n5,
         sbox_Inst_L_XORInst8_n6, sbox_Inst_L_XORInst8_n5, sbox_KS_n18,
         sbox_KS_n17, sbox_KS_n16, sbox_KS_n15, sbox_KS_n14, sbox_KS_n13,
         sbox_KS_n12, sbox_KS_n11, sbox_KS_n10, sbox_KS_n9, sbox_KS_n8,
         sbox_KS_n7, sbox_KS_n6, sbox_KS_n5;
  wire   [4:0] counter;
  wire   [3:0] share1;
  wire   [3:0] state;
  wire   [3:0] share2;
  wire   [3:0] sboxKS;
  wire   [3:0] roundkey;
  wire   [3:1] keyRegKS;
  wire   [3:0] fsm_countSerial;
  wire   [62:1] stateFF_inputPar;
  wire   [6:48] stateFF_n;
  wire   [62:1] md1FF_inputPar;
  wire   [14:56] md1FF_n;
  wire   [4:0] keyFF_counterAdd;
  wire   [75:3] keyFF_outputPar;
  wire   [8:1] sbox_h_reg;
  wire   [8:1] sbox_g_reg;
  wire   [4:1] sbox_e_reg;
  wire   [8:1] sbox_f_reg;
  wire   [8:1] sbox_h;
  wire   [8:1] sbox_g;
  wire   [8:1] sbox_f;
  wire   [4:1] sbox_e;

  XOR2_X2 U9 ( .A(roundkey[3]), .B(state[3]), .Z(dataOut1[3]) );
  XOR2_X2 U10 ( .A(roundkey[2]), .B(state[2]), .Z(dataOut1[2]) );
  XOR2_X1 U11 ( .A(roundkey[0]), .B(state[0]), .Z(dataOut1[0]) );
  XOR2_X2 U12 ( .A(roundkey[1]), .B(state[1]), .Z(dataOut1[1]) );
  OAI211_X1 fsm_U19 ( .C1(fsm_n7), .C2(fsm_n20), .A(enKey), .B(nReset), .ZN(
        fsm_n21) );
  AOI221_X1 fsm_U18 ( .B1(fsm_n19), .B2(fsm_n18), .C1(fsm_n20), .C2(fsm_n18), 
        .A(fsm_n15), .ZN(fsm_n17) );
  NAND3_X1 fsm_U17 ( .A1(fsm_ps_state_2_), .A2(fsm_n9), .A3(fsm_n7), .ZN(
        fsm_n18) );
  AOI21_X1 fsm_U16 ( .B1(fsm_n14), .B2(fsm_n12), .A(fsm_n15), .ZN(fsm_n16) );
  INV_X1 fsm_U15 ( .A(nReset), .ZN(fsm_n15) );
  NAND3_X1 fsm_U14 ( .A1(selP), .A2(counter[3]), .A3(fsm_n11), .ZN(fsm_n12) );
  AND4_X1 fsm_U13 ( .A1(counter[4]), .A2(counter[1]), .A3(counter[0]), .A4(
        counter[2]), .ZN(fsm_n11) );
  AOI21_X1 fsm_U12 ( .B1(done), .B2(fsm_n20), .A(fsm_en_countRound), .ZN(
        fsm_n14) );
  NOR3_X1 fsm_U11 ( .A1(fsm_ps_state_1_), .A2(fsm_n20), .A3(fsm_n10), .ZN(
        fsm_en_countRound) );
  NAND4_X1 fsm_U10 ( .A1(fsm_countSerial[2]), .A2(fsm_countSerial[3]), .A3(
        fsm_countSerial[0]), .A4(fsm_countSerial[1]), .ZN(fsm_n20) );
  INV_X1 fsm_U9 ( .A(fsm_n19), .ZN(done) );
  NAND2_X1 fsm_U8 ( .A1(fsm_ps_state_1_), .A2(fsm_n13), .ZN(fsm_n19) );
  INV_X1 fsm_U7 ( .A(fsm_n10), .ZN(fsm_n13) );
  NAND2_X1 fsm_U6 ( .A1(enKey), .A2(fsm_ps_state_0_), .ZN(fsm_n10) );
  NAND2_X1 fsm_U5 ( .A1(fsm_n7), .A2(enKey), .ZN(fsm_rst_countSerial) );
  NOR2_X1 fsm_U4 ( .A1(fsm_n9), .A2(fsm_rst_countSerial), .ZN(selP) );
  NOR2_X2 fsm_U3 ( .A1(fsm_rst_countSerial), .A2(fsm_ps_state_1_), .ZN(selInit) );
  DFF_X1 fsm_ps_state_reg_0_ ( .D(fsm_n21), .CK(clk), .Q(fsm_n7), .QN(
        fsm_ps_state_0_) );
  DFF_X1 fsm_ps_state_reg_1_ ( .D(fsm_n16), .CK(clk), .Q(fsm_ps_state_1_), 
        .QN(fsm_n9) );
  DFF_X1 fsm_ps_state_reg_2_ ( .D(fsm_n17), .CK(clk), .Q(fsm_ps_state_2_), 
        .QN(enKey) );
  AOI22_X1 fsm_cnt_rnd_U23 ( .A1(counter[0]), .A2(fsm_cnt_rnd_n40), .B1(
        fsm_cnt_rnd_n39), .B2(fsm_cnt_rnd_n27), .ZN(fsm_cnt_rnd_n5) );
  OR2_X1 fsm_cnt_rnd_U22 ( .A1(selInit), .A2(fsm_en_countRound), .ZN(
        fsm_cnt_rnd_n40) );
  OAI21_X1 fsm_cnt_rnd_U21 ( .B1(fsm_cnt_rnd_n38), .B2(counter[4]), .A(
        fsm_cnt_rnd_n37), .ZN(fsm_cnt_rnd_n20) );
  OAI21_X1 fsm_cnt_rnd_U20 ( .B1(fsm_cnt_rnd_n36), .B2(fsm_cnt_rnd_n35), .A(
        counter[4]), .ZN(fsm_cnt_rnd_n37) );
  NAND3_X1 fsm_cnt_rnd_U19 ( .A1(fsm_cnt_rnd_n34), .A2(counter[3]), .A3(
        fsm_cnt_rnd_n33), .ZN(fsm_cnt_rnd_n38) );
  INV_X1 fsm_cnt_rnd_U18 ( .A(fsm_cnt_rnd_n32), .ZN(fsm_cnt_rnd_n21) );
  AOI22_X1 fsm_cnt_rnd_U17 ( .A1(counter[3]), .A2(fsm_cnt_rnd_n36), .B1(
        fsm_cnt_rnd_n35), .B2(fsm_cnt_rnd_n33), .ZN(fsm_cnt_rnd_n32) );
  NOR2_X1 fsm_cnt_rnd_U16 ( .A1(counter[3]), .A2(fsm_cnt_rnd_n39), .ZN(
        fsm_cnt_rnd_n35) );
  AOI21_X1 fsm_cnt_rnd_U15 ( .B1(fsm_en_countRound), .B2(fsm_cnt_rnd_n33), .A(
        selInit), .ZN(fsm_cnt_rnd_n36) );
  NOR3_X1 fsm_cnt_rnd_U14 ( .A1(fsm_cnt_rnd_n27), .A2(fsm_cnt_rnd_n28), .A3(
        fsm_cnt_rnd_n26), .ZN(fsm_cnt_rnd_n33) );
  AOI22_X1 fsm_cnt_rnd_U13 ( .A1(counter[1]), .A2(fsm_cnt_rnd_n29), .B1(
        fsm_cnt_rnd_n31), .B2(fsm_cnt_rnd_n26), .ZN(fsm_cnt_rnd_n23) );
  NAND2_X1 fsm_cnt_rnd_U12 ( .A1(fsm_cnt_rnd_n34), .A2(counter[0]), .ZN(
        fsm_cnt_rnd_n31) );
  INV_X1 fsm_cnt_rnd_U11 ( .A(fsm_cnt_rnd_n39), .ZN(fsm_cnt_rnd_n34) );
  INV_X1 fsm_cnt_rnd_U10 ( .A(fsm_cnt_rnd_n30), .ZN(fsm_cnt_rnd_n29) );
  AOI21_X1 fsm_cnt_rnd_U9 ( .B1(fsm_en_countRound), .B2(counter[0]), .A(
        selInit), .ZN(fsm_cnt_rnd_n30) );
  INV_X1 fsm_cnt_rnd_U7 ( .A(fsm_cnt_rnd_n28), .ZN(fsm_cnt_rnd_n24) );
  AOI21_X1 fsm_cnt_rnd_U6 ( .B1(fsm_cnt_rnd_n26), .B2(fsm_cnt_rnd_n34), .A(
        fsm_cnt_rnd_n30), .ZN(fsm_cnt_rnd_n19) );
  NAND2_X1 fsm_cnt_rnd_U5 ( .A1(fsm_en_countRound), .A2(fsm_cnt_rnd_n18), .ZN(
        fsm_cnt_rnd_n39) );
  INV_X1 fsm_cnt_rnd_U4 ( .A(selInit), .ZN(fsm_cnt_rnd_n18) );
  OAI33_X1 fsm_cnt_rnd_U3 ( .A1(1'b0), .A2(fsm_cnt_rnd_n28), .A3(
        fsm_cnt_rnd_n19), .B1(fsm_cnt_rnd_n24), .B2(fsm_cnt_rnd_n26), .B3(
        fsm_cnt_rnd_n31), .ZN(fsm_cnt_rnd_n22) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_0_ ( .D(fsm_cnt_rnd_n5), .CK(clk), .Q(
        counter[0]), .QN(fsm_cnt_rnd_n27) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_1_ ( .D(fsm_cnt_rnd_n23), .CK(clk), .Q(
        counter[1]), .QN(fsm_cnt_rnd_n26) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_2_ ( .D(fsm_cnt_rnd_n22), .CK(clk), .Q(
        counter[2]), .QN(fsm_cnt_rnd_n28) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_3_ ( .D(fsm_cnt_rnd_n21), .CK(clk), .Q(
        counter[3]), .QN() );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_4_ ( .D(fsm_cnt_rnd_n20), .CK(clk), .Q(
        counter[4]), .QN() );
  INV_X1 fsm_cnt_ser_U13 ( .A(fsm_cnt_ser_n21), .ZN(fsm_cnt_ser_n20) );
  OAI211_X1 fsm_cnt_ser_U12 ( .C1(fsm_n13), .C2(fsm_countSerial[0]), .A(
        fsm_rst_countSerial), .B(fsm_cnt_ser_n16), .ZN(fsm_cnt_ser_n21) );
  AOI211_X1 fsm_cnt_ser_U11 ( .C1(fsm_cnt_ser_n16), .C2(fsm_cnt_ser_n10), .A(
        fsm_cnt_ser_n15), .B(fsm_cnt_ser_n14), .ZN(fsm_cnt_ser_n19) );
  INV_X1 fsm_cnt_ser_U10 ( .A(fsm_cnt_ser_n13), .ZN(fsm_cnt_ser_n15) );
  NAND2_X1 fsm_cnt_ser_U9 ( .A1(fsm_n13), .A2(fsm_countSerial[0]), .ZN(
        fsm_cnt_ser_n16) );
  AOI211_X1 fsm_cnt_ser_U8 ( .C1(fsm_cnt_ser_n13), .C2(fsm_cnt_ser_n9), .A(
        fsm_cnt_ser_n12), .B(fsm_cnt_ser_n14), .ZN(fsm_cnt_ser_n18) );
  INV_X1 fsm_cnt_ser_U7 ( .A(fsm_rst_countSerial), .ZN(fsm_cnt_ser_n14) );
  AOI21_X1 fsm_cnt_ser_U6 ( .B1(fsm_cnt_ser_n12), .B2(fsm_countSerial[3]), .A(
        fsm_cnt_ser_n11), .ZN(fsm_cnt_ser_n17) );
  OAI21_X1 fsm_cnt_ser_U5 ( .B1(fsm_cnt_ser_n12), .B2(fsm_countSerial[3]), .A(
        fsm_rst_countSerial), .ZN(fsm_cnt_ser_n11) );
  NOR2_X1 fsm_cnt_ser_U4 ( .A1(fsm_cnt_ser_n13), .A2(fsm_cnt_ser_n9), .ZN(
        fsm_cnt_ser_n12) );
  NAND3_X1 fsm_cnt_ser_U3 ( .A1(fsm_n13), .A2(fsm_countSerial[0]), .A3(
        fsm_countSerial[1]), .ZN(fsm_cnt_ser_n13) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_3_ ( .D(fsm_cnt_ser_n17), .CK(clk), .Q(
        fsm_countSerial[3]), .QN() );
  DFF_X1 fsm_cnt_ser_count_reg_reg_2_ ( .D(fsm_cnt_ser_n18), .CK(clk), .Q(
        fsm_countSerial[2]), .QN(fsm_cnt_ser_n9) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_1_ ( .D(fsm_cnt_ser_n19), .CK(clk), .Q(
        fsm_countSerial[1]), .QN(fsm_cnt_ser_n10) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_0_ ( .D(fsm_cnt_ser_n20), .CK(clk), .Q(
        fsm_countSerial[0]), .QN() );
  MUX2_X1 stateFF_U5 ( .A(share1[0]), .B(dataIn1[0]), .S(selInit), .Z(
        stateFF_n1) );
  MUX2_X1 stateFF_U4 ( .A(share1[2]), .B(dataIn1[2]), .S(selInit), .Z(
        stateFF_inputPar[32]) );
  MUX2_X1 stateFF_U3 ( .A(share1[1]), .B(dataIn1[1]), .S(selInit), .Z(
        stateFF_inputPar[16]) );
  MUX2_X1 stateFF_U2 ( .A(share1[3]), .B(dataIn1[3]), .S(selInit), .Z(
        stateFF_inputPar[48]) );
  BUF_X1 stateFF_state_U6 ( .A(selP), .Z(stateFF_state_n9) );
  BUF_X1 stateFF_state_U5 ( .A(selP), .Z(stateFF_state_n10) );
  BUF_X1 stateFF_state_U4 ( .A(selP), .Z(stateFF_state_n11) );
  BUF_X2 stateFF_state_U3 ( .A(enKey), .Z(stateFF_state_n6) );
  BUF_X2 stateFF_state_U2 ( .A(enKey), .Z(stateFF_state_n8) );
  BUF_X2 stateFF_state_U1 ( .A(enKey), .Z(stateFF_state_n7) );
  BUF_X1 stateFF_state_gff_1_U2 ( .A(stateFF_state_n10), .Z(
        stateFF_state_gff_1_n2) );
  OAI21_X1 stateFF_state_gff_1_SFF_0_U3 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_1_SFF_0_n7), .A(stateFF_state_gff_1_SFF_0_n9), .ZN(
        stateFF_state_gff_1_SFF_0_n6) );
  NAND2_X1 stateFF_state_gff_1_SFF_0_U2 ( .A1(stateFF_state_n7), .A2(
        stateFF_n1), .ZN(stateFF_state_gff_1_SFF_0_n9) );
  DFF_X1 stateFF_state_gff_1_SFF_0_Cell_reg ( .D(stateFF_state_gff_1_SFF_0_n6), 
        .CK(clk), .Q(stateFF_inputPar[1]), .QN(stateFF_state_gff_1_SFF_0_n7)
         );
  OAI21_X1 stateFF_state_gff_1_SFF_1_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_1_SFF_1_n8), .A(stateFF_state_gff_1_SFF_1_n11), .ZN(
        stateFF_state_gff_1_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_1_SFF_1_U3 ( .B1(stateFF_state_gff_1_n2), .B2(
        stateFF_inputPar[16]), .C1(stateFF_state_gff_1_SFF_1_n10), .C2(
        stateFF_inputPar[1]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_1_SFF_1_n11) );
  INV_X1 stateFF_state_gff_1_SFF_1_U2 ( .A(stateFF_state_gff_1_n2), .ZN(
        stateFF_state_gff_1_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_1_SFF_1_Cell_reg ( .D(stateFF_state_gff_1_SFF_1_n7), 
        .CK(clk), .Q(stateFF_inputPar[17]), .QN(stateFF_state_gff_1_SFF_1_n8)
         );
  OAI21_X1 stateFF_state_gff_1_SFF_2_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_1_SFF_2_n8), .A(stateFF_state_gff_1_SFF_2_n11), .ZN(
        stateFF_state_gff_1_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_1_SFF_2_U3 ( .B1(stateFF_state_gff_1_n2), .B2(
        stateFF_inputPar[32]), .C1(stateFF_state_gff_1_SFF_2_n10), .C2(
        stateFF_inputPar[2]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_1_SFF_2_n11) );
  INV_X1 stateFF_state_gff_1_SFF_2_U2 ( .A(stateFF_state_gff_1_n2), .ZN(
        stateFF_state_gff_1_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_1_SFF_2_Cell_reg ( .D(stateFF_state_gff_1_SFF_2_n7), 
        .CK(clk), .Q(stateFF_inputPar[33]), .QN(stateFF_state_gff_1_SFF_2_n8)
         );
  OAI21_X1 stateFF_state_gff_1_SFF_3_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_1_SFF_3_n8), .A(stateFF_state_gff_1_SFF_3_n11), .ZN(
        stateFF_state_gff_1_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_1_SFF_3_U3 ( .B1(stateFF_state_gff_1_n2), .B2(
        stateFF_inputPar[48]), .C1(stateFF_state_gff_1_SFF_3_n10), .C2(
        stateFF_inputPar[3]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_1_SFF_3_n11) );
  INV_X1 stateFF_state_gff_1_SFF_3_U2 ( .A(stateFF_state_gff_1_n2), .ZN(
        stateFF_state_gff_1_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_1_SFF_3_Cell_reg ( .D(stateFF_state_gff_1_SFF_3_n7), 
        .CK(clk), .Q(stateFF_inputPar[49]), .QN(stateFF_state_gff_1_SFF_3_n8)
         );
  OAI21_X1 stateFF_state_gff_2_SFF_0_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_2_SFF_0_n8), .A(stateFF_state_gff_2_SFF_0_n12), .ZN(
        stateFF_state_gff_2_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_2_SFF_0_U4 ( .B1(stateFF_state_gff_2_SFF_0_n10), 
        .B2(stateFF_inputPar[1]), .C1(stateFF_state_gff_2_SFF_0_n11), .C2(
        stateFF_inputPar[4]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_2_SFF_0_n12) );
  INV_X1 stateFF_state_gff_2_SFF_0_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_2_SFF_0_n11) );
  INV_X1 stateFF_state_gff_2_SFF_0_U2 ( .A(stateFF_state_gff_2_SFF_0_n11), 
        .ZN(stateFF_state_gff_2_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_2_SFF_0_Cell_reg ( .D(stateFF_state_gff_2_SFF_0_n7), 
        .CK(clk), .Q(stateFF_inputPar[2]), .QN(stateFF_state_gff_2_SFF_0_n8)
         );
  OAI21_X1 stateFF_state_gff_2_SFF_1_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_2_SFF_1_n8), .A(stateFF_state_gff_2_SFF_1_n12), .ZN(
        stateFF_state_gff_2_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_2_SFF_1_U4 ( .B1(stateFF_state_gff_2_SFF_1_n10), 
        .B2(stateFF_inputPar[17]), .C1(stateFF_state_gff_2_SFF_1_n11), .C2(
        stateFF_inputPar[5]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_2_SFF_1_n12) );
  INV_X1 stateFF_state_gff_2_SFF_1_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_2_SFF_1_n11) );
  INV_X1 stateFF_state_gff_2_SFF_1_U2 ( .A(stateFF_state_gff_2_SFF_1_n11), 
        .ZN(stateFF_state_gff_2_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_2_SFF_1_Cell_reg ( .D(stateFF_state_gff_2_SFF_1_n7), 
        .CK(clk), .Q(stateFF_inputPar[18]), .QN(stateFF_state_gff_2_SFF_1_n8)
         );
  OAI21_X1 stateFF_state_gff_2_SFF_2_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_2_SFF_2_n8), .A(stateFF_state_gff_2_SFF_2_n12), .ZN(
        stateFF_state_gff_2_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_2_SFF_2_U4 ( .B1(stateFF_state_gff_2_SFF_2_n10), 
        .B2(stateFF_inputPar[33]), .C1(stateFF_state_gff_2_SFF_2_n11), .C2(
        stateFF_inputPar[6]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_2_SFF_2_n12) );
  INV_X1 stateFF_state_gff_2_SFF_2_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_2_SFF_2_n11) );
  INV_X1 stateFF_state_gff_2_SFF_2_U2 ( .A(stateFF_state_gff_2_SFF_2_n11), 
        .ZN(stateFF_state_gff_2_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_2_SFF_2_Cell_reg ( .D(stateFF_state_gff_2_SFF_2_n7), 
        .CK(clk), .Q(stateFF_inputPar[34]), .QN(stateFF_state_gff_2_SFF_2_n8)
         );
  OAI21_X1 stateFF_state_gff_2_SFF_3_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_2_SFF_3_n8), .A(stateFF_state_gff_2_SFF_3_n12), .ZN(
        stateFF_state_gff_2_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_2_SFF_3_U4 ( .B1(stateFF_state_gff_2_SFF_3_n10), 
        .B2(stateFF_inputPar[49]), .C1(stateFF_state_gff_2_SFF_3_n11), .C2(
        stateFF_inputPar[7]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_2_SFF_3_n12) );
  INV_X1 stateFF_state_gff_2_SFF_3_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_2_SFF_3_n11) );
  INV_X1 stateFF_state_gff_2_SFF_3_U2 ( .A(stateFF_state_gff_2_SFF_3_n11), 
        .ZN(stateFF_state_gff_2_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_2_SFF_3_Cell_reg ( .D(stateFF_state_gff_2_SFF_3_n7), 
        .CK(clk), .Q(stateFF_inputPar[50]), .QN(stateFF_state_gff_2_SFF_3_n8)
         );
  OAI21_X1 stateFF_state_gff_3_SFF_0_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_3_SFF_0_n8), .A(stateFF_state_gff_3_SFF_0_n11), .ZN(
        stateFF_state_gff_3_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_3_SFF_0_U3 ( .B1(stateFF_state_n9), .B2(
        stateFF_inputPar[2]), .C1(stateFF_state_gff_3_SFF_0_n10), .C2(
        stateFF_inputPar[8]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_3_SFF_0_n11) );
  INV_X1 stateFF_state_gff_3_SFF_0_U2 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_3_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_3_SFF_0_Cell_reg ( .D(stateFF_state_gff_3_SFF_0_n7), 
        .CK(clk), .Q(stateFF_inputPar[3]), .QN(stateFF_state_gff_3_SFF_0_n8)
         );
  OAI21_X1 stateFF_state_gff_3_SFF_1_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_3_SFF_1_n8), .A(stateFF_state_gff_3_SFF_1_n11), .ZN(
        stateFF_state_gff_3_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_3_SFF_1_U3 ( .B1(stateFF_state_n9), .B2(
        stateFF_inputPar[18]), .C1(stateFF_state_gff_3_SFF_1_n10), .C2(
        stateFF_inputPar[9]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_3_SFF_1_n11) );
  INV_X1 stateFF_state_gff_3_SFF_1_U2 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_3_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_3_SFF_1_Cell_reg ( .D(stateFF_state_gff_3_SFF_1_n7), 
        .CK(clk), .Q(stateFF_inputPar[19]), .QN(stateFF_state_gff_3_SFF_1_n8)
         );
  OAI21_X1 stateFF_state_gff_3_SFF_2_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_3_SFF_2_n8), .A(stateFF_state_gff_3_SFF_2_n11), .ZN(
        stateFF_state_gff_3_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_3_SFF_2_U3 ( .B1(stateFF_state_n9), .B2(
        stateFF_inputPar[34]), .C1(stateFF_state_gff_3_SFF_2_n10), .C2(
        stateFF_inputPar[10]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_3_SFF_2_n11) );
  INV_X1 stateFF_state_gff_3_SFF_2_U2 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_3_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_3_SFF_2_Cell_reg ( .D(stateFF_state_gff_3_SFF_2_n7), 
        .CK(clk), .Q(stateFF_inputPar[35]), .QN(stateFF_state_gff_3_SFF_2_n8)
         );
  OAI21_X1 stateFF_state_gff_3_SFF_3_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_3_SFF_3_n8), .A(stateFF_state_gff_3_SFF_3_n11), .ZN(
        stateFF_state_gff_3_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_3_SFF_3_U3 ( .B1(stateFF_state_n9), .B2(
        stateFF_inputPar[50]), .C1(stateFF_state_gff_3_SFF_3_n10), .C2(
        stateFF_inputPar[11]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_3_SFF_3_n11) );
  INV_X1 stateFF_state_gff_3_SFF_3_U2 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_3_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_3_SFF_3_Cell_reg ( .D(stateFF_state_gff_3_SFF_3_n7), 
        .CK(clk), .Q(stateFF_inputPar[51]), .QN(stateFF_state_gff_3_SFF_3_n8)
         );
  OAI21_X1 stateFF_state_gff_4_SFF_0_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_4_SFF_0_n8), .A(stateFF_state_gff_4_SFF_0_n11), .ZN(
        stateFF_state_gff_4_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_4_SFF_0_U3 ( .B1(stateFF_state_n9), .B2(
        stateFF_inputPar[3]), .C1(stateFF_state_gff_4_SFF_0_n10), .C2(
        stateFF_inputPar[12]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_4_SFF_0_n11) );
  INV_X1 stateFF_state_gff_4_SFF_0_U2 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_4_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_4_SFF_0_Cell_reg ( .D(stateFF_state_gff_4_SFF_0_n7), 
        .CK(clk), .Q(stateFF_inputPar[4]), .QN(stateFF_state_gff_4_SFF_0_n8)
         );
  OAI21_X1 stateFF_state_gff_4_SFF_1_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_4_SFF_1_n8), .A(stateFF_state_gff_4_SFF_1_n11), .ZN(
        stateFF_state_gff_4_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_4_SFF_1_U3 ( .B1(stateFF_state_n9), .B2(
        stateFF_inputPar[19]), .C1(stateFF_state_gff_4_SFF_1_n10), .C2(
        stateFF_inputPar[13]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_4_SFF_1_n11) );
  INV_X1 stateFF_state_gff_4_SFF_1_U2 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_4_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_4_SFF_1_Cell_reg ( .D(stateFF_state_gff_4_SFF_1_n7), 
        .CK(clk), .Q(stateFF_inputPar[20]), .QN(stateFF_state_gff_4_SFF_1_n8)
         );
  OAI21_X1 stateFF_state_gff_4_SFF_2_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_4_SFF_2_n7), .A(stateFF_state_gff_4_SFF_2_n11), .ZN(
        stateFF_state_gff_4_SFF_2_n6) );
  OAI221_X1 stateFF_state_gff_4_SFF_2_U4 ( .B1(stateFF_state_gff_4_SFF_2_n9), 
        .B2(stateFF_inputPar[35]), .C1(stateFF_state_gff_4_SFF_2_n10), .C2(
        stateFF_inputPar[14]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_4_SFF_2_n11) );
  INV_X1 stateFF_state_gff_4_SFF_2_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_4_SFF_2_n10) );
  INV_X1 stateFF_state_gff_4_SFF_2_U2 ( .A(stateFF_state_gff_4_SFF_2_n10), 
        .ZN(stateFF_state_gff_4_SFF_2_n9) );
  DFF_X1 stateFF_state_gff_4_SFF_2_Cell_reg ( .D(stateFF_state_gff_4_SFF_2_n6), 
        .CK(clk), .Q(stateFF_inputPar[36]), .QN(stateFF_state_gff_4_SFF_2_n7)
         );
  OAI21_X1 stateFF_state_gff_4_SFF_3_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_4_SFF_3_n7), .A(stateFF_state_gff_4_SFF_3_n11), .ZN(
        stateFF_state_gff_4_SFF_3_n6) );
  OAI221_X1 stateFF_state_gff_4_SFF_3_U4 ( .B1(stateFF_state_gff_4_SFF_3_n9), 
        .B2(stateFF_inputPar[51]), .C1(stateFF_state_gff_4_SFF_3_n10), .C2(
        stateFF_inputPar[15]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_4_SFF_3_n11) );
  INV_X1 stateFF_state_gff_4_SFF_3_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_4_SFF_3_n10) );
  INV_X1 stateFF_state_gff_4_SFF_3_U2 ( .A(stateFF_state_gff_4_SFF_3_n10), 
        .ZN(stateFF_state_gff_4_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_4_SFF_3_Cell_reg ( .D(stateFF_state_gff_4_SFF_3_n6), 
        .CK(clk), .Q(stateFF_inputPar[52]), .QN(stateFF_state_gff_4_SFF_3_n7)
         );
  OAI21_X1 stateFF_state_gff_5_SFF_0_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_5_SFF_0_n7), .A(stateFF_state_gff_5_SFF_0_n11), .ZN(
        stateFF_state_gff_5_SFF_0_n6) );
  OAI221_X1 stateFF_state_gff_5_SFF_0_U4 ( .B1(stateFF_state_gff_5_SFF_0_n9), 
        .B2(stateFF_inputPar[4]), .C1(stateFF_state_gff_5_SFF_0_n10), .C2(
        stateFF_inputPar[16]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_5_SFF_0_n11) );
  INV_X1 stateFF_state_gff_5_SFF_0_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_5_SFF_0_n10) );
  INV_X1 stateFF_state_gff_5_SFF_0_U2 ( .A(stateFF_state_gff_5_SFF_0_n10), 
        .ZN(stateFF_state_gff_5_SFF_0_n9) );
  DFF_X1 stateFF_state_gff_5_SFF_0_Cell_reg ( .D(stateFF_state_gff_5_SFF_0_n6), 
        .CK(clk), .Q(stateFF_inputPar[5]), .QN(stateFF_state_gff_5_SFF_0_n7)
         );
  OAI21_X1 stateFF_state_gff_5_SFF_1_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_5_SFF_1_n7), .A(stateFF_state_gff_5_SFF_1_n11), .ZN(
        stateFF_state_gff_5_SFF_1_n6) );
  OAI221_X1 stateFF_state_gff_5_SFF_1_U4 ( .B1(stateFF_state_gff_5_SFF_1_n9), 
        .B2(stateFF_inputPar[20]), .C1(stateFF_state_gff_5_SFF_1_n10), .C2(
        stateFF_inputPar[17]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_5_SFF_1_n11) );
  INV_X1 stateFF_state_gff_5_SFF_1_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_5_SFF_1_n10) );
  INV_X1 stateFF_state_gff_5_SFF_1_U2 ( .A(stateFF_state_gff_5_SFF_1_n10), 
        .ZN(stateFF_state_gff_5_SFF_1_n9) );
  DFF_X1 stateFF_state_gff_5_SFF_1_Cell_reg ( .D(stateFF_state_gff_5_SFF_1_n6), 
        .CK(clk), .Q(stateFF_n[48]), .QN(stateFF_state_gff_5_SFF_1_n7) );
  OAI21_X1 stateFF_state_gff_5_SFF_2_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_5_SFF_2_n7), .A(stateFF_state_gff_5_SFF_2_n11), .ZN(
        stateFF_state_gff_5_SFF_2_n6) );
  OAI221_X1 stateFF_state_gff_5_SFF_2_U4 ( .B1(stateFF_state_gff_5_SFF_2_n9), 
        .B2(stateFF_inputPar[36]), .C1(stateFF_state_gff_5_SFF_2_n10), .C2(
        stateFF_inputPar[18]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_5_SFF_2_n11) );
  INV_X1 stateFF_state_gff_5_SFF_2_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_5_SFF_2_n10) );
  INV_X1 stateFF_state_gff_5_SFF_2_U2 ( .A(stateFF_state_gff_5_SFF_2_n10), 
        .ZN(stateFF_state_gff_5_SFF_2_n9) );
  DFF_X1 stateFF_state_gff_5_SFF_2_Cell_reg ( .D(stateFF_state_gff_5_SFF_2_n6), 
        .CK(clk), .Q(stateFF_inputPar[37]), .QN(stateFF_state_gff_5_SFF_2_n7)
         );
  OAI21_X1 stateFF_state_gff_5_SFF_3_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_5_SFF_3_n7), .A(stateFF_state_gff_5_SFF_3_n11), .ZN(
        stateFF_state_gff_5_SFF_3_n6) );
  OAI221_X1 stateFF_state_gff_5_SFF_3_U4 ( .B1(stateFF_state_gff_5_SFF_3_n9), 
        .B2(stateFF_inputPar[52]), .C1(stateFF_state_gff_5_SFF_3_n10), .C2(
        stateFF_inputPar[19]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_5_SFF_3_n11) );
  INV_X1 stateFF_state_gff_5_SFF_3_U3 ( .A(stateFF_state_n9), .ZN(
        stateFF_state_gff_5_SFF_3_n10) );
  INV_X1 stateFF_state_gff_5_SFF_3_U2 ( .A(stateFF_state_gff_5_SFF_3_n10), 
        .ZN(stateFF_state_gff_5_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_5_SFF_3_Cell_reg ( .D(stateFF_state_gff_5_SFF_3_n6), 
        .CK(clk), .Q(stateFF_inputPar[53]), .QN(stateFF_state_gff_5_SFF_3_n7)
         );
  BUF_X1 stateFF_state_gff_6_U2 ( .A(selP), .Z(stateFF_state_gff_6_n2) );
  OAI21_X1 stateFF_state_gff_6_SFF_0_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_6_SFF_0_n8), .A(stateFF_state_gff_6_SFF_0_n11), .ZN(
        stateFF_state_gff_6_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_6_SFF_0_U3 ( .B1(stateFF_state_gff_6_n2), .B2(
        stateFF_inputPar[5]), .C1(stateFF_state_gff_6_SFF_0_n10), .C2(
        stateFF_inputPar[20]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_6_SFF_0_n11) );
  INV_X1 stateFF_state_gff_6_SFF_0_U2 ( .A(stateFF_state_gff_6_n2), .ZN(
        stateFF_state_gff_6_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_6_SFF_0_Cell_reg ( .D(stateFF_state_gff_6_SFF_0_n7), 
        .CK(clk), .Q(stateFF_inputPar[6]), .QN(stateFF_state_gff_6_SFF_0_n8)
         );
  OAI21_X1 stateFF_state_gff_6_SFF_1_U3 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_6_SFF_1_n8), .A(stateFF_state_gff_6_SFF_1_n10), .ZN(
        stateFF_state_gff_6_SFF_1_n7) );
  NAND2_X1 stateFF_state_gff_6_SFF_1_U2 ( .A1(stateFF_state_n7), .A2(
        stateFF_n[48]), .ZN(stateFF_state_gff_6_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_6_SFF_1_Cell_reg ( .D(stateFF_state_gff_6_SFF_1_n7), 
        .CK(clk), .Q(stateFF_inputPar[22]), .QN(stateFF_state_gff_6_SFF_1_n8)
         );
  OAI21_X1 stateFF_state_gff_6_SFF_2_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_6_SFF_2_n8), .A(stateFF_state_gff_6_SFF_2_n11), .ZN(
        stateFF_state_gff_6_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_6_SFF_2_U3 ( .B1(stateFF_state_gff_6_n2), .B2(
        stateFF_inputPar[37]), .C1(stateFF_state_gff_6_SFF_2_n10), .C2(
        stateFF_inputPar[22]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_6_SFF_2_n11) );
  INV_X1 stateFF_state_gff_6_SFF_2_U2 ( .A(stateFF_state_gff_6_n2), .ZN(
        stateFF_state_gff_6_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_6_SFF_2_Cell_reg ( .D(stateFF_state_gff_6_SFF_2_n7), 
        .CK(clk), .Q(stateFF_inputPar[38]), .QN(stateFF_state_gff_6_SFF_2_n8)
         );
  OAI21_X1 stateFF_state_gff_6_SFF_3_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_6_SFF_3_n8), .A(stateFF_state_gff_6_SFF_3_n11), .ZN(
        stateFF_state_gff_6_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_6_SFF_3_U3 ( .B1(stateFF_state_gff_6_n2), .B2(
        stateFF_inputPar[53]), .C1(stateFF_state_gff_6_SFF_3_n10), .C2(
        stateFF_inputPar[23]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_6_SFF_3_n11) );
  INV_X1 stateFF_state_gff_6_SFF_3_U2 ( .A(stateFF_state_gff_6_n2), .ZN(
        stateFF_state_gff_6_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_6_SFF_3_Cell_reg ( .D(stateFF_state_gff_6_SFF_3_n7), 
        .CK(clk), .Q(stateFF_inputPar[54]), .QN(stateFF_state_gff_6_SFF_3_n8)
         );
  OAI21_X1 stateFF_state_gff_7_SFF_0_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_7_SFF_0_n8), .A(stateFF_state_gff_7_SFF_0_n12), .ZN(
        stateFF_state_gff_7_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_7_SFF_0_U4 ( .B1(stateFF_state_gff_7_SFF_0_n10), 
        .B2(stateFF_inputPar[6]), .C1(stateFF_state_gff_7_SFF_0_n11), .C2(
        stateFF_inputPar[24]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_7_SFF_0_n12) );
  INV_X1 stateFF_state_gff_7_SFF_0_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_7_SFF_0_n11) );
  INV_X1 stateFF_state_gff_7_SFF_0_U2 ( .A(stateFF_state_gff_7_SFF_0_n11), 
        .ZN(stateFF_state_gff_7_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_7_SFF_0_Cell_reg ( .D(stateFF_state_gff_7_SFF_0_n7), 
        .CK(clk), .Q(stateFF_inputPar[7]), .QN(stateFF_state_gff_7_SFF_0_n8)
         );
  OAI21_X1 stateFF_state_gff_7_SFF_1_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_7_SFF_1_n8), .A(stateFF_state_gff_7_SFF_1_n12), .ZN(
        stateFF_state_gff_7_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_7_SFF_1_U4 ( .B1(stateFF_state_gff_7_SFF_1_n10), 
        .B2(stateFF_inputPar[22]), .C1(stateFF_state_gff_7_SFF_1_n11), .C2(
        stateFF_inputPar[25]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_7_SFF_1_n12) );
  INV_X1 stateFF_state_gff_7_SFF_1_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_7_SFF_1_n11) );
  INV_X1 stateFF_state_gff_7_SFF_1_U2 ( .A(stateFF_state_gff_7_SFF_1_n11), 
        .ZN(stateFF_state_gff_7_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_7_SFF_1_Cell_reg ( .D(stateFF_state_gff_7_SFF_1_n7), 
        .CK(clk), .Q(stateFF_inputPar[23]), .QN(stateFF_state_gff_7_SFF_1_n8)
         );
  OAI21_X1 stateFF_state_gff_7_SFF_2_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_7_SFF_2_n8), .A(stateFF_state_gff_7_SFF_2_n12), .ZN(
        stateFF_state_gff_7_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_7_SFF_2_U4 ( .B1(stateFF_state_gff_7_SFF_2_n10), 
        .B2(stateFF_inputPar[38]), .C1(stateFF_state_gff_7_SFF_2_n11), .C2(
        stateFF_inputPar[26]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_7_SFF_2_n12) );
  INV_X1 stateFF_state_gff_7_SFF_2_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_7_SFF_2_n11) );
  INV_X1 stateFF_state_gff_7_SFF_2_U2 ( .A(stateFF_state_gff_7_SFF_2_n11), 
        .ZN(stateFF_state_gff_7_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_7_SFF_2_Cell_reg ( .D(stateFF_state_gff_7_SFF_2_n7), 
        .CK(clk), .Q(stateFF_inputPar[39]), .QN(stateFF_state_gff_7_SFF_2_n8)
         );
  OAI21_X1 stateFF_state_gff_7_SFF_3_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_7_SFF_3_n8), .A(stateFF_state_gff_7_SFF_3_n12), .ZN(
        stateFF_state_gff_7_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_7_SFF_3_U4 ( .B1(stateFF_state_gff_7_SFF_3_n10), 
        .B2(stateFF_inputPar[54]), .C1(stateFF_state_gff_7_SFF_3_n11), .C2(
        stateFF_inputPar[27]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_7_SFF_3_n12) );
  INV_X1 stateFF_state_gff_7_SFF_3_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_7_SFF_3_n11) );
  INV_X1 stateFF_state_gff_7_SFF_3_U2 ( .A(stateFF_state_gff_7_SFF_3_n11), 
        .ZN(stateFF_state_gff_7_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_7_SFF_3_Cell_reg ( .D(stateFF_state_gff_7_SFF_3_n7), 
        .CK(clk), .Q(stateFF_inputPar[55]), .QN(stateFF_state_gff_7_SFF_3_n8)
         );
  OAI21_X1 stateFF_state_gff_8_SFF_0_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_8_SFF_0_n8), .A(stateFF_state_gff_8_SFF_0_n12), .ZN(
        stateFF_state_gff_8_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_8_SFF_0_U4 ( .B1(stateFF_state_gff_8_SFF_0_n10), 
        .B2(stateFF_inputPar[7]), .C1(stateFF_state_gff_8_SFF_0_n11), .C2(
        stateFF_inputPar[28]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_8_SFF_0_n12) );
  INV_X1 stateFF_state_gff_8_SFF_0_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_8_SFF_0_n11) );
  INV_X1 stateFF_state_gff_8_SFF_0_U2 ( .A(stateFF_state_gff_8_SFF_0_n11), 
        .ZN(stateFF_state_gff_8_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_8_SFF_0_Cell_reg ( .D(stateFF_state_gff_8_SFF_0_n7), 
        .CK(clk), .Q(stateFF_inputPar[8]), .QN(stateFF_state_gff_8_SFF_0_n8)
         );
  OAI21_X1 stateFF_state_gff_8_SFF_1_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_8_SFF_1_n8), .A(stateFF_state_gff_8_SFF_1_n12), .ZN(
        stateFF_state_gff_8_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_8_SFF_1_U4 ( .B1(stateFF_state_gff_8_SFF_1_n10), 
        .B2(stateFF_inputPar[23]), .C1(stateFF_state_gff_8_SFF_1_n11), .C2(
        stateFF_inputPar[29]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_8_SFF_1_n12) );
  INV_X1 stateFF_state_gff_8_SFF_1_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_8_SFF_1_n11) );
  INV_X1 stateFF_state_gff_8_SFF_1_U2 ( .A(stateFF_state_gff_8_SFF_1_n11), 
        .ZN(stateFF_state_gff_8_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_8_SFF_1_Cell_reg ( .D(stateFF_state_gff_8_SFF_1_n7), 
        .CK(clk), .Q(stateFF_inputPar[24]), .QN(stateFF_state_gff_8_SFF_1_n8)
         );
  OAI21_X1 stateFF_state_gff_8_SFF_2_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_8_SFF_2_n7), .A(stateFF_state_gff_8_SFF_2_n11), .ZN(
        stateFF_state_gff_8_SFF_2_n6) );
  OAI221_X1 stateFF_state_gff_8_SFF_2_U4 ( .B1(stateFF_state_gff_8_SFF_2_n9), 
        .B2(stateFF_inputPar[39]), .C1(stateFF_state_gff_8_SFF_2_n10), .C2(
        stateFF_inputPar[30]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_8_SFF_2_n11) );
  INV_X1 stateFF_state_gff_8_SFF_2_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_8_SFF_2_n10) );
  INV_X1 stateFF_state_gff_8_SFF_2_U2 ( .A(stateFF_state_gff_8_SFF_2_n10), 
        .ZN(stateFF_state_gff_8_SFF_2_n9) );
  DFF_X1 stateFF_state_gff_8_SFF_2_Cell_reg ( .D(stateFF_state_gff_8_SFF_2_n6), 
        .CK(clk), .Q(stateFF_inputPar[40]), .QN(stateFF_state_gff_8_SFF_2_n7)
         );
  OAI21_X1 stateFF_state_gff_8_SFF_3_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_8_SFF_3_n7), .A(stateFF_state_gff_8_SFF_3_n11), .ZN(
        stateFF_state_gff_8_SFF_3_n6) );
  OAI221_X1 stateFF_state_gff_8_SFF_3_U4 ( .B1(stateFF_state_gff_8_SFF_3_n9), 
        .B2(stateFF_inputPar[55]), .C1(stateFF_state_gff_8_SFF_3_n10), .C2(
        stateFF_inputPar[31]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_8_SFF_3_n11) );
  INV_X1 stateFF_state_gff_8_SFF_3_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_8_SFF_3_n10) );
  INV_X1 stateFF_state_gff_8_SFF_3_U2 ( .A(stateFF_state_gff_8_SFF_3_n10), 
        .ZN(stateFF_state_gff_8_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_8_SFF_3_Cell_reg ( .D(stateFF_state_gff_8_SFF_3_n6), 
        .CK(clk), .Q(stateFF_inputPar[56]), .QN(stateFF_state_gff_8_SFF_3_n7)
         );
  OAI21_X1 stateFF_state_gff_9_SFF_0_U5 ( .B1(enKey), .B2(
        stateFF_state_gff_9_SFF_0_n7), .A(stateFF_state_gff_9_SFF_0_n11), .ZN(
        stateFF_state_gff_9_SFF_0_n6) );
  OAI221_X1 stateFF_state_gff_9_SFF_0_U4 ( .B1(stateFF_state_gff_9_SFF_0_n9), 
        .B2(stateFF_inputPar[8]), .C1(stateFF_state_gff_9_SFF_0_n10), .C2(
        stateFF_inputPar[32]), .A(enKey), .ZN(stateFF_state_gff_9_SFF_0_n11)
         );
  INV_X1 stateFF_state_gff_9_SFF_0_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_9_SFF_0_n10) );
  INV_X1 stateFF_state_gff_9_SFF_0_U2 ( .A(stateFF_state_gff_9_SFF_0_n10), 
        .ZN(stateFF_state_gff_9_SFF_0_n9) );
  DFF_X1 stateFF_state_gff_9_SFF_0_Cell_reg ( .D(stateFF_state_gff_9_SFF_0_n6), 
        .CK(clk), .Q(stateFF_inputPar[9]), .QN(stateFF_state_gff_9_SFF_0_n7)
         );
  OAI21_X1 stateFF_state_gff_9_SFF_1_U5 ( .B1(enKey), .B2(
        stateFF_state_gff_9_SFF_1_n7), .A(stateFF_state_gff_9_SFF_1_n11), .ZN(
        stateFF_state_gff_9_SFF_1_n6) );
  OAI221_X1 stateFF_state_gff_9_SFF_1_U4 ( .B1(stateFF_state_gff_9_SFF_1_n9), 
        .B2(stateFF_inputPar[24]), .C1(stateFF_state_gff_9_SFF_1_n10), .C2(
        stateFF_inputPar[33]), .A(enKey), .ZN(stateFF_state_gff_9_SFF_1_n11)
         );
  INV_X1 stateFF_state_gff_9_SFF_1_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_9_SFF_1_n10) );
  INV_X1 stateFF_state_gff_9_SFF_1_U2 ( .A(stateFF_state_gff_9_SFF_1_n10), 
        .ZN(stateFF_state_gff_9_SFF_1_n9) );
  DFF_X1 stateFF_state_gff_9_SFF_1_Cell_reg ( .D(stateFF_state_gff_9_SFF_1_n6), 
        .CK(clk), .Q(stateFF_inputPar[25]), .QN(stateFF_state_gff_9_SFF_1_n7)
         );
  OAI21_X1 stateFF_state_gff_9_SFF_2_U5 ( .B1(enKey), .B2(
        stateFF_state_gff_9_SFF_2_n7), .A(stateFF_state_gff_9_SFF_2_n11), .ZN(
        stateFF_state_gff_9_SFF_2_n6) );
  OAI221_X1 stateFF_state_gff_9_SFF_2_U4 ( .B1(stateFF_state_gff_9_SFF_2_n9), 
        .B2(stateFF_inputPar[40]), .C1(stateFF_state_gff_9_SFF_2_n10), .C2(
        stateFF_inputPar[34]), .A(enKey), .ZN(stateFF_state_gff_9_SFF_2_n11)
         );
  INV_X1 stateFF_state_gff_9_SFF_2_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_9_SFF_2_n10) );
  INV_X1 stateFF_state_gff_9_SFF_2_U2 ( .A(stateFF_state_gff_9_SFF_2_n10), 
        .ZN(stateFF_state_gff_9_SFF_2_n9) );
  DFF_X1 stateFF_state_gff_9_SFF_2_Cell_reg ( .D(stateFF_state_gff_9_SFF_2_n6), 
        .CK(clk), .Q(stateFF_inputPar[41]), .QN(stateFF_state_gff_9_SFF_2_n7)
         );
  OAI21_X1 stateFF_state_gff_9_SFF_3_U5 ( .B1(enKey), .B2(
        stateFF_state_gff_9_SFF_3_n7), .A(stateFF_state_gff_9_SFF_3_n11), .ZN(
        stateFF_state_gff_9_SFF_3_n6) );
  OAI221_X1 stateFF_state_gff_9_SFF_3_U4 ( .B1(stateFF_state_gff_9_SFF_3_n9), 
        .B2(stateFF_inputPar[56]), .C1(stateFF_state_gff_9_SFF_3_n10), .C2(
        stateFF_inputPar[35]), .A(enKey), .ZN(stateFF_state_gff_9_SFF_3_n11)
         );
  INV_X1 stateFF_state_gff_9_SFF_3_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_9_SFF_3_n10) );
  INV_X1 stateFF_state_gff_9_SFF_3_U2 ( .A(stateFF_state_gff_9_SFF_3_n10), 
        .ZN(stateFF_state_gff_9_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_9_SFF_3_Cell_reg ( .D(stateFF_state_gff_9_SFF_3_n6), 
        .CK(clk), .Q(stateFF_inputPar[57]), .QN(stateFF_state_gff_9_SFF_3_n7)
         );
  OAI21_X1 stateFF_state_gff_10_SFF_0_U5 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_10_SFF_0_n8), .A(stateFF_state_gff_10_SFF_0_n12), 
        .ZN(stateFF_state_gff_10_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_10_SFF_0_U4 ( .B1(stateFF_state_gff_10_SFF_0_n10), .B2(stateFF_inputPar[9]), .C1(stateFF_state_gff_10_SFF_0_n11), .C2(
        stateFF_inputPar[36]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_10_SFF_0_n12) );
  INV_X1 stateFF_state_gff_10_SFF_0_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_10_SFF_0_n11) );
  INV_X1 stateFF_state_gff_10_SFF_0_U2 ( .A(stateFF_state_gff_10_SFF_0_n11), 
        .ZN(stateFF_state_gff_10_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_10_SFF_0_Cell_reg ( .D(
        stateFF_state_gff_10_SFF_0_n7), .CK(clk), .Q(stateFF_inputPar[10]), 
        .QN(stateFF_state_gff_10_SFF_0_n8) );
  OAI21_X1 stateFF_state_gff_10_SFF_1_U5 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_10_SFF_1_n8), .A(stateFF_state_gff_10_SFF_1_n12), 
        .ZN(stateFF_state_gff_10_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_10_SFF_1_U4 ( .B1(stateFF_state_gff_10_SFF_1_n10), .B2(stateFF_inputPar[25]), .C1(stateFF_state_gff_10_SFF_1_n11), .C2(
        stateFF_inputPar[37]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_10_SFF_1_n12) );
  INV_X1 stateFF_state_gff_10_SFF_1_U3 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_10_SFF_1_n11) );
  INV_X1 stateFF_state_gff_10_SFF_1_U2 ( .A(stateFF_state_gff_10_SFF_1_n11), 
        .ZN(stateFF_state_gff_10_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_10_SFF_1_Cell_reg ( .D(
        stateFF_state_gff_10_SFF_1_n7), .CK(clk), .Q(stateFF_inputPar[26]), 
        .QN(stateFF_state_gff_10_SFF_1_n8) );
  OAI21_X1 stateFF_state_gff_10_SFF_2_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_10_SFF_2_n8), .A(stateFF_state_gff_10_SFF_2_n11), 
        .ZN(stateFF_state_gff_10_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_10_SFF_2_U3 ( .B1(stateFF_state_n11), .B2(
        stateFF_inputPar[41]), .C1(stateFF_state_gff_10_SFF_2_n10), .C2(
        stateFF_inputPar[38]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_10_SFF_2_n11) );
  INV_X1 stateFF_state_gff_10_SFF_2_U2 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_10_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_10_SFF_2_Cell_reg ( .D(
        stateFF_state_gff_10_SFF_2_n7), .CK(clk), .Q(stateFF_n[27]), .QN(
        stateFF_state_gff_10_SFF_2_n8) );
  OAI21_X1 stateFF_state_gff_10_SFF_3_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_10_SFF_3_n8), .A(stateFF_state_gff_10_SFF_3_n11), 
        .ZN(stateFF_state_gff_10_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_10_SFF_3_U3 ( .B1(stateFF_state_n11), .B2(
        stateFF_inputPar[57]), .C1(stateFF_state_gff_10_SFF_3_n10), .C2(
        stateFF_inputPar[39]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_10_SFF_3_n11) );
  INV_X1 stateFF_state_gff_10_SFF_3_U2 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_10_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_10_SFF_3_Cell_reg ( .D(
        stateFF_state_gff_10_SFF_3_n7), .CK(clk), .Q(stateFF_inputPar[58]), 
        .QN(stateFF_state_gff_10_SFF_3_n8) );
  BUF_X1 stateFF_state_gff_11_U2 ( .A(stateFF_state_n11), .Z(
        stateFF_state_gff_11_n2) );
  OAI21_X1 stateFF_state_gff_11_SFF_0_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_11_SFF_0_n8), .A(stateFF_state_gff_11_SFF_0_n11), 
        .ZN(stateFF_state_gff_11_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_11_SFF_0_U3 ( .B1(stateFF_state_gff_11_n2), .B2(
        stateFF_inputPar[10]), .C1(stateFF_state_gff_11_SFF_0_n10), .C2(
        stateFF_inputPar[40]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_11_SFF_0_n11) );
  INV_X1 stateFF_state_gff_11_SFF_0_U2 ( .A(stateFF_state_gff_11_n2), .ZN(
        stateFF_state_gff_11_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_11_SFF_0_Cell_reg ( .D(
        stateFF_state_gff_11_SFF_0_n7), .CK(clk), .Q(stateFF_inputPar[11]), 
        .QN(stateFF_state_gff_11_SFF_0_n8) );
  OAI21_X1 stateFF_state_gff_11_SFF_1_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_11_SFF_1_n8), .A(stateFF_state_gff_11_SFF_1_n11), 
        .ZN(stateFF_state_gff_11_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_11_SFF_1_U3 ( .B1(stateFF_state_gff_11_n2), .B2(
        stateFF_inputPar[26]), .C1(stateFF_state_gff_11_SFF_1_n10), .C2(
        stateFF_inputPar[41]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_11_SFF_1_n11) );
  INV_X1 stateFF_state_gff_11_SFF_1_U2 ( .A(stateFF_state_gff_11_n2), .ZN(
        stateFF_state_gff_11_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_11_SFF_1_Cell_reg ( .D(
        stateFF_state_gff_11_SFF_1_n7), .CK(clk), .Q(stateFF_inputPar[27]), 
        .QN(stateFF_state_gff_11_SFF_1_n8) );
  OAI21_X1 stateFF_state_gff_11_SFF_2_U3 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_11_SFF_2_n8), .A(stateFF_state_gff_11_SFF_2_n10), 
        .ZN(stateFF_state_gff_11_SFF_2_n7) );
  NAND2_X1 stateFF_state_gff_11_SFF_2_U2 ( .A1(stateFF_state_n7), .A2(
        stateFF_n[27]), .ZN(stateFF_state_gff_11_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_11_SFF_2_Cell_reg ( .D(
        stateFF_state_gff_11_SFF_2_n7), .CK(clk), .Q(stateFF_inputPar[43]), 
        .QN(stateFF_state_gff_11_SFF_2_n8) );
  OAI21_X1 stateFF_state_gff_11_SFF_3_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_11_SFF_3_n8), .A(stateFF_state_gff_11_SFF_3_n11), 
        .ZN(stateFF_state_gff_11_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_11_SFF_3_U3 ( .B1(stateFF_state_gff_11_n2), .B2(
        stateFF_inputPar[58]), .C1(stateFF_state_gff_11_SFF_3_n10), .C2(
        stateFF_inputPar[43]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_11_SFF_3_n11) );
  INV_X1 stateFF_state_gff_11_SFF_3_U2 ( .A(stateFF_state_gff_11_n2), .ZN(
        stateFF_state_gff_11_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_11_SFF_3_Cell_reg ( .D(
        stateFF_state_gff_11_SFF_3_n7), .CK(clk), .Q(stateFF_inputPar[59]), 
        .QN(stateFF_state_gff_11_SFF_3_n8) );
  OAI21_X1 stateFF_state_gff_12_SFF_0_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_12_SFF_0_n8), .A(stateFF_state_gff_12_SFF_0_n11), 
        .ZN(stateFF_state_gff_12_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_12_SFF_0_U3 ( .B1(stateFF_state_n10), .B2(
        stateFF_inputPar[11]), .C1(stateFF_state_gff_12_SFF_0_n10), .C2(
        stateFF_inputPar[44]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_12_SFF_0_n11) );
  INV_X1 stateFF_state_gff_12_SFF_0_U2 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_12_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_12_SFF_0_Cell_reg ( .D(
        stateFF_state_gff_12_SFF_0_n7), .CK(clk), .Q(stateFF_inputPar[12]), 
        .QN(stateFF_state_gff_12_SFF_0_n8) );
  OAI21_X1 stateFF_state_gff_12_SFF_1_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_12_SFF_1_n8), .A(stateFF_state_gff_12_SFF_1_n11), 
        .ZN(stateFF_state_gff_12_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_12_SFF_1_U3 ( .B1(stateFF_state_n10), .B2(
        stateFF_inputPar[27]), .C1(stateFF_state_gff_12_SFF_1_n10), .C2(
        stateFF_inputPar[45]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_12_SFF_1_n11) );
  INV_X1 stateFF_state_gff_12_SFF_1_U2 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_12_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_12_SFF_1_Cell_reg ( .D(
        stateFF_state_gff_12_SFF_1_n7), .CK(clk), .Q(stateFF_inputPar[28]), 
        .QN(stateFF_state_gff_12_SFF_1_n8) );
  OAI21_X1 stateFF_state_gff_12_SFF_2_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_12_SFF_2_n7), .A(stateFF_state_gff_12_SFF_2_n11), 
        .ZN(stateFF_state_gff_12_SFF_2_n6) );
  OAI221_X1 stateFF_state_gff_12_SFF_2_U4 ( .B1(stateFF_state_gff_12_SFF_2_n9), 
        .B2(stateFF_inputPar[43]), .C1(stateFF_state_gff_12_SFF_2_n10), .C2(
        stateFF_inputPar[46]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_12_SFF_2_n11) );
  INV_X1 stateFF_state_gff_12_SFF_2_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_12_SFF_2_n10) );
  INV_X1 stateFF_state_gff_12_SFF_2_U2 ( .A(stateFF_state_gff_12_SFF_2_n10), 
        .ZN(stateFF_state_gff_12_SFF_2_n9) );
  DFF_X1 stateFF_state_gff_12_SFF_2_Cell_reg ( .D(
        stateFF_state_gff_12_SFF_2_n6), .CK(clk), .Q(stateFF_inputPar[44]), 
        .QN(stateFF_state_gff_12_SFF_2_n7) );
  OAI21_X1 stateFF_state_gff_12_SFF_3_U5 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_12_SFF_3_n7), .A(stateFF_state_gff_12_SFF_3_n11), 
        .ZN(stateFF_state_gff_12_SFF_3_n6) );
  OAI221_X1 stateFF_state_gff_12_SFF_3_U4 ( .B1(stateFF_state_gff_12_SFF_3_n9), 
        .B2(stateFF_inputPar[59]), .C1(stateFF_state_gff_12_SFF_3_n10), .C2(
        stateFF_inputPar[47]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_12_SFF_3_n11) );
  INV_X1 stateFF_state_gff_12_SFF_3_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_12_SFF_3_n10) );
  INV_X1 stateFF_state_gff_12_SFF_3_U2 ( .A(stateFF_state_gff_12_SFF_3_n10), 
        .ZN(stateFF_state_gff_12_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_12_SFF_3_Cell_reg ( .D(
        stateFF_state_gff_12_SFF_3_n6), .CK(clk), .Q(stateFF_inputPar[60]), 
        .QN(stateFF_state_gff_12_SFF_3_n7) );
  OAI21_X1 stateFF_state_gff_13_SFF_0_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_13_SFF_0_n7), .A(stateFF_state_gff_13_SFF_0_n11), 
        .ZN(stateFF_state_gff_13_SFF_0_n6) );
  OAI221_X1 stateFF_state_gff_13_SFF_0_U4 ( .B1(stateFF_state_gff_13_SFF_0_n9), 
        .B2(stateFF_inputPar[12]), .C1(stateFF_state_gff_13_SFF_0_n10), .C2(
        stateFF_inputPar[48]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_13_SFF_0_n11) );
  INV_X1 stateFF_state_gff_13_SFF_0_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_13_SFF_0_n10) );
  INV_X1 stateFF_state_gff_13_SFF_0_U2 ( .A(stateFF_state_gff_13_SFF_0_n10), 
        .ZN(stateFF_state_gff_13_SFF_0_n9) );
  DFF_X1 stateFF_state_gff_13_SFF_0_Cell_reg ( .D(
        stateFF_state_gff_13_SFF_0_n6), .CK(clk), .Q(stateFF_inputPar[13]), 
        .QN(stateFF_state_gff_13_SFF_0_n7) );
  OAI21_X1 stateFF_state_gff_13_SFF_1_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_13_SFF_1_n7), .A(stateFF_state_gff_13_SFF_1_n11), 
        .ZN(stateFF_state_gff_13_SFF_1_n6) );
  OAI221_X1 stateFF_state_gff_13_SFF_1_U4 ( .B1(stateFF_state_gff_13_SFF_1_n9), 
        .B2(stateFF_inputPar[28]), .C1(stateFF_state_gff_13_SFF_1_n10), .C2(
        stateFF_inputPar[49]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_13_SFF_1_n11) );
  INV_X1 stateFF_state_gff_13_SFF_1_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_13_SFF_1_n10) );
  INV_X1 stateFF_state_gff_13_SFF_1_U2 ( .A(stateFF_state_gff_13_SFF_1_n10), 
        .ZN(stateFF_state_gff_13_SFF_1_n9) );
  DFF_X1 stateFF_state_gff_13_SFF_1_Cell_reg ( .D(
        stateFF_state_gff_13_SFF_1_n6), .CK(clk), .Q(stateFF_inputPar[29]), 
        .QN(stateFF_state_gff_13_SFF_1_n7) );
  OAI21_X1 stateFF_state_gff_13_SFF_2_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_13_SFF_2_n7), .A(stateFF_state_gff_13_SFF_2_n11), 
        .ZN(stateFF_state_gff_13_SFF_2_n6) );
  OAI221_X1 stateFF_state_gff_13_SFF_2_U4 ( .B1(stateFF_state_gff_13_SFF_2_n9), 
        .B2(stateFF_inputPar[44]), .C1(stateFF_state_gff_13_SFF_2_n10), .C2(
        stateFF_inputPar[50]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_13_SFF_2_n11) );
  INV_X1 stateFF_state_gff_13_SFF_2_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_13_SFF_2_n10) );
  INV_X1 stateFF_state_gff_13_SFF_2_U2 ( .A(stateFF_state_gff_13_SFF_2_n10), 
        .ZN(stateFF_state_gff_13_SFF_2_n9) );
  DFF_X1 stateFF_state_gff_13_SFF_2_Cell_reg ( .D(
        stateFF_state_gff_13_SFF_2_n6), .CK(clk), .Q(stateFF_inputPar[45]), 
        .QN(stateFF_state_gff_13_SFF_2_n7) );
  OAI21_X1 stateFF_state_gff_13_SFF_3_U5 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_13_SFF_3_n7), .A(stateFF_state_gff_13_SFF_3_n11), 
        .ZN(stateFF_state_gff_13_SFF_3_n6) );
  OAI221_X1 stateFF_state_gff_13_SFF_3_U4 ( .B1(stateFF_state_gff_13_SFF_3_n9), 
        .B2(stateFF_inputPar[60]), .C1(stateFF_state_gff_13_SFF_3_n10), .C2(
        stateFF_inputPar[51]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_13_SFF_3_n11) );
  INV_X1 stateFF_state_gff_13_SFF_3_U3 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_13_SFF_3_n10) );
  INV_X1 stateFF_state_gff_13_SFF_3_U2 ( .A(stateFF_state_gff_13_SFF_3_n10), 
        .ZN(stateFF_state_gff_13_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_13_SFF_3_Cell_reg ( .D(
        stateFF_state_gff_13_SFF_3_n6), .CK(clk), .Q(stateFF_inputPar[61]), 
        .QN(stateFF_state_gff_13_SFF_3_n7) );
  OAI21_X1 stateFF_state_gff_14_SFF_0_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_14_SFF_0_n8), .A(stateFF_state_gff_14_SFF_0_n11), 
        .ZN(stateFF_state_gff_14_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_14_SFF_0_U3 ( .B1(stateFF_state_n11), .B2(
        stateFF_inputPar[13]), .C1(stateFF_state_gff_14_SFF_0_n10), .C2(
        stateFF_inputPar[52]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_14_SFF_0_n11) );
  INV_X1 stateFF_state_gff_14_SFF_0_U2 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_14_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_14_SFF_0_Cell_reg ( .D(
        stateFF_state_gff_14_SFF_0_n7), .CK(clk), .Q(stateFF_inputPar[14]), 
        .QN(stateFF_state_gff_14_SFF_0_n8) );
  OAI21_X1 stateFF_state_gff_14_SFF_1_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_14_SFF_1_n8), .A(stateFF_state_gff_14_SFF_1_n11), 
        .ZN(stateFF_state_gff_14_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_14_SFF_1_U3 ( .B1(stateFF_state_n11), .B2(
        stateFF_inputPar[29]), .C1(stateFF_state_gff_14_SFF_1_n10), .C2(
        stateFF_inputPar[53]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_14_SFF_1_n11) );
  INV_X1 stateFF_state_gff_14_SFF_1_U2 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_14_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_14_SFF_1_Cell_reg ( .D(
        stateFF_state_gff_14_SFF_1_n7), .CK(clk), .Q(stateFF_inputPar[30]), 
        .QN(stateFF_state_gff_14_SFF_1_n8) );
  OAI21_X1 stateFF_state_gff_14_SFF_2_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_14_SFF_2_n8), .A(stateFF_state_gff_14_SFF_2_n11), 
        .ZN(stateFF_state_gff_14_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_14_SFF_2_U3 ( .B1(stateFF_state_n11), .B2(
        stateFF_inputPar[45]), .C1(stateFF_state_gff_14_SFF_2_n10), .C2(
        stateFF_inputPar[54]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_14_SFF_2_n11) );
  INV_X1 stateFF_state_gff_14_SFF_2_U2 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_14_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_14_SFF_2_Cell_reg ( .D(
        stateFF_state_gff_14_SFF_2_n7), .CK(clk), .Q(stateFF_inputPar[46]), 
        .QN(stateFF_state_gff_14_SFF_2_n8) );
  OAI21_X1 stateFF_state_gff_14_SFF_3_U4 ( .B1(stateFF_state_n8), .B2(
        stateFF_state_gff_14_SFF_3_n8), .A(stateFF_state_gff_14_SFF_3_n11), 
        .ZN(stateFF_state_gff_14_SFF_3_n7) );
  OAI221_X1 stateFF_state_gff_14_SFF_3_U3 ( .B1(stateFF_state_n11), .B2(
        stateFF_inputPar[61]), .C1(stateFF_state_gff_14_SFF_3_n10), .C2(
        stateFF_inputPar[55]), .A(stateFF_state_n8), .ZN(
        stateFF_state_gff_14_SFF_3_n11) );
  INV_X1 stateFF_state_gff_14_SFF_3_U2 ( .A(stateFF_state_n11), .ZN(
        stateFF_state_gff_14_SFF_3_n10) );
  DFF_X1 stateFF_state_gff_14_SFF_3_Cell_reg ( .D(
        stateFF_state_gff_14_SFF_3_n7), .CK(clk), .Q(stateFF_inputPar[62]), 
        .QN(stateFF_state_gff_14_SFF_3_n8) );
  OAI21_X1 stateFF_state_gff_15_SFF_0_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_15_SFF_0_n8), .A(stateFF_state_gff_15_SFF_0_n11), 
        .ZN(stateFF_state_gff_15_SFF_0_n7) );
  OAI221_X1 stateFF_state_gff_15_SFF_0_U3 ( .B1(stateFF_state_n10), .B2(
        stateFF_inputPar[14]), .C1(stateFF_state_gff_15_SFF_0_n10), .C2(
        stateFF_inputPar[56]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_15_SFF_0_n11) );
  INV_X1 stateFF_state_gff_15_SFF_0_U2 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_15_SFF_0_n10) );
  DFF_X1 stateFF_state_gff_15_SFF_0_Cell_reg ( .D(
        stateFF_state_gff_15_SFF_0_n7), .CK(clk), .Q(stateFF_inputPar[15]), 
        .QN(stateFF_state_gff_15_SFF_0_n8) );
  OAI21_X1 stateFF_state_gff_15_SFF_1_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_15_SFF_1_n8), .A(stateFF_state_gff_15_SFF_1_n11), 
        .ZN(stateFF_state_gff_15_SFF_1_n7) );
  OAI221_X1 stateFF_state_gff_15_SFF_1_U3 ( .B1(stateFF_state_n10), .B2(
        stateFF_inputPar[30]), .C1(stateFF_state_gff_15_SFF_1_n10), .C2(
        stateFF_inputPar[57]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_15_SFF_1_n11) );
  INV_X1 stateFF_state_gff_15_SFF_1_U2 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_15_SFF_1_n10) );
  DFF_X1 stateFF_state_gff_15_SFF_1_Cell_reg ( .D(
        stateFF_state_gff_15_SFF_1_n7), .CK(clk), .Q(stateFF_inputPar[31]), 
        .QN(stateFF_state_gff_15_SFF_1_n8) );
  OAI21_X1 stateFF_state_gff_15_SFF_2_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_15_SFF_2_n8), .A(stateFF_state_gff_15_SFF_2_n11), 
        .ZN(stateFF_state_gff_15_SFF_2_n7) );
  OAI221_X1 stateFF_state_gff_15_SFF_2_U3 ( .B1(stateFF_state_n10), .B2(
        stateFF_inputPar[46]), .C1(stateFF_state_gff_15_SFF_2_n10), .C2(
        stateFF_inputPar[58]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_15_SFF_2_n11) );
  INV_X1 stateFF_state_gff_15_SFF_2_U2 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_15_SFF_2_n10) );
  DFF_X1 stateFF_state_gff_15_SFF_2_Cell_reg ( .D(
        stateFF_state_gff_15_SFF_2_n7), .CK(clk), .Q(stateFF_inputPar[47]), 
        .QN(stateFF_state_gff_15_SFF_2_n8) );
  OAI21_X1 stateFF_state_gff_15_SFF_3_U4 ( .B1(stateFF_state_n6), .B2(
        stateFF_state_gff_15_SFF_3_n7), .A(stateFF_state_gff_15_SFF_3_n10), 
        .ZN(stateFF_state_gff_15_SFF_3_n6) );
  OAI221_X1 stateFF_state_gff_15_SFF_3_U3 ( .B1(stateFF_state_n10), .B2(
        stateFF_inputPar[62]), .C1(stateFF_state_gff_15_SFF_3_n9), .C2(
        stateFF_inputPar[59]), .A(stateFF_state_n6), .ZN(
        stateFF_state_gff_15_SFF_3_n10) );
  INV_X1 stateFF_state_gff_15_SFF_3_U2 ( .A(stateFF_state_n10), .ZN(
        stateFF_state_gff_15_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_15_SFF_3_Cell_reg ( .D(
        stateFF_state_gff_15_SFF_3_n6), .CK(clk), .Q(stateFF_n[6]), .QN(
        stateFF_state_gff_15_SFF_3_n7) );
  BUF_X1 stateFF_state_gff_16_U2 ( .A(stateFF_state_n9), .Z(
        stateFF_state_gff_16_n2) );
  OAI21_X1 stateFF_state_gff_16_SFF_0_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_16_SFF_0_n7), .A(stateFF_state_gff_16_SFF_0_n10), 
        .ZN(stateFF_state_gff_16_SFF_0_n6) );
  OAI221_X1 stateFF_state_gff_16_SFF_0_U3 ( .B1(stateFF_state_gff_16_n2), .B2(
        stateFF_inputPar[15]), .C1(stateFF_state_gff_16_SFF_0_n9), .C2(
        stateFF_inputPar[60]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_16_SFF_0_n10) );
  INV_X1 stateFF_state_gff_16_SFF_0_U2 ( .A(stateFF_state_gff_16_n2), .ZN(
        stateFF_state_gff_16_SFF_0_n9) );
  DFF_X1 stateFF_state_gff_16_SFF_0_Cell_reg ( .D(
        stateFF_state_gff_16_SFF_0_n6), .CK(clk), .Q(state[0]), .QN(
        stateFF_state_gff_16_SFF_0_n7) );
  OAI21_X1 stateFF_state_gff_16_SFF_1_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_16_SFF_1_n7), .A(stateFF_state_gff_16_SFF_1_n10), 
        .ZN(stateFF_state_gff_16_SFF_1_n6) );
  OAI221_X1 stateFF_state_gff_16_SFF_1_U3 ( .B1(stateFF_state_gff_16_n2), .B2(
        stateFF_inputPar[31]), .C1(stateFF_state_gff_16_SFF_1_n9), .C2(
        stateFF_inputPar[61]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_16_SFF_1_n10) );
  INV_X1 stateFF_state_gff_16_SFF_1_U2 ( .A(stateFF_state_gff_16_n2), .ZN(
        stateFF_state_gff_16_SFF_1_n9) );
  DFF_X1 stateFF_state_gff_16_SFF_1_Cell_reg ( .D(
        stateFF_state_gff_16_SFF_1_n6), .CK(clk), .Q(state[1]), .QN(
        stateFF_state_gff_16_SFF_1_n7) );
  OAI21_X1 stateFF_state_gff_16_SFF_2_U4 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_16_SFF_2_n7), .A(stateFF_state_gff_16_SFF_2_n10), 
        .ZN(stateFF_state_gff_16_SFF_2_n6) );
  OAI221_X1 stateFF_state_gff_16_SFF_2_U3 ( .B1(stateFF_state_gff_16_n2), .B2(
        stateFF_inputPar[47]), .C1(stateFF_state_gff_16_SFF_2_n9), .C2(
        stateFF_inputPar[62]), .A(stateFF_state_n7), .ZN(
        stateFF_state_gff_16_SFF_2_n10) );
  INV_X1 stateFF_state_gff_16_SFF_2_U2 ( .A(stateFF_state_gff_16_n2), .ZN(
        stateFF_state_gff_16_SFF_2_n9) );
  DFF_X1 stateFF_state_gff_16_SFF_2_Cell_reg ( .D(
        stateFF_state_gff_16_SFF_2_n6), .CK(clk), .Q(state[2]), .QN(
        stateFF_state_gff_16_SFF_2_n7) );
  OAI21_X1 stateFF_state_gff_16_SFF_3_U3 ( .B1(stateFF_state_n7), .B2(
        stateFF_state_gff_16_SFF_3_n7), .A(stateFF_state_gff_16_SFF_3_n9), 
        .ZN(stateFF_state_gff_16_SFF_3_n6) );
  NAND2_X1 stateFF_state_gff_16_SFF_3_U2 ( .A1(stateFF_state_n7), .A2(
        stateFF_n[6]), .ZN(stateFF_state_gff_16_SFF_3_n9) );
  DFF_X1 stateFF_state_gff_16_SFF_3_Cell_reg ( .D(
        stateFF_state_gff_16_SFF_3_n6), .CK(clk), .Q(state[3]), .QN(
        stateFF_state_gff_16_SFF_3_n7) );
  MUX2_X1 md1FF_U5 ( .A(share2[2]), .B(dataIn2[2]), .S(selInit), .Z(
        md1FF_inputPar[32]) );
  MUX2_X1 md1FF_U4 ( .A(share2[1]), .B(dataIn2[1]), .S(selInit), .Z(
        md1FF_inputPar[16]) );
  MUX2_X1 md1FF_U3 ( .A(share2[0]), .B(dataIn2[0]), .S(selInit), .Z(md1FF_n3)
         );
  MUX2_X1 md1FF_U2 ( .A(share2[3]), .B(dataIn2[3]), .S(selInit), .Z(
        md1FF_inputPar[48]) );
  BUF_X1 md1FF_state_U7 ( .A(selP), .Z(md1FF_state_n11) );
  BUF_X1 md1FF_state_U6 ( .A(selP), .Z(md1FF_state_n12) );
  BUF_X1 md1FF_state_U5 ( .A(selP), .Z(md1FF_state_n10) );
  BUF_X2 md1FF_state_U4 ( .A(enKey), .Z(md1FF_state_n9) );
  BUF_X2 md1FF_state_U3 ( .A(enKey), .Z(md1FF_state_n8) );
  BUF_X2 md1FF_state_U2 ( .A(enKey), .Z(md1FF_state_n6) );
  BUF_X2 md1FF_state_U1 ( .A(enKey), .Z(md1FF_state_n7) );
  BUF_X1 md1FF_state_gff_1_U2 ( .A(selP), .Z(md1FF_state_gff_1_n2) );
  OAI21_X1 md1FF_state_gff_1_SFF_0_U3 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_1_SFF_0_n8), .A(md1FF_state_gff_1_SFF_0_n10), .ZN(
        md1FF_state_gff_1_SFF_0_n7) );
  NAND2_X1 md1FF_state_gff_1_SFF_0_U2 ( .A1(md1FF_state_n7), .A2(md1FF_n3), 
        .ZN(md1FF_state_gff_1_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_1_SFF_0_Cell_reg ( .D(md1FF_state_gff_1_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[1]), .QN(md1FF_state_gff_1_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_1_SFF_1_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_1_SFF_1_n8), .A(md1FF_state_gff_1_SFF_1_n11), .ZN(
        md1FF_state_gff_1_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_1_SFF_1_U3 ( .B1(md1FF_state_gff_1_n2), .B2(
        md1FF_inputPar[16]), .C1(md1FF_state_gff_1_SFF_1_n10), .C2(
        md1FF_inputPar[1]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_1_SFF_1_n11) );
  INV_X1 md1FF_state_gff_1_SFF_1_U2 ( .A(md1FF_state_gff_1_n2), .ZN(
        md1FF_state_gff_1_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_1_SFF_1_Cell_reg ( .D(md1FF_state_gff_1_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[17]), .QN(md1FF_state_gff_1_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_1_SFF_2_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_1_SFF_2_n8), .A(md1FF_state_gff_1_SFF_2_n11), .ZN(
        md1FF_state_gff_1_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_1_SFF_2_U3 ( .B1(md1FF_state_gff_1_n2), .B2(
        md1FF_inputPar[32]), .C1(md1FF_state_gff_1_SFF_2_n10), .C2(
        md1FF_inputPar[2]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_1_SFF_2_n11) );
  INV_X1 md1FF_state_gff_1_SFF_2_U2 ( .A(md1FF_state_gff_1_n2), .ZN(
        md1FF_state_gff_1_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_1_SFF_2_Cell_reg ( .D(md1FF_state_gff_1_SFF_2_n7), 
        .CK(clk), .Q(md1FF_inputPar[33]), .QN(md1FF_state_gff_1_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_1_SFF_3_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_1_SFF_3_n8), .A(md1FF_state_gff_1_SFF_3_n11), .ZN(
        md1FF_state_gff_1_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_1_SFF_3_U3 ( .B1(md1FF_state_gff_1_n2), .B2(
        md1FF_inputPar[48]), .C1(md1FF_state_gff_1_SFF_3_n10), .C2(
        md1FF_inputPar[3]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_1_SFF_3_n11) );
  INV_X1 md1FF_state_gff_1_SFF_3_U2 ( .A(md1FF_state_gff_1_n2), .ZN(
        md1FF_state_gff_1_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_1_SFF_3_Cell_reg ( .D(md1FF_state_gff_1_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[49]), .QN(md1FF_state_gff_1_SFF_3_n8) );
  OAI21_X1 md1FF_state_gff_2_SFF_0_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_2_SFF_0_n8), .A(md1FF_state_gff_2_SFF_0_n12), .ZN(
        md1FF_state_gff_2_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_2_SFF_0_U4 ( .B1(md1FF_state_gff_2_SFF_0_n10), 
        .B2(md1FF_inputPar[1]), .C1(md1FF_state_gff_2_SFF_0_n11), .C2(
        md1FF_inputPar[4]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_2_SFF_0_n12) );
  INV_X1 md1FF_state_gff_2_SFF_0_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_2_SFF_0_n11) );
  INV_X1 md1FF_state_gff_2_SFF_0_U2 ( .A(md1FF_state_gff_2_SFF_0_n11), .ZN(
        md1FF_state_gff_2_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_2_SFF_0_Cell_reg ( .D(md1FF_state_gff_2_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[2]), .QN(md1FF_state_gff_2_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_2_SFF_1_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_2_SFF_1_n8), .A(md1FF_state_gff_2_SFF_1_n12), .ZN(
        md1FF_state_gff_2_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_2_SFF_1_U4 ( .B1(md1FF_state_gff_2_SFF_1_n10), 
        .B2(md1FF_inputPar[17]), .C1(md1FF_state_gff_2_SFF_1_n11), .C2(
        md1FF_inputPar[5]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_2_SFF_1_n12) );
  INV_X1 md1FF_state_gff_2_SFF_1_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_2_SFF_1_n11) );
  INV_X1 md1FF_state_gff_2_SFF_1_U2 ( .A(md1FF_state_gff_2_SFF_1_n11), .ZN(
        md1FF_state_gff_2_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_2_SFF_1_Cell_reg ( .D(md1FF_state_gff_2_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[18]), .QN(md1FF_state_gff_2_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_2_SFF_2_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_2_SFF_2_n8), .A(md1FF_state_gff_2_SFF_2_n12), .ZN(
        md1FF_state_gff_2_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_2_SFF_2_U4 ( .B1(md1FF_state_gff_2_SFF_2_n10), 
        .B2(md1FF_inputPar[33]), .C1(md1FF_state_gff_2_SFF_2_n11), .C2(
        md1FF_inputPar[6]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_2_SFF_2_n12) );
  INV_X1 md1FF_state_gff_2_SFF_2_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_2_SFF_2_n11) );
  INV_X1 md1FF_state_gff_2_SFF_2_U2 ( .A(md1FF_state_gff_2_SFF_2_n11), .ZN(
        md1FF_state_gff_2_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_2_SFF_2_Cell_reg ( .D(md1FF_state_gff_2_SFF_2_n7), 
        .CK(clk), .Q(md1FF_inputPar[34]), .QN(md1FF_state_gff_2_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_2_SFF_3_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_2_SFF_3_n8), .A(md1FF_state_gff_2_SFF_3_n12), .ZN(
        md1FF_state_gff_2_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_2_SFF_3_U4 ( .B1(md1FF_state_gff_2_SFF_3_n10), 
        .B2(md1FF_inputPar[49]), .C1(md1FF_state_gff_2_SFF_3_n11), .C2(
        md1FF_inputPar[7]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_2_SFF_3_n12) );
  INV_X1 md1FF_state_gff_2_SFF_3_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_2_SFF_3_n11) );
  INV_X1 md1FF_state_gff_2_SFF_3_U2 ( .A(md1FF_state_gff_2_SFF_3_n11), .ZN(
        md1FF_state_gff_2_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_2_SFF_3_Cell_reg ( .D(md1FF_state_gff_2_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[50]), .QN(md1FF_state_gff_2_SFF_3_n8) );
  OAI21_X1 md1FF_state_gff_3_SFF_0_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_3_SFF_0_n8), .A(md1FF_state_gff_3_SFF_0_n12), .ZN(
        md1FF_state_gff_3_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_3_SFF_0_U4 ( .B1(md1FF_state_gff_3_SFF_0_n10), 
        .B2(md1FF_inputPar[2]), .C1(md1FF_state_gff_3_SFF_0_n11), .C2(
        md1FF_inputPar[8]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_3_SFF_0_n12) );
  INV_X1 md1FF_state_gff_3_SFF_0_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_3_SFF_0_n11) );
  INV_X1 md1FF_state_gff_3_SFF_0_U2 ( .A(md1FF_state_gff_3_SFF_0_n11), .ZN(
        md1FF_state_gff_3_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_3_SFF_0_Cell_reg ( .D(md1FF_state_gff_3_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[3]), .QN(md1FF_state_gff_3_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_3_SFF_1_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_3_SFF_1_n8), .A(md1FF_state_gff_3_SFF_1_n12), .ZN(
        md1FF_state_gff_3_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_3_SFF_1_U4 ( .B1(md1FF_state_gff_3_SFF_1_n10), 
        .B2(md1FF_inputPar[18]), .C1(md1FF_state_gff_3_SFF_1_n11), .C2(
        md1FF_inputPar[9]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_3_SFF_1_n12) );
  INV_X1 md1FF_state_gff_3_SFF_1_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_3_SFF_1_n11) );
  INV_X1 md1FF_state_gff_3_SFF_1_U2 ( .A(md1FF_state_gff_3_SFF_1_n11), .ZN(
        md1FF_state_gff_3_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_3_SFF_1_Cell_reg ( .D(md1FF_state_gff_3_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[19]), .QN(md1FF_state_gff_3_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_3_SFF_2_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_3_SFF_2_n7), .A(md1FF_state_gff_3_SFF_2_n11), .ZN(
        md1FF_state_gff_3_SFF_2_n6) );
  OAI221_X1 md1FF_state_gff_3_SFF_2_U4 ( .B1(md1FF_state_gff_3_SFF_2_n9), .B2(
        md1FF_inputPar[34]), .C1(md1FF_state_gff_3_SFF_2_n10), .C2(
        md1FF_inputPar[10]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_3_SFF_2_n11) );
  INV_X1 md1FF_state_gff_3_SFF_2_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_3_SFF_2_n10) );
  INV_X1 md1FF_state_gff_3_SFF_2_U2 ( .A(md1FF_state_gff_3_SFF_2_n10), .ZN(
        md1FF_state_gff_3_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_3_SFF_2_Cell_reg ( .D(md1FF_state_gff_3_SFF_2_n6), 
        .CK(clk), .Q(md1FF_inputPar[35]), .QN(md1FF_state_gff_3_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_3_SFF_3_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_3_SFF_3_n7), .A(md1FF_state_gff_3_SFF_3_n11), .ZN(
        md1FF_state_gff_3_SFF_3_n6) );
  OAI221_X1 md1FF_state_gff_3_SFF_3_U4 ( .B1(md1FF_state_gff_3_SFF_3_n9), .B2(
        md1FF_inputPar[50]), .C1(md1FF_state_gff_3_SFF_3_n10), .C2(
        md1FF_inputPar[11]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_3_SFF_3_n11) );
  INV_X1 md1FF_state_gff_3_SFF_3_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_3_SFF_3_n10) );
  INV_X1 md1FF_state_gff_3_SFF_3_U2 ( .A(md1FF_state_gff_3_SFF_3_n10), .ZN(
        md1FF_state_gff_3_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_3_SFF_3_Cell_reg ( .D(md1FF_state_gff_3_SFF_3_n6), 
        .CK(clk), .Q(md1FF_inputPar[51]), .QN(md1FF_state_gff_3_SFF_3_n7) );
  OAI21_X1 md1FF_state_gff_4_SFF_0_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_4_SFF_0_n7), .A(md1FF_state_gff_4_SFF_0_n11), .ZN(
        md1FF_state_gff_4_SFF_0_n6) );
  OAI221_X1 md1FF_state_gff_4_SFF_0_U4 ( .B1(md1FF_state_gff_4_SFF_0_n9), .B2(
        md1FF_inputPar[3]), .C1(md1FF_state_gff_4_SFF_0_n10), .C2(
        md1FF_inputPar[12]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_4_SFF_0_n11) );
  INV_X1 md1FF_state_gff_4_SFF_0_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_4_SFF_0_n10) );
  INV_X1 md1FF_state_gff_4_SFF_0_U2 ( .A(md1FF_state_gff_4_SFF_0_n10), .ZN(
        md1FF_state_gff_4_SFF_0_n9) );
  DFF_X1 md1FF_state_gff_4_SFF_0_Cell_reg ( .D(md1FF_state_gff_4_SFF_0_n6), 
        .CK(clk), .Q(md1FF_inputPar[4]), .QN(md1FF_state_gff_4_SFF_0_n7) );
  OAI21_X1 md1FF_state_gff_4_SFF_1_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_4_SFF_1_n7), .A(md1FF_state_gff_4_SFF_1_n11), .ZN(
        md1FF_state_gff_4_SFF_1_n6) );
  OAI221_X1 md1FF_state_gff_4_SFF_1_U4 ( .B1(md1FF_state_gff_4_SFF_1_n9), .B2(
        md1FF_inputPar[19]), .C1(md1FF_state_gff_4_SFF_1_n10), .C2(
        md1FF_inputPar[13]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_4_SFF_1_n11) );
  INV_X1 md1FF_state_gff_4_SFF_1_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_4_SFF_1_n10) );
  INV_X1 md1FF_state_gff_4_SFF_1_U2 ( .A(md1FF_state_gff_4_SFF_1_n10), .ZN(
        md1FF_state_gff_4_SFF_1_n9) );
  DFF_X1 md1FF_state_gff_4_SFF_1_Cell_reg ( .D(md1FF_state_gff_4_SFF_1_n6), 
        .CK(clk), .Q(md1FF_inputPar[20]), .QN(md1FF_state_gff_4_SFF_1_n7) );
  OAI21_X1 md1FF_state_gff_4_SFF_2_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_4_SFF_2_n7), .A(md1FF_state_gff_4_SFF_2_n11), .ZN(
        md1FF_state_gff_4_SFF_2_n6) );
  OAI221_X1 md1FF_state_gff_4_SFF_2_U4 ( .B1(md1FF_state_gff_4_SFF_2_n9), .B2(
        md1FF_inputPar[35]), .C1(md1FF_state_gff_4_SFF_2_n10), .C2(
        md1FF_inputPar[14]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_4_SFF_2_n11) );
  INV_X1 md1FF_state_gff_4_SFF_2_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_4_SFF_2_n10) );
  INV_X1 md1FF_state_gff_4_SFF_2_U2 ( .A(md1FF_state_gff_4_SFF_2_n10), .ZN(
        md1FF_state_gff_4_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_4_SFF_2_Cell_reg ( .D(md1FF_state_gff_4_SFF_2_n6), 
        .CK(clk), .Q(md1FF_inputPar[36]), .QN(md1FF_state_gff_4_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_4_SFF_3_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_4_SFF_3_n7), .A(md1FF_state_gff_4_SFF_3_n11), .ZN(
        md1FF_state_gff_4_SFF_3_n6) );
  OAI221_X1 md1FF_state_gff_4_SFF_3_U4 ( .B1(md1FF_state_gff_4_SFF_3_n9), .B2(
        md1FF_inputPar[51]), .C1(md1FF_state_gff_4_SFF_3_n10), .C2(
        md1FF_inputPar[15]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_4_SFF_3_n11) );
  INV_X1 md1FF_state_gff_4_SFF_3_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_4_SFF_3_n10) );
  INV_X1 md1FF_state_gff_4_SFF_3_U2 ( .A(md1FF_state_gff_4_SFF_3_n10), .ZN(
        md1FF_state_gff_4_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_4_SFF_3_Cell_reg ( .D(md1FF_state_gff_4_SFF_3_n6), 
        .CK(clk), .Q(md1FF_inputPar[52]), .QN(md1FF_state_gff_4_SFF_3_n7) );
  OAI21_X1 md1FF_state_gff_5_SFF_0_U5 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_5_SFF_0_n8), .A(md1FF_state_gff_5_SFF_0_n12), .ZN(
        md1FF_state_gff_5_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_5_SFF_0_U4 ( .B1(md1FF_state_gff_5_SFF_0_n10), 
        .B2(md1FF_inputPar[4]), .C1(md1FF_state_gff_5_SFF_0_n11), .C2(
        md1FF_inputPar[16]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_5_SFF_0_n12) );
  INV_X1 md1FF_state_gff_5_SFF_0_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_5_SFF_0_n11) );
  INV_X1 md1FF_state_gff_5_SFF_0_U2 ( .A(md1FF_state_gff_5_SFF_0_n11), .ZN(
        md1FF_state_gff_5_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_5_SFF_0_Cell_reg ( .D(md1FF_state_gff_5_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[5]), .QN(md1FF_state_gff_5_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_5_SFF_1_U5 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_5_SFF_1_n8), .A(md1FF_state_gff_5_SFF_1_n12), .ZN(
        md1FF_state_gff_5_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_5_SFF_1_U4 ( .B1(md1FF_state_gff_5_SFF_1_n10), 
        .B2(md1FF_inputPar[20]), .C1(md1FF_state_gff_5_SFF_1_n11), .C2(
        md1FF_inputPar[17]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_5_SFF_1_n12) );
  INV_X1 md1FF_state_gff_5_SFF_1_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_5_SFF_1_n11) );
  INV_X1 md1FF_state_gff_5_SFF_1_U2 ( .A(md1FF_state_gff_5_SFF_1_n11), .ZN(
        md1FF_state_gff_5_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_5_SFF_1_Cell_reg ( .D(md1FF_state_gff_5_SFF_1_n7), 
        .CK(clk), .Q(md1FF_n[56]), .QN(md1FF_state_gff_5_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_5_SFF_2_U5 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_5_SFF_2_n8), .A(md1FF_state_gff_5_SFF_2_n12), .ZN(
        md1FF_state_gff_5_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_5_SFF_2_U4 ( .B1(md1FF_state_gff_5_SFF_2_n10), 
        .B2(md1FF_inputPar[36]), .C1(md1FF_state_gff_5_SFF_2_n11), .C2(
        md1FF_inputPar[18]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_5_SFF_2_n12) );
  INV_X1 md1FF_state_gff_5_SFF_2_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_5_SFF_2_n11) );
  INV_X1 md1FF_state_gff_5_SFF_2_U2 ( .A(md1FF_state_gff_5_SFF_2_n11), .ZN(
        md1FF_state_gff_5_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_5_SFF_2_Cell_reg ( .D(md1FF_state_gff_5_SFF_2_n7), 
        .CK(clk), .Q(md1FF_inputPar[37]), .QN(md1FF_state_gff_5_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_5_SFF_3_U5 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_5_SFF_3_n8), .A(md1FF_state_gff_5_SFF_3_n12), .ZN(
        md1FF_state_gff_5_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_5_SFF_3_U4 ( .B1(md1FF_state_gff_5_SFF_3_n10), 
        .B2(md1FF_inputPar[52]), .C1(md1FF_state_gff_5_SFF_3_n11), .C2(
        md1FF_inputPar[19]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_5_SFF_3_n12) );
  INV_X1 md1FF_state_gff_5_SFF_3_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_5_SFF_3_n11) );
  INV_X1 md1FF_state_gff_5_SFF_3_U2 ( .A(md1FF_state_gff_5_SFF_3_n11), .ZN(
        md1FF_state_gff_5_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_5_SFF_3_Cell_reg ( .D(md1FF_state_gff_5_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[53]), .QN(md1FF_state_gff_5_SFF_3_n8) );
  BUF_X1 md1FF_state_gff_6_U2 ( .A(selP), .Z(md1FF_state_gff_6_n2) );
  OAI21_X1 md1FF_state_gff_6_SFF_0_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_6_SFF_0_n8), .A(md1FF_state_gff_6_SFF_0_n11), .ZN(
        md1FF_state_gff_6_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_6_SFF_0_U3 ( .B1(md1FF_state_gff_6_n2), .B2(
        md1FF_inputPar[5]), .C1(md1FF_state_gff_6_SFF_0_n10), .C2(
        md1FF_inputPar[20]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_6_SFF_0_n11) );
  INV_X1 md1FF_state_gff_6_SFF_0_U2 ( .A(md1FF_state_gff_6_n2), .ZN(
        md1FF_state_gff_6_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_6_SFF_0_Cell_reg ( .D(md1FF_state_gff_6_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[6]), .QN(md1FF_state_gff_6_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_6_SFF_1_U3 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_6_SFF_1_n8), .A(md1FF_state_gff_6_SFF_1_n10), .ZN(
        md1FF_state_gff_6_SFF_1_n7) );
  NAND2_X1 md1FF_state_gff_6_SFF_1_U2 ( .A1(md1FF_state_n7), .A2(md1FF_n[56]), 
        .ZN(md1FF_state_gff_6_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_6_SFF_1_Cell_reg ( .D(md1FF_state_gff_6_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[22]), .QN(md1FF_state_gff_6_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_6_SFF_2_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_6_SFF_2_n8), .A(md1FF_state_gff_6_SFF_2_n11), .ZN(
        md1FF_state_gff_6_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_6_SFF_2_U3 ( .B1(md1FF_state_gff_6_n2), .B2(
        md1FF_inputPar[37]), .C1(md1FF_state_gff_6_SFF_2_n10), .C2(
        md1FF_inputPar[22]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_6_SFF_2_n11) );
  INV_X1 md1FF_state_gff_6_SFF_2_U2 ( .A(md1FF_state_gff_6_n2), .ZN(
        md1FF_state_gff_6_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_6_SFF_2_Cell_reg ( .D(md1FF_state_gff_6_SFF_2_n7), 
        .CK(clk), .Q(md1FF_inputPar[38]), .QN(md1FF_state_gff_6_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_6_SFF_3_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_6_SFF_3_n8), .A(md1FF_state_gff_6_SFF_3_n11), .ZN(
        md1FF_state_gff_6_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_6_SFF_3_U3 ( .B1(md1FF_state_gff_6_n2), .B2(
        md1FF_inputPar[53]), .C1(md1FF_state_gff_6_SFF_3_n10), .C2(
        md1FF_inputPar[23]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_6_SFF_3_n11) );
  INV_X1 md1FF_state_gff_6_SFF_3_U2 ( .A(md1FF_state_gff_6_n2), .ZN(
        md1FF_state_gff_6_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_6_SFF_3_Cell_reg ( .D(md1FF_state_gff_6_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[54]), .QN(md1FF_state_gff_6_SFF_3_n8) );
  OAI21_X1 md1FF_state_gff_7_SFF_0_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_7_SFF_0_n8), .A(md1FF_state_gff_7_SFF_0_n11), .ZN(
        md1FF_state_gff_7_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_7_SFF_0_U3 ( .B1(md1FF_state_n10), .B2(
        md1FF_inputPar[6]), .C1(md1FF_state_gff_7_SFF_0_n10), .C2(
        md1FF_inputPar[24]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_7_SFF_0_n11) );
  INV_X1 md1FF_state_gff_7_SFF_0_U2 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_7_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_7_SFF_0_Cell_reg ( .D(md1FF_state_gff_7_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[7]), .QN(md1FF_state_gff_7_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_7_SFF_1_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_7_SFF_1_n8), .A(md1FF_state_gff_7_SFF_1_n11), .ZN(
        md1FF_state_gff_7_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_7_SFF_1_U3 ( .B1(md1FF_state_n10), .B2(
        md1FF_inputPar[22]), .C1(md1FF_state_gff_7_SFF_1_n10), .C2(
        md1FF_inputPar[25]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_7_SFF_1_n11) );
  INV_X1 md1FF_state_gff_7_SFF_1_U2 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_7_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_7_SFF_1_Cell_reg ( .D(md1FF_state_gff_7_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[23]), .QN(md1FF_state_gff_7_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_7_SFF_2_U5 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_7_SFF_2_n7), .A(md1FF_state_gff_7_SFF_2_n11), .ZN(
        md1FF_state_gff_7_SFF_2_n6) );
  OAI221_X1 md1FF_state_gff_7_SFF_2_U4 ( .B1(md1FF_state_gff_7_SFF_2_n9), .B2(
        md1FF_inputPar[38]), .C1(md1FF_state_gff_7_SFF_2_n10), .C2(
        md1FF_inputPar[26]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_7_SFF_2_n11) );
  INV_X1 md1FF_state_gff_7_SFF_2_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_7_SFF_2_n10) );
  INV_X1 md1FF_state_gff_7_SFF_2_U2 ( .A(md1FF_state_gff_7_SFF_2_n10), .ZN(
        md1FF_state_gff_7_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_7_SFF_2_Cell_reg ( .D(md1FF_state_gff_7_SFF_2_n6), 
        .CK(clk), .Q(md1FF_inputPar[39]), .QN(md1FF_state_gff_7_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_7_SFF_3_U5 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_7_SFF_3_n7), .A(md1FF_state_gff_7_SFF_3_n11), .ZN(
        md1FF_state_gff_7_SFF_3_n6) );
  OAI221_X1 md1FF_state_gff_7_SFF_3_U4 ( .B1(md1FF_state_gff_7_SFF_3_n9), .B2(
        md1FF_inputPar[54]), .C1(md1FF_state_gff_7_SFF_3_n10), .C2(
        md1FF_inputPar[27]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_7_SFF_3_n11) );
  INV_X1 md1FF_state_gff_7_SFF_3_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_7_SFF_3_n10) );
  INV_X1 md1FF_state_gff_7_SFF_3_U2 ( .A(md1FF_state_gff_7_SFF_3_n10), .ZN(
        md1FF_state_gff_7_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_7_SFF_3_Cell_reg ( .D(md1FF_state_gff_7_SFF_3_n6), 
        .CK(clk), .Q(md1FF_inputPar[55]), .QN(md1FF_state_gff_7_SFF_3_n7) );
  OAI21_X1 md1FF_state_gff_8_SFF_0_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_8_SFF_0_n7), .A(md1FF_state_gff_8_SFF_0_n11), .ZN(
        md1FF_state_gff_8_SFF_0_n6) );
  OAI221_X1 md1FF_state_gff_8_SFF_0_U4 ( .B1(md1FF_state_gff_8_SFF_0_n9), .B2(
        md1FF_inputPar[7]), .C1(md1FF_state_gff_8_SFF_0_n10), .C2(
        md1FF_inputPar[28]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_8_SFF_0_n11) );
  INV_X1 md1FF_state_gff_8_SFF_0_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_8_SFF_0_n10) );
  INV_X1 md1FF_state_gff_8_SFF_0_U2 ( .A(md1FF_state_gff_8_SFF_0_n10), .ZN(
        md1FF_state_gff_8_SFF_0_n9) );
  DFF_X1 md1FF_state_gff_8_SFF_0_Cell_reg ( .D(md1FF_state_gff_8_SFF_0_n6), 
        .CK(clk), .Q(md1FF_inputPar[8]), .QN(md1FF_state_gff_8_SFF_0_n7) );
  OAI21_X1 md1FF_state_gff_8_SFF_1_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_8_SFF_1_n7), .A(md1FF_state_gff_8_SFF_1_n11), .ZN(
        md1FF_state_gff_8_SFF_1_n6) );
  OAI221_X1 md1FF_state_gff_8_SFF_1_U4 ( .B1(md1FF_state_gff_8_SFF_1_n9), .B2(
        md1FF_inputPar[23]), .C1(md1FF_state_gff_8_SFF_1_n10), .C2(
        md1FF_inputPar[29]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_8_SFF_1_n11) );
  INV_X1 md1FF_state_gff_8_SFF_1_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_8_SFF_1_n10) );
  INV_X1 md1FF_state_gff_8_SFF_1_U2 ( .A(md1FF_state_gff_8_SFF_1_n10), .ZN(
        md1FF_state_gff_8_SFF_1_n9) );
  DFF_X1 md1FF_state_gff_8_SFF_1_Cell_reg ( .D(md1FF_state_gff_8_SFF_1_n6), 
        .CK(clk), .Q(md1FF_inputPar[24]), .QN(md1FF_state_gff_8_SFF_1_n7) );
  OAI21_X1 md1FF_state_gff_8_SFF_2_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_8_SFF_2_n7), .A(md1FF_state_gff_8_SFF_2_n11), .ZN(
        md1FF_state_gff_8_SFF_2_n6) );
  OAI221_X1 md1FF_state_gff_8_SFF_2_U4 ( .B1(md1FF_state_gff_8_SFF_2_n9), .B2(
        md1FF_inputPar[39]), .C1(md1FF_state_gff_8_SFF_2_n10), .C2(
        md1FF_inputPar[30]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_8_SFF_2_n11) );
  INV_X1 md1FF_state_gff_8_SFF_2_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_8_SFF_2_n10) );
  INV_X1 md1FF_state_gff_8_SFF_2_U2 ( .A(md1FF_state_gff_8_SFF_2_n10), .ZN(
        md1FF_state_gff_8_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_8_SFF_2_Cell_reg ( .D(md1FF_state_gff_8_SFF_2_n6), 
        .CK(clk), .Q(md1FF_inputPar[40]), .QN(md1FF_state_gff_8_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_8_SFF_3_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_8_SFF_3_n7), .A(md1FF_state_gff_8_SFF_3_n11), .ZN(
        md1FF_state_gff_8_SFF_3_n6) );
  OAI221_X1 md1FF_state_gff_8_SFF_3_U4 ( .B1(md1FF_state_gff_8_SFF_3_n9), .B2(
        md1FF_inputPar[55]), .C1(md1FF_state_gff_8_SFF_3_n10), .C2(
        md1FF_inputPar[31]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_8_SFF_3_n11) );
  INV_X1 md1FF_state_gff_8_SFF_3_U3 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_8_SFF_3_n10) );
  INV_X1 md1FF_state_gff_8_SFF_3_U2 ( .A(md1FF_state_gff_8_SFF_3_n10), .ZN(
        md1FF_state_gff_8_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_8_SFF_3_Cell_reg ( .D(md1FF_state_gff_8_SFF_3_n6), 
        .CK(clk), .Q(md1FF_inputPar[56]), .QN(md1FF_state_gff_8_SFF_3_n7) );
  OAI21_X1 md1FF_state_gff_9_SFF_0_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_9_SFF_0_n8), .A(md1FF_state_gff_9_SFF_0_n12), .ZN(
        md1FF_state_gff_9_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_9_SFF_0_U4 ( .B1(md1FF_state_gff_9_SFF_0_n10), 
        .B2(md1FF_inputPar[8]), .C1(md1FF_state_gff_9_SFF_0_n11), .C2(
        md1FF_inputPar[32]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_9_SFF_0_n12) );
  INV_X1 md1FF_state_gff_9_SFF_0_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_9_SFF_0_n11) );
  INV_X1 md1FF_state_gff_9_SFF_0_U2 ( .A(md1FF_state_gff_9_SFF_0_n11), .ZN(
        md1FF_state_gff_9_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_9_SFF_0_Cell_reg ( .D(md1FF_state_gff_9_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[9]), .QN(md1FF_state_gff_9_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_9_SFF_1_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_9_SFF_1_n8), .A(md1FF_state_gff_9_SFF_1_n12), .ZN(
        md1FF_state_gff_9_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_9_SFF_1_U4 ( .B1(md1FF_state_gff_9_SFF_1_n10), 
        .B2(md1FF_inputPar[24]), .C1(md1FF_state_gff_9_SFF_1_n11), .C2(
        md1FF_inputPar[33]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_9_SFF_1_n12) );
  INV_X1 md1FF_state_gff_9_SFF_1_U3 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_9_SFF_1_n11) );
  INV_X1 md1FF_state_gff_9_SFF_1_U2 ( .A(md1FF_state_gff_9_SFF_1_n11), .ZN(
        md1FF_state_gff_9_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_9_SFF_1_Cell_reg ( .D(md1FF_state_gff_9_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[25]), .QN(md1FF_state_gff_9_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_9_SFF_2_U4 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_9_SFF_2_n8), .A(md1FF_state_gff_9_SFF_2_n11), .ZN(
        md1FF_state_gff_9_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_9_SFF_2_U3 ( .B1(md1FF_state_n12), .B2(
        md1FF_inputPar[40]), .C1(md1FF_state_gff_9_SFF_2_n10), .C2(
        md1FF_inputPar[34]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_9_SFF_2_n11) );
  INV_X1 md1FF_state_gff_9_SFF_2_U2 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_9_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_9_SFF_2_Cell_reg ( .D(md1FF_state_gff_9_SFF_2_n7), 
        .CK(clk), .Q(md1FF_inputPar[41]), .QN(md1FF_state_gff_9_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_9_SFF_3_U4 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_9_SFF_3_n8), .A(md1FF_state_gff_9_SFF_3_n11), .ZN(
        md1FF_state_gff_9_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_9_SFF_3_U3 ( .B1(md1FF_state_n12), .B2(
        md1FF_inputPar[56]), .C1(md1FF_state_gff_9_SFF_3_n10), .C2(
        md1FF_inputPar[35]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_9_SFF_3_n11) );
  INV_X1 md1FF_state_gff_9_SFF_3_U2 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_9_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_9_SFF_3_Cell_reg ( .D(md1FF_state_gff_9_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[57]), .QN(md1FF_state_gff_9_SFF_3_n8) );
  OAI21_X1 md1FF_state_gff_10_SFF_0_U4 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_10_SFF_0_n8), .A(md1FF_state_gff_10_SFF_0_n11), .ZN(
        md1FF_state_gff_10_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_10_SFF_0_U3 ( .B1(md1FF_state_n12), .B2(
        md1FF_inputPar[9]), .C1(md1FF_state_gff_10_SFF_0_n10), .C2(
        md1FF_inputPar[36]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_10_SFF_0_n11) );
  INV_X1 md1FF_state_gff_10_SFF_0_U2 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_10_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_10_SFF_0_Cell_reg ( .D(md1FF_state_gff_10_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[10]), .QN(md1FF_state_gff_10_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_10_SFF_1_U4 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_10_SFF_1_n8), .A(md1FF_state_gff_10_SFF_1_n11), .ZN(
        md1FF_state_gff_10_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_10_SFF_1_U3 ( .B1(md1FF_state_n12), .B2(
        md1FF_inputPar[25]), .C1(md1FF_state_gff_10_SFF_1_n10), .C2(
        md1FF_inputPar[37]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_10_SFF_1_n11) );
  INV_X1 md1FF_state_gff_10_SFF_1_U2 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_10_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_10_SFF_1_Cell_reg ( .D(md1FF_state_gff_10_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[26]), .QN(md1FF_state_gff_10_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_10_SFF_2_U4 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_10_SFF_2_n8), .A(md1FF_state_gff_10_SFF_2_n11), .ZN(
        md1FF_state_gff_10_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_10_SFF_2_U3 ( .B1(md1FF_state_n12), .B2(
        md1FF_inputPar[41]), .C1(md1FF_state_gff_10_SFF_2_n10), .C2(
        md1FF_inputPar[38]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_10_SFF_2_n11) );
  INV_X1 md1FF_state_gff_10_SFF_2_U2 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_10_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_10_SFF_2_Cell_reg ( .D(md1FF_state_gff_10_SFF_2_n7), 
        .CK(clk), .Q(md1FF_n[35]), .QN(md1FF_state_gff_10_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_10_SFF_3_U4 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_10_SFF_3_n8), .A(md1FF_state_gff_10_SFF_3_n11), .ZN(
        md1FF_state_gff_10_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_10_SFF_3_U3 ( .B1(md1FF_state_n12), .B2(
        md1FF_inputPar[57]), .C1(md1FF_state_gff_10_SFF_3_n10), .C2(
        md1FF_inputPar[39]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_10_SFF_3_n11) );
  INV_X1 md1FF_state_gff_10_SFF_3_U2 ( .A(md1FF_state_n12), .ZN(
        md1FF_state_gff_10_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_10_SFF_3_Cell_reg ( .D(md1FF_state_gff_10_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[58]), .QN(md1FF_state_gff_10_SFF_3_n8) );
  BUF_X1 md1FF_state_gff_11_U2 ( .A(md1FF_state_n11), .Z(md1FF_state_gff_11_n2) );
  OAI21_X1 md1FF_state_gff_11_SFF_0_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_11_SFF_0_n8), .A(md1FF_state_gff_11_SFF_0_n11), .ZN(
        md1FF_state_gff_11_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_11_SFF_0_U3 ( .B1(md1FF_state_gff_11_n2), .B2(
        md1FF_inputPar[10]), .C1(md1FF_state_gff_11_SFF_0_n10), .C2(
        md1FF_inputPar[40]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_11_SFF_0_n11) );
  INV_X1 md1FF_state_gff_11_SFF_0_U2 ( .A(md1FF_state_gff_11_n2), .ZN(
        md1FF_state_gff_11_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_11_SFF_0_Cell_reg ( .D(md1FF_state_gff_11_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[11]), .QN(md1FF_state_gff_11_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_11_SFF_1_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_11_SFF_1_n8), .A(md1FF_state_gff_11_SFF_1_n11), .ZN(
        md1FF_state_gff_11_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_11_SFF_1_U3 ( .B1(md1FF_state_gff_11_n2), .B2(
        md1FF_inputPar[26]), .C1(md1FF_state_gff_11_SFF_1_n10), .C2(
        md1FF_inputPar[41]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_11_SFF_1_n11) );
  INV_X1 md1FF_state_gff_11_SFF_1_U2 ( .A(md1FF_state_gff_11_n2), .ZN(
        md1FF_state_gff_11_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_11_SFF_1_Cell_reg ( .D(md1FF_state_gff_11_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[27]), .QN(md1FF_state_gff_11_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_11_SFF_2_U3 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_11_SFF_2_n7), .A(md1FF_state_gff_11_SFF_2_n9), .ZN(
        md1FF_state_gff_11_SFF_2_n6) );
  NAND2_X1 md1FF_state_gff_11_SFF_2_U2 ( .A1(md1FF_state_n7), .A2(md1FF_n[35]), 
        .ZN(md1FF_state_gff_11_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_11_SFF_2_Cell_reg ( .D(md1FF_state_gff_11_SFF_2_n6), 
        .CK(clk), .Q(md1FF_inputPar[43]), .QN(md1FF_state_gff_11_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_11_SFF_3_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_11_SFF_3_n7), .A(md1FF_state_gff_11_SFF_3_n10), .ZN(
        md1FF_state_gff_11_SFF_3_n6) );
  OAI221_X1 md1FF_state_gff_11_SFF_3_U3 ( .B1(md1FF_state_gff_11_n2), .B2(
        md1FF_inputPar[58]), .C1(md1FF_state_gff_11_SFF_3_n9), .C2(
        md1FF_inputPar[43]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_11_SFF_3_n10) );
  INV_X1 md1FF_state_gff_11_SFF_3_U2 ( .A(md1FF_state_gff_11_n2), .ZN(
        md1FF_state_gff_11_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_11_SFF_3_Cell_reg ( .D(md1FF_state_gff_11_SFF_3_n6), 
        .CK(clk), .Q(md1FF_inputPar[59]), .QN(md1FF_state_gff_11_SFF_3_n7) );
  OAI21_X1 md1FF_state_gff_12_SFF_0_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_12_SFF_0_n7), .A(md1FF_state_gff_12_SFF_0_n10), .ZN(
        md1FF_state_gff_12_SFF_0_n6) );
  OAI221_X1 md1FF_state_gff_12_SFF_0_U3 ( .B1(md1FF_state_n10), .B2(
        md1FF_inputPar[11]), .C1(md1FF_state_gff_12_SFF_0_n9), .C2(
        md1FF_inputPar[44]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_12_SFF_0_n10) );
  INV_X1 md1FF_state_gff_12_SFF_0_U2 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_12_SFF_0_n9) );
  DFF_X1 md1FF_state_gff_12_SFF_0_Cell_reg ( .D(md1FF_state_gff_12_SFF_0_n6), 
        .CK(clk), .Q(md1FF_inputPar[12]), .QN(md1FF_state_gff_12_SFF_0_n7) );
  OAI21_X1 md1FF_state_gff_12_SFF_1_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_12_SFF_1_n7), .A(md1FF_state_gff_12_SFF_1_n10), .ZN(
        md1FF_state_gff_12_SFF_1_n6) );
  OAI221_X1 md1FF_state_gff_12_SFF_1_U3 ( .B1(md1FF_state_n10), .B2(
        md1FF_inputPar[27]), .C1(md1FF_state_gff_12_SFF_1_n9), .C2(
        md1FF_inputPar[45]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_12_SFF_1_n10) );
  INV_X1 md1FF_state_gff_12_SFF_1_U2 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_12_SFF_1_n9) );
  DFF_X1 md1FF_state_gff_12_SFF_1_Cell_reg ( .D(md1FF_state_gff_12_SFF_1_n6), 
        .CK(clk), .Q(md1FF_inputPar[28]), .QN(md1FF_state_gff_12_SFF_1_n7) );
  OAI21_X1 md1FF_state_gff_12_SFF_2_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_12_SFF_2_n7), .A(md1FF_state_gff_12_SFF_2_n10), .ZN(
        md1FF_state_gff_12_SFF_2_n6) );
  OAI221_X1 md1FF_state_gff_12_SFF_2_U3 ( .B1(md1FF_state_n10), .B2(
        md1FF_inputPar[43]), .C1(md1FF_state_gff_12_SFF_2_n9), .C2(
        md1FF_inputPar[46]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_12_SFF_2_n10) );
  INV_X1 md1FF_state_gff_12_SFF_2_U2 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_12_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_12_SFF_2_Cell_reg ( .D(md1FF_state_gff_12_SFF_2_n6), 
        .CK(clk), .Q(md1FF_inputPar[44]), .QN(md1FF_state_gff_12_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_12_SFF_3_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_12_SFF_3_n7), .A(md1FF_state_gff_12_SFF_3_n10), .ZN(
        md1FF_state_gff_12_SFF_3_n6) );
  OAI221_X1 md1FF_state_gff_12_SFF_3_U3 ( .B1(md1FF_state_n10), .B2(
        md1FF_inputPar[59]), .C1(md1FF_state_gff_12_SFF_3_n9), .C2(
        md1FF_inputPar[47]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_12_SFF_3_n10) );
  INV_X1 md1FF_state_gff_12_SFF_3_U2 ( .A(md1FF_state_n10), .ZN(
        md1FF_state_gff_12_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_12_SFF_3_Cell_reg ( .D(md1FF_state_gff_12_SFF_3_n6), 
        .CK(clk), .Q(md1FF_inputPar[60]), .QN(md1FF_state_gff_12_SFF_3_n7) );
  OAI21_X1 md1FF_state_gff_13_SFF_0_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_13_SFF_0_n8), .A(md1FF_state_gff_13_SFF_0_n12), .ZN(
        md1FF_state_gff_13_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_13_SFF_0_U4 ( .B1(md1FF_state_gff_13_SFF_0_n10), 
        .B2(md1FF_inputPar[12]), .C1(md1FF_state_gff_13_SFF_0_n11), .C2(
        md1FF_inputPar[48]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_13_SFF_0_n12) );
  INV_X1 md1FF_state_gff_13_SFF_0_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_13_SFF_0_n11) );
  INV_X1 md1FF_state_gff_13_SFF_0_U2 ( .A(md1FF_state_gff_13_SFF_0_n11), .ZN(
        md1FF_state_gff_13_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_13_SFF_0_Cell_reg ( .D(md1FF_state_gff_13_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[13]), .QN(md1FF_state_gff_13_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_13_SFF_1_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_13_SFF_1_n8), .A(md1FF_state_gff_13_SFF_1_n12), .ZN(
        md1FF_state_gff_13_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_13_SFF_1_U4 ( .B1(md1FF_state_gff_13_SFF_1_n10), 
        .B2(md1FF_inputPar[28]), .C1(md1FF_state_gff_13_SFF_1_n11), .C2(
        md1FF_inputPar[49]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_13_SFF_1_n12) );
  INV_X1 md1FF_state_gff_13_SFF_1_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_13_SFF_1_n11) );
  INV_X1 md1FF_state_gff_13_SFF_1_U2 ( .A(md1FF_state_gff_13_SFF_1_n11), .ZN(
        md1FF_state_gff_13_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_13_SFF_1_Cell_reg ( .D(md1FF_state_gff_13_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[29]), .QN(md1FF_state_gff_13_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_13_SFF_2_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_13_SFF_2_n8), .A(md1FF_state_gff_13_SFF_2_n12), .ZN(
        md1FF_state_gff_13_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_13_SFF_2_U4 ( .B1(md1FF_state_gff_13_SFF_2_n10), 
        .B2(md1FF_inputPar[44]), .C1(md1FF_state_gff_13_SFF_2_n11), .C2(
        md1FF_inputPar[50]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_13_SFF_2_n12) );
  INV_X1 md1FF_state_gff_13_SFF_2_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_13_SFF_2_n11) );
  INV_X1 md1FF_state_gff_13_SFF_2_U2 ( .A(md1FF_state_gff_13_SFF_2_n11), .ZN(
        md1FF_state_gff_13_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_13_SFF_2_Cell_reg ( .D(md1FF_state_gff_13_SFF_2_n7), 
        .CK(clk), .Q(md1FF_inputPar[45]), .QN(md1FF_state_gff_13_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_13_SFF_3_U5 ( .B1(md1FF_state_n6), .B2(
        md1FF_state_gff_13_SFF_3_n8), .A(md1FF_state_gff_13_SFF_3_n12), .ZN(
        md1FF_state_gff_13_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_13_SFF_3_U4 ( .B1(md1FF_state_gff_13_SFF_3_n10), 
        .B2(md1FF_inputPar[60]), .C1(md1FF_state_gff_13_SFF_3_n11), .C2(
        md1FF_inputPar[51]), .A(md1FF_state_n6), .ZN(
        md1FF_state_gff_13_SFF_3_n12) );
  INV_X1 md1FF_state_gff_13_SFF_3_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_13_SFF_3_n11) );
  INV_X1 md1FF_state_gff_13_SFF_3_U2 ( .A(md1FF_state_gff_13_SFF_3_n11), .ZN(
        md1FF_state_gff_13_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_13_SFF_3_Cell_reg ( .D(md1FF_state_gff_13_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[61]), .QN(md1FF_state_gff_13_SFF_3_n8) );
  OAI21_X1 md1FF_state_gff_14_SFF_0_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_14_SFF_0_n8), .A(md1FF_state_gff_14_SFF_0_n11), .ZN(
        md1FF_state_gff_14_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_14_SFF_0_U3 ( .B1(md1FF_state_n11), .B2(
        md1FF_inputPar[13]), .C1(md1FF_state_gff_14_SFF_0_n10), .C2(
        md1FF_inputPar[52]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_14_SFF_0_n11) );
  INV_X1 md1FF_state_gff_14_SFF_0_U2 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_14_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_14_SFF_0_Cell_reg ( .D(md1FF_state_gff_14_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[14]), .QN(md1FF_state_gff_14_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_14_SFF_1_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_14_SFF_1_n8), .A(md1FF_state_gff_14_SFF_1_n11), .ZN(
        md1FF_state_gff_14_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_14_SFF_1_U3 ( .B1(md1FF_state_n11), .B2(
        md1FF_inputPar[29]), .C1(md1FF_state_gff_14_SFF_1_n10), .C2(
        md1FF_inputPar[53]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_14_SFF_1_n11) );
  INV_X1 md1FF_state_gff_14_SFF_1_U2 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_14_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_14_SFF_1_Cell_reg ( .D(md1FF_state_gff_14_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[30]), .QN(md1FF_state_gff_14_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_14_SFF_2_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_14_SFF_2_n8), .A(md1FF_state_gff_14_SFF_2_n11), .ZN(
        md1FF_state_gff_14_SFF_2_n7) );
  OAI221_X1 md1FF_state_gff_14_SFF_2_U3 ( .B1(md1FF_state_n11), .B2(
        md1FF_inputPar[45]), .C1(md1FF_state_gff_14_SFF_2_n10), .C2(
        md1FF_inputPar[54]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_14_SFF_2_n11) );
  INV_X1 md1FF_state_gff_14_SFF_2_U2 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_14_SFF_2_n10) );
  DFF_X1 md1FF_state_gff_14_SFF_2_Cell_reg ( .D(md1FF_state_gff_14_SFF_2_n7), 
        .CK(clk), .Q(md1FF_inputPar[46]), .QN(md1FF_state_gff_14_SFF_2_n8) );
  OAI21_X1 md1FF_state_gff_14_SFF_3_U4 ( .B1(md1FF_state_n8), .B2(
        md1FF_state_gff_14_SFF_3_n8), .A(md1FF_state_gff_14_SFF_3_n11), .ZN(
        md1FF_state_gff_14_SFF_3_n7) );
  OAI221_X1 md1FF_state_gff_14_SFF_3_U3 ( .B1(md1FF_state_n11), .B2(
        md1FF_inputPar[61]), .C1(md1FF_state_gff_14_SFF_3_n10), .C2(
        md1FF_inputPar[55]), .A(md1FF_state_n8), .ZN(
        md1FF_state_gff_14_SFF_3_n11) );
  INV_X1 md1FF_state_gff_14_SFF_3_U2 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_14_SFF_3_n10) );
  DFF_X1 md1FF_state_gff_14_SFF_3_Cell_reg ( .D(md1FF_state_gff_14_SFF_3_n7), 
        .CK(clk), .Q(md1FF_inputPar[62]), .QN(md1FF_state_gff_14_SFF_3_n8) );
  OAI21_X1 md1FF_state_gff_15_SFF_0_U4 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_15_SFF_0_n8), .A(md1FF_state_gff_15_SFF_0_n11), .ZN(
        md1FF_state_gff_15_SFF_0_n7) );
  OAI221_X1 md1FF_state_gff_15_SFF_0_U3 ( .B1(md1FF_state_n11), .B2(
        md1FF_inputPar[14]), .C1(md1FF_state_gff_15_SFF_0_n10), .C2(
        md1FF_inputPar[56]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_15_SFF_0_n11) );
  INV_X1 md1FF_state_gff_15_SFF_0_U2 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_15_SFF_0_n10) );
  DFF_X1 md1FF_state_gff_15_SFF_0_Cell_reg ( .D(md1FF_state_gff_15_SFF_0_n7), 
        .CK(clk), .Q(md1FF_inputPar[15]), .QN(md1FF_state_gff_15_SFF_0_n8) );
  OAI21_X1 md1FF_state_gff_15_SFF_1_U4 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_15_SFF_1_n8), .A(md1FF_state_gff_15_SFF_1_n11), .ZN(
        md1FF_state_gff_15_SFF_1_n7) );
  OAI221_X1 md1FF_state_gff_15_SFF_1_U3 ( .B1(md1FF_state_n11), .B2(
        md1FF_inputPar[30]), .C1(md1FF_state_gff_15_SFF_1_n10), .C2(
        md1FF_inputPar[57]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_15_SFF_1_n11) );
  INV_X1 md1FF_state_gff_15_SFF_1_U2 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_15_SFF_1_n10) );
  DFF_X1 md1FF_state_gff_15_SFF_1_Cell_reg ( .D(md1FF_state_gff_15_SFF_1_n7), 
        .CK(clk), .Q(md1FF_inputPar[31]), .QN(md1FF_state_gff_15_SFF_1_n8) );
  OAI21_X1 md1FF_state_gff_15_SFF_2_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_15_SFF_2_n7), .A(md1FF_state_gff_15_SFF_2_n11), .ZN(
        md1FF_state_gff_15_SFF_2_n6) );
  OAI221_X1 md1FF_state_gff_15_SFF_2_U4 ( .B1(md1FF_state_gff_15_SFF_2_n9), 
        .B2(md1FF_inputPar[46]), .C1(md1FF_state_gff_15_SFF_2_n10), .C2(
        md1FF_inputPar[58]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_15_SFF_2_n11) );
  INV_X1 md1FF_state_gff_15_SFF_2_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_15_SFF_2_n10) );
  INV_X1 md1FF_state_gff_15_SFF_2_U2 ( .A(md1FF_state_gff_15_SFF_2_n10), .ZN(
        md1FF_state_gff_15_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_15_SFF_2_Cell_reg ( .D(md1FF_state_gff_15_SFF_2_n6), 
        .CK(clk), .Q(md1FF_inputPar[47]), .QN(md1FF_state_gff_15_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_15_SFF_3_U5 ( .B1(md1FF_state_n9), .B2(
        md1FF_state_gff_15_SFF_3_n7), .A(md1FF_state_gff_15_SFF_3_n11), .ZN(
        md1FF_state_gff_15_SFF_3_n6) );
  OAI221_X1 md1FF_state_gff_15_SFF_3_U4 ( .B1(md1FF_state_gff_15_SFF_3_n9), 
        .B2(md1FF_inputPar[62]), .C1(md1FF_state_gff_15_SFF_3_n10), .C2(
        md1FF_inputPar[59]), .A(md1FF_state_n9), .ZN(
        md1FF_state_gff_15_SFF_3_n11) );
  INV_X1 md1FF_state_gff_15_SFF_3_U3 ( .A(md1FF_state_n11), .ZN(
        md1FF_state_gff_15_SFF_3_n10) );
  INV_X1 md1FF_state_gff_15_SFF_3_U2 ( .A(md1FF_state_gff_15_SFF_3_n10), .ZN(
        md1FF_state_gff_15_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_15_SFF_3_Cell_reg ( .D(md1FF_state_gff_15_SFF_3_n6), 
        .CK(clk), .Q(md1FF_n[14]), .QN(md1FF_state_gff_15_SFF_3_n7) );
  BUF_X1 md1FF_state_gff_16_U2 ( .A(md1FF_state_n12), .Z(md1FF_state_gff_16_n2) );
  OAI21_X1 md1FF_state_gff_16_SFF_0_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_16_SFF_0_n7), .A(md1FF_state_gff_16_SFF_0_n10), .ZN(
        md1FF_state_gff_16_SFF_0_n6) );
  OAI221_X1 md1FF_state_gff_16_SFF_0_U3 ( .B1(md1FF_state_gff_16_n2), .B2(
        md1FF_inputPar[15]), .C1(md1FF_state_gff_16_SFF_0_n9), .C2(
        md1FF_inputPar[60]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_16_SFF_0_n10) );
  INV_X1 md1FF_state_gff_16_SFF_0_U2 ( .A(md1FF_state_gff_16_n2), .ZN(
        md1FF_state_gff_16_SFF_0_n9) );
  DFF_X1 md1FF_state_gff_16_SFF_0_Cell_reg ( .D(md1FF_state_gff_16_SFF_0_n6), 
        .CK(clk), .Q(dataOut2[0]), .QN(md1FF_state_gff_16_SFF_0_n7) );
  OAI21_X1 md1FF_state_gff_16_SFF_1_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_16_SFF_1_n7), .A(md1FF_state_gff_16_SFF_1_n10), .ZN(
        md1FF_state_gff_16_SFF_1_n6) );
  OAI221_X1 md1FF_state_gff_16_SFF_1_U3 ( .B1(md1FF_state_gff_16_n2), .B2(
        md1FF_inputPar[31]), .C1(md1FF_state_gff_16_SFF_1_n9), .C2(
        md1FF_inputPar[61]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_16_SFF_1_n10) );
  INV_X1 md1FF_state_gff_16_SFF_1_U2 ( .A(md1FF_state_gff_16_n2), .ZN(
        md1FF_state_gff_16_SFF_1_n9) );
  DFF_X1 md1FF_state_gff_16_SFF_1_Cell_reg ( .D(md1FF_state_gff_16_SFF_1_n6), 
        .CK(clk), .Q(dataOut2[1]), .QN(md1FF_state_gff_16_SFF_1_n7) );
  OAI21_X1 md1FF_state_gff_16_SFF_2_U4 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_16_SFF_2_n7), .A(md1FF_state_gff_16_SFF_2_n10), .ZN(
        md1FF_state_gff_16_SFF_2_n6) );
  OAI221_X1 md1FF_state_gff_16_SFF_2_U3 ( .B1(md1FF_state_gff_16_n2), .B2(
        md1FF_inputPar[47]), .C1(md1FF_state_gff_16_SFF_2_n9), .C2(
        md1FF_inputPar[62]), .A(md1FF_state_n7), .ZN(
        md1FF_state_gff_16_SFF_2_n10) );
  INV_X1 md1FF_state_gff_16_SFF_2_U2 ( .A(md1FF_state_gff_16_n2), .ZN(
        md1FF_state_gff_16_SFF_2_n9) );
  DFF_X1 md1FF_state_gff_16_SFF_2_Cell_reg ( .D(md1FF_state_gff_16_SFF_2_n6), 
        .CK(clk), .Q(dataOut2[2]), .QN(md1FF_state_gff_16_SFF_2_n7) );
  OAI21_X1 md1FF_state_gff_16_SFF_3_U3 ( .B1(md1FF_state_n7), .B2(
        md1FF_state_gff_16_SFF_3_n7), .A(md1FF_state_gff_16_SFF_3_n9), .ZN(
        md1FF_state_gff_16_SFF_3_n6) );
  NAND2_X1 md1FF_state_gff_16_SFF_3_U2 ( .A1(md1FF_state_n7), .A2(md1FF_n[14]), 
        .ZN(md1FF_state_gff_16_SFF_3_n9) );
  DFF_X1 md1FF_state_gff_16_SFF_3_Cell_reg ( .D(md1FF_state_gff_16_SFF_3_n6), 
        .CK(clk), .Q(dataOut2[3]), .QN(md1FF_state_gff_16_SFF_3_n7) );
  MUX2_X1 keyFF_U10 ( .A(roundkey[0]), .B(key[0]), .S(selInit), .Z(keyFF_n1)
         );
  MUX2_X1 keyFF_U9 ( .A(roundkey[1]), .B(key[1]), .S(selInit), .Z(keyFF_n2) );
  MUX2_X1 keyFF_U8 ( .A(roundkey[2]), .B(key[2]), .S(selInit), .Z(keyFF_n3) );
  MUX2_X1 keyFF_U7 ( .A(roundkey[3]), .B(key[3]), .S(selInit), .Z(keyFF_n4) );
  XOR2_X1 keyFF_U6 ( .A(counter[4]), .B(keyFF_outputPar[22]), .Z(
        keyFF_counterAdd[4]) );
  XOR2_X1 keyFF_U5 ( .A(counter[3]), .B(keyFF_outputPar[21]), .Z(
        keyFF_counterAdd[3]) );
  XOR2_X1 keyFF_U4 ( .A(counter[2]), .B(keyFF_outputPar[20]), .Z(
        keyFF_counterAdd[2]) );
  XOR2_X1 keyFF_U3 ( .A(counter[1]), .B(keyFF_outputPar[19]), .Z(
        keyFF_counterAdd[1]) );
  XOR2_X1 keyFF_U2 ( .A(counter[0]), .B(keyFF_outputPar[18]), .Z(
        keyFF_counterAdd[0]) );
  BUF_X2 keyFF_keystate_U9 ( .A(enKey), .Z(keyFF_keystate_n13) );
  BUF_X2 keyFF_keystate_U8 ( .A(enKey), .Z(keyFF_keystate_n12) );
  BUF_X2 keyFF_keystate_U7 ( .A(enKey), .Z(keyFF_keystate_n11) );
  BUF_X2 keyFF_keystate_U6 ( .A(enKey), .Z(keyFF_keystate_n10) );
  BUF_X1 keyFF_keystate_U5 ( .A(selP), .Z(keyFF_keystate_n18) );
  BUF_X1 keyFF_keystate_U4 ( .A(selP), .Z(keyFF_keystate_n17) );
  BUF_X1 keyFF_keystate_U3 ( .A(selP), .Z(keyFF_keystate_n16) );
  BUF_X1 keyFF_keystate_U2 ( .A(selP), .Z(keyFF_keystate_n15) );
  BUF_X1 keyFF_keystate_U1 ( .A(selP), .Z(keyFF_keystate_n14) );
  OAI21_X1 keyFF_keystate_gff_1_SFF_0_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_1_SFF_0_n8), .A(keyFF_keystate_gff_1_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_1_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_1_SFF_0_U4 ( .B1(keyFF_keystate_gff_1_SFF_0_n10), .B2(keyFF_n1), .C1(keyFF_keystate_gff_1_SFF_0_n11), .C2(keyFF_outputPar[3]), 
        .A(keyFF_keystate_n10), .ZN(keyFF_keystate_gff_1_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_1_SFF_0_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_1_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_1_SFF_0_U2 ( .A(keyFF_keystate_gff_1_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_1_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_1_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_1_SFF_0_n7), .CK(clk), .Q(keyRegKS[1]), .QN(
        keyFF_keystate_gff_1_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_1_SFF_1_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_1_SFF_1_n8), .A(keyFF_keystate_gff_1_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_1_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_1_SFF_1_U4 ( .B1(keyFF_keystate_gff_1_SFF_1_n10), .B2(keyFF_n2), .C1(keyFF_keystate_gff_1_SFF_1_n11), .C2(keyFF_outputPar[4]), 
        .A(keyFF_keystate_n10), .ZN(keyFF_keystate_gff_1_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_1_SFF_1_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_1_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_1_SFF_1_U2 ( .A(keyFF_keystate_gff_1_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_1_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_1_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_1_SFF_1_n7), .CK(clk), .Q(keyRegKS[2]), .QN(
        keyFF_keystate_gff_1_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_1_SFF_2_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_1_SFF_2_n8), .A(keyFF_keystate_gff_1_SFF_2_n12), 
        .ZN(keyFF_keystate_gff_1_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_1_SFF_2_U4 ( .B1(keyFF_keystate_gff_1_SFF_2_n10), .B2(keyFF_n3), .C1(keyFF_keystate_gff_1_SFF_2_n11), .C2(keyFF_outputPar[5]), 
        .A(keyFF_keystate_n10), .ZN(keyFF_keystate_gff_1_SFF_2_n12) );
  INV_X1 keyFF_keystate_gff_1_SFF_2_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_1_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_1_SFF_2_U2 ( .A(keyFF_keystate_gff_1_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_1_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_1_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_1_SFF_2_n7), .CK(clk), .Q(keyRegKS[3]), .QN(
        keyFF_keystate_gff_1_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_1_SFF_3_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_1_SFF_3_n8), .A(keyFF_keystate_gff_1_SFF_3_n12), 
        .ZN(keyFF_keystate_gff_1_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_1_SFF_3_U4 ( .B1(keyFF_keystate_gff_1_SFF_3_n10), .B2(keyFF_n4), .C1(keyFF_keystate_gff_1_SFF_3_n11), .C2(keyFF_outputPar[6]), 
        .A(keyFF_keystate_n10), .ZN(keyFF_keystate_gff_1_SFF_3_n12) );
  INV_X1 keyFF_keystate_gff_1_SFF_3_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_1_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_1_SFF_3_U2 ( .A(keyFF_keystate_gff_1_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_1_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_1_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_1_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[3]), .QN(
        keyFF_keystate_gff_1_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_2_SFF_0_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_2_SFF_0_n8), .A(keyFF_keystate_gff_2_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_2_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_2_SFF_0_U4 ( .B1(keyFF_keystate_gff_2_SFF_0_n10), .B2(keyRegKS[1]), .C1(keyFF_keystate_gff_2_SFF_0_n11), .C2(
        keyFF_outputPar[7]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_2_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_2_SFF_0_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_2_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_2_SFF_0_U2 ( .A(keyFF_keystate_gff_2_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_2_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_2_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_2_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[4]), .QN(
        keyFF_keystate_gff_2_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_2_SFF_1_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_2_SFF_1_n8), .A(keyFF_keystate_gff_2_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_2_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_2_SFF_1_U4 ( .B1(keyFF_keystate_gff_2_SFF_1_n10), .B2(keyRegKS[2]), .C1(keyFF_keystate_gff_2_SFF_1_n11), .C2(
        keyFF_outputPar[8]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_2_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_2_SFF_1_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_2_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_2_SFF_1_U2 ( .A(keyFF_keystate_gff_2_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_2_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_2_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_2_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[5]), .QN(
        keyFF_keystate_gff_2_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_2_SFF_2_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_2_SFF_2_n8), .A(keyFF_keystate_gff_2_SFF_2_n12), 
        .ZN(keyFF_keystate_gff_2_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_2_SFF_2_U4 ( .B1(keyFF_keystate_gff_2_SFF_2_n10), .B2(keyRegKS[3]), .C1(keyFF_keystate_gff_2_SFF_2_n11), .C2(
        keyFF_outputPar[9]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_2_SFF_2_n12) );
  INV_X1 keyFF_keystate_gff_2_SFF_2_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_2_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_2_SFF_2_U2 ( .A(keyFF_keystate_gff_2_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_2_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_2_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_2_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[6]), .QN(
        keyFF_keystate_gff_2_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_2_SFF_3_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_2_SFF_3_n8), .A(keyFF_keystate_gff_2_SFF_3_n12), 
        .ZN(keyFF_keystate_gff_2_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_2_SFF_3_U4 ( .B1(keyFF_keystate_gff_2_SFF_3_n10), .B2(keyFF_outputPar[3]), .C1(keyFF_keystate_gff_2_SFF_3_n11), .C2(
        keyFF_outputPar[10]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_2_SFF_3_n12) );
  INV_X1 keyFF_keystate_gff_2_SFF_3_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_2_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_2_SFF_3_U2 ( .A(keyFF_keystate_gff_2_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_2_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_2_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_2_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[7]), .QN(
        keyFF_keystate_gff_2_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_3_SFF_0_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_3_SFF_0_n8), .A(keyFF_keystate_gff_3_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_3_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_3_SFF_0_U4 ( .B1(keyFF_keystate_gff_3_SFF_0_n10), .B2(keyFF_outputPar[4]), .C1(keyFF_keystate_gff_3_SFF_0_n11), .C2(
        keyFF_outputPar[11]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_3_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_3_SFF_0_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_3_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_3_SFF_0_U2 ( .A(keyFF_keystate_gff_3_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_3_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_3_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_3_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[8]), .QN(
        keyFF_keystate_gff_3_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_3_SFF_1_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_3_SFF_1_n8), .A(keyFF_keystate_gff_3_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_3_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_3_SFF_1_U4 ( .B1(keyFF_keystate_gff_3_SFF_1_n10), .B2(keyFF_outputPar[5]), .C1(keyFF_keystate_gff_3_SFF_1_n11), .C2(
        keyFF_outputPar[12]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_3_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_3_SFF_1_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_3_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_3_SFF_1_U2 ( .A(keyFF_keystate_gff_3_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_3_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_3_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_3_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[9]), .QN(
        keyFF_keystate_gff_3_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_3_SFF_2_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_3_SFF_2_n7), .A(keyFF_keystate_gff_3_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_3_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_3_SFF_2_U4 ( .B1(keyFF_keystate_gff_3_SFF_2_n9), 
        .B2(keyFF_outputPar[6]), .C1(keyFF_keystate_gff_3_SFF_2_n10), .C2(
        keyFF_outputPar[13]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_3_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_3_SFF_2_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_3_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_3_SFF_2_U2 ( .A(keyFF_keystate_gff_3_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_3_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_3_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_3_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[10]), 
        .QN(keyFF_keystate_gff_3_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_3_SFF_3_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_3_SFF_3_n7), .A(keyFF_keystate_gff_3_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_3_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_3_SFF_3_U4 ( .B1(keyFF_keystate_gff_3_SFF_3_n9), 
        .B2(keyFF_outputPar[7]), .C1(keyFF_keystate_gff_3_SFF_3_n10), .C2(
        keyFF_outputPar[14]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_3_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_3_SFF_3_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_3_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_3_SFF_3_U2 ( .A(keyFF_keystate_gff_3_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_3_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_3_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_3_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[11]), 
        .QN(keyFF_keystate_gff_3_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_4_SFF_0_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_4_SFF_0_n7), .A(keyFF_keystate_gff_4_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_4_SFF_0_n6) );
  OAI221_X1 keyFF_keystate_gff_4_SFF_0_U4 ( .B1(keyFF_keystate_gff_4_SFF_0_n9), 
        .B2(keyFF_outputPar[8]), .C1(keyFF_keystate_gff_4_SFF_0_n10), .C2(
        keyFF_outputPar[15]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_4_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_4_SFF_0_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_4_SFF_0_n10) );
  INV_X1 keyFF_keystate_gff_4_SFF_0_U2 ( .A(keyFF_keystate_gff_4_SFF_0_n10), 
        .ZN(keyFF_keystate_gff_4_SFF_0_n9) );
  DFF_X1 keyFF_keystate_gff_4_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_4_SFF_0_n6), .CK(clk), .Q(keyFF_outputPar[12]), 
        .QN(keyFF_keystate_gff_4_SFF_0_n7) );
  OAI21_X1 keyFF_keystate_gff_4_SFF_1_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_4_SFF_1_n7), .A(keyFF_keystate_gff_4_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_4_SFF_1_n6) );
  OAI221_X1 keyFF_keystate_gff_4_SFF_1_U4 ( .B1(keyFF_keystate_gff_4_SFF_1_n9), 
        .B2(keyFF_outputPar[9]), .C1(keyFF_keystate_gff_4_SFF_1_n10), .C2(
        keyFF_outputPar[16]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_4_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_4_SFF_1_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_4_SFF_1_n10) );
  INV_X1 keyFF_keystate_gff_4_SFF_1_U2 ( .A(keyFF_keystate_gff_4_SFF_1_n10), 
        .ZN(keyFF_keystate_gff_4_SFF_1_n9) );
  DFF_X1 keyFF_keystate_gff_4_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_4_SFF_1_n6), .CK(clk), .Q(keyFF_outputPar[13]), 
        .QN(keyFF_keystate_gff_4_SFF_1_n7) );
  OAI21_X1 keyFF_keystate_gff_4_SFF_2_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_4_SFF_2_n7), .A(keyFF_keystate_gff_4_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_4_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_4_SFF_2_U4 ( .B1(keyFF_keystate_gff_4_SFF_2_n9), 
        .B2(keyFF_outputPar[10]), .C1(keyFF_keystate_gff_4_SFF_2_n10), .C2(
        keyFF_outputPar[17]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_4_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_4_SFF_2_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_4_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_4_SFF_2_U2 ( .A(keyFF_keystate_gff_4_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_4_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_4_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_4_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[14]), 
        .QN(keyFF_keystate_gff_4_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_4_SFF_3_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_4_SFF_3_n7), .A(keyFF_keystate_gff_4_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_4_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_4_SFF_3_U4 ( .B1(keyFF_keystate_gff_4_SFF_3_n9), 
        .B2(keyFF_outputPar[11]), .C1(keyFF_keystate_gff_4_SFF_3_n10), .C2(
        keyFF_counterAdd[0]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_4_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_4_SFF_3_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_4_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_4_SFF_3_U2 ( .A(keyFF_keystate_gff_4_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_4_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_4_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_4_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[15]), 
        .QN(keyFF_keystate_gff_4_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_5_SFF_0_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_5_SFF_0_n8), .A(keyFF_keystate_gff_5_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_5_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_5_SFF_0_U4 ( .B1(keyFF_keystate_gff_5_SFF_0_n10), .B2(keyFF_outputPar[12]), .C1(keyFF_keystate_gff_5_SFF_0_n11), .C2(
        keyFF_counterAdd[1]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_5_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_5_SFF_0_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_5_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_5_SFF_0_U2 ( .A(keyFF_keystate_gff_5_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_5_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_5_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_5_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[16]), 
        .QN(keyFF_keystate_gff_5_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_5_SFF_1_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_5_SFF_1_n8), .A(keyFF_keystate_gff_5_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_5_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_5_SFF_1_U4 ( .B1(keyFF_keystate_gff_5_SFF_1_n10), .B2(keyFF_outputPar[13]), .C1(keyFF_keystate_gff_5_SFF_1_n11), .C2(
        keyFF_counterAdd[2]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_5_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_5_SFF_1_U3 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_5_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_5_SFF_1_U2 ( .A(keyFF_keystate_gff_5_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_5_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_5_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_5_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[17]), 
        .QN(keyFF_keystate_gff_5_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_5_SFF_2_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_5_SFF_2_n8), .A(keyFF_keystate_gff_5_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_5_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_5_SFF_2_U3 ( .B1(keyFF_keystate_n14), .B2(
        keyFF_outputPar[14]), .C1(keyFF_keystate_gff_5_SFF_2_n10), .C2(
        keyFF_counterAdd[3]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_5_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_5_SFF_2_U2 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_5_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_5_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_5_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[18]), 
        .QN(keyFF_keystate_gff_5_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_5_SFF_3_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_5_SFF_3_n8), .A(keyFF_keystate_gff_5_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_5_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_5_SFF_3_U3 ( .B1(keyFF_keystate_n14), .B2(
        keyFF_outputPar[15]), .C1(keyFF_keystate_gff_5_SFF_3_n10), .C2(
        keyFF_counterAdd[4]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_5_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_5_SFF_3_U2 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_5_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_5_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_5_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[19]), 
        .QN(keyFF_keystate_gff_5_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_6_SFF_0_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_6_SFF_0_n8), .A(keyFF_keystate_gff_6_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_6_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_6_SFF_0_U3 ( .B1(keyFF_keystate_n14), .B2(
        keyFF_outputPar[16]), .C1(keyFF_keystate_gff_6_SFF_0_n10), .C2(
        keyFF_outputPar[23]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_6_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_6_SFF_0_U2 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_6_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_6_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_6_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[20]), 
        .QN(keyFF_keystate_gff_6_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_6_SFF_1_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_6_SFF_1_n8), .A(keyFF_keystate_gff_6_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_6_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_6_SFF_1_U3 ( .B1(keyFF_keystate_n14), .B2(
        keyFF_outputPar[17]), .C1(keyFF_keystate_gff_6_SFF_1_n10), .C2(
        keyFF_outputPar[24]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_6_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_6_SFF_1_U2 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_6_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_6_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_6_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[21]), 
        .QN(keyFF_keystate_gff_6_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_6_SFF_2_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_6_SFF_2_n8), .A(keyFF_keystate_gff_6_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_6_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_6_SFF_2_U3 ( .B1(keyFF_keystate_n14), .B2(
        keyFF_outputPar[18]), .C1(keyFF_keystate_gff_6_SFF_2_n10), .C2(
        keyFF_outputPar[25]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_6_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_6_SFF_2_U2 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_6_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_6_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_6_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[22]), 
        .QN(keyFF_keystate_gff_6_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_6_SFF_3_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_6_SFF_3_n8), .A(keyFF_keystate_gff_6_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_6_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_6_SFF_3_U3 ( .B1(keyFF_keystate_n14), .B2(
        keyFF_outputPar[19]), .C1(keyFF_keystate_gff_6_SFF_3_n10), .C2(
        keyFF_outputPar[26]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_6_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_6_SFF_3_U2 ( .A(keyFF_keystate_n14), .ZN(
        keyFF_keystate_gff_6_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_6_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_6_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[23]), 
        .QN(keyFF_keystate_gff_6_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_7_SFF_0_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_7_SFF_0_n8), .A(keyFF_keystate_gff_7_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_7_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_7_SFF_0_U4 ( .B1(keyFF_keystate_gff_7_SFF_0_n10), .B2(keyFF_outputPar[20]), .C1(keyFF_keystate_gff_7_SFF_0_n11), .C2(
        keyFF_outputPar[27]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_7_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_7_SFF_0_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_7_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_7_SFF_0_U2 ( .A(keyFF_keystate_gff_7_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_7_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_7_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_7_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[24]), 
        .QN(keyFF_keystate_gff_7_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_7_SFF_1_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_7_SFF_1_n8), .A(keyFF_keystate_gff_7_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_7_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_7_SFF_1_U4 ( .B1(keyFF_keystate_gff_7_SFF_1_n10), .B2(keyFF_outputPar[21]), .C1(keyFF_keystate_gff_7_SFF_1_n11), .C2(
        keyFF_outputPar[28]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_7_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_7_SFF_1_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_7_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_7_SFF_1_U2 ( .A(keyFF_keystate_gff_7_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_7_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_7_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_7_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[25]), 
        .QN(keyFF_keystate_gff_7_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_7_SFF_2_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_7_SFF_2_n7), .A(keyFF_keystate_gff_7_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_7_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_7_SFF_2_U4 ( .B1(keyFF_keystate_gff_7_SFF_2_n9), 
        .B2(keyFF_outputPar[22]), .C1(keyFF_keystate_gff_7_SFF_2_n10), .C2(
        keyFF_outputPar[29]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_7_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_7_SFF_2_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_7_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_7_SFF_2_U2 ( .A(keyFF_keystate_gff_7_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_7_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_7_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_7_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[26]), 
        .QN(keyFF_keystate_gff_7_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_7_SFF_3_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_7_SFF_3_n7), .A(keyFF_keystate_gff_7_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_7_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_7_SFF_3_U4 ( .B1(keyFF_keystate_gff_7_SFF_3_n9), 
        .B2(keyFF_outputPar[23]), .C1(keyFF_keystate_gff_7_SFF_3_n10), .C2(
        keyFF_outputPar[30]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_7_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_7_SFF_3_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_7_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_7_SFF_3_U2 ( .A(keyFF_keystate_gff_7_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_7_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_7_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_7_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[27]), 
        .QN(keyFF_keystate_gff_7_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_8_SFF_0_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_8_SFF_0_n7), .A(keyFF_keystate_gff_8_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_8_SFF_0_n6) );
  OAI221_X1 keyFF_keystate_gff_8_SFF_0_U4 ( .B1(keyFF_keystate_gff_8_SFF_0_n9), 
        .B2(keyFF_outputPar[24]), .C1(keyFF_keystate_gff_8_SFF_0_n10), .C2(
        keyFF_outputPar[31]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_8_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_8_SFF_0_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_8_SFF_0_n10) );
  INV_X1 keyFF_keystate_gff_8_SFF_0_U2 ( .A(keyFF_keystate_gff_8_SFF_0_n10), 
        .ZN(keyFF_keystate_gff_8_SFF_0_n9) );
  DFF_X1 keyFF_keystate_gff_8_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_8_SFF_0_n6), .CK(clk), .Q(keyFF_outputPar[28]), 
        .QN(keyFF_keystate_gff_8_SFF_0_n7) );
  OAI21_X1 keyFF_keystate_gff_8_SFF_1_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_8_SFF_1_n7), .A(keyFF_keystate_gff_8_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_8_SFF_1_n6) );
  OAI221_X1 keyFF_keystate_gff_8_SFF_1_U4 ( .B1(keyFF_keystate_gff_8_SFF_1_n9), 
        .B2(keyFF_outputPar[25]), .C1(keyFF_keystate_gff_8_SFF_1_n10), .C2(
        keyFF_outputPar[32]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_8_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_8_SFF_1_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_8_SFF_1_n10) );
  INV_X1 keyFF_keystate_gff_8_SFF_1_U2 ( .A(keyFF_keystate_gff_8_SFF_1_n10), 
        .ZN(keyFF_keystate_gff_8_SFF_1_n9) );
  DFF_X1 keyFF_keystate_gff_8_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_8_SFF_1_n6), .CK(clk), .Q(keyFF_outputPar[29]), 
        .QN(keyFF_keystate_gff_8_SFF_1_n7) );
  OAI21_X1 keyFF_keystate_gff_8_SFF_2_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_8_SFF_2_n7), .A(keyFF_keystate_gff_8_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_8_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_8_SFF_2_U4 ( .B1(keyFF_keystate_gff_8_SFF_2_n9), 
        .B2(keyFF_outputPar[26]), .C1(keyFF_keystate_gff_8_SFF_2_n10), .C2(
        keyFF_outputPar[33]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_8_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_8_SFF_2_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_8_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_8_SFF_2_U2 ( .A(keyFF_keystate_gff_8_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_8_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_8_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_8_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[30]), 
        .QN(keyFF_keystate_gff_8_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_8_SFF_3_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_8_SFF_3_n7), .A(keyFF_keystate_gff_8_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_8_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_8_SFF_3_U4 ( .B1(keyFF_keystate_gff_8_SFF_3_n9), 
        .B2(keyFF_outputPar[27]), .C1(keyFF_keystate_gff_8_SFF_3_n10), .C2(
        keyFF_outputPar[34]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_8_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_8_SFF_3_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_8_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_8_SFF_3_U2 ( .A(keyFF_keystate_gff_8_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_8_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_8_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_8_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[31]), 
        .QN(keyFF_keystate_gff_8_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_9_SFF_0_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_9_SFF_0_n8), .A(keyFF_keystate_gff_9_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_9_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_9_SFF_0_U4 ( .B1(keyFF_keystate_gff_9_SFF_0_n10), .B2(keyFF_outputPar[28]), .C1(keyFF_keystate_gff_9_SFF_0_n11), .C2(
        keyFF_outputPar[35]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_9_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_9_SFF_0_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_9_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_9_SFF_0_U2 ( .A(keyFF_keystate_gff_9_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_9_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_9_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_9_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[32]), 
        .QN(keyFF_keystate_gff_9_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_9_SFF_1_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_9_SFF_1_n8), .A(keyFF_keystate_gff_9_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_9_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_9_SFF_1_U4 ( .B1(keyFF_keystate_gff_9_SFF_1_n10), .B2(keyFF_outputPar[29]), .C1(keyFF_keystate_gff_9_SFF_1_n11), .C2(
        keyFF_outputPar[36]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_9_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_9_SFF_1_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_9_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_9_SFF_1_U2 ( .A(keyFF_keystate_gff_9_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_9_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_9_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_9_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[33]), 
        .QN(keyFF_keystate_gff_9_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_9_SFF_2_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_9_SFF_2_n8), .A(keyFF_keystate_gff_9_SFF_2_n12), 
        .ZN(keyFF_keystate_gff_9_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_9_SFF_2_U4 ( .B1(keyFF_keystate_gff_9_SFF_2_n10), .B2(keyFF_outputPar[30]), .C1(keyFF_keystate_gff_9_SFF_2_n11), .C2(
        keyFF_outputPar[37]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_9_SFF_2_n12) );
  INV_X1 keyFF_keystate_gff_9_SFF_2_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_9_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_9_SFF_2_U2 ( .A(keyFF_keystate_gff_9_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_9_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_9_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_9_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[34]), 
        .QN(keyFF_keystate_gff_9_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_9_SFF_3_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_9_SFF_3_n8), .A(keyFF_keystate_gff_9_SFF_3_n12), 
        .ZN(keyFF_keystate_gff_9_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_9_SFF_3_U4 ( .B1(keyFF_keystate_gff_9_SFF_3_n10), .B2(keyFF_outputPar[31]), .C1(keyFF_keystate_gff_9_SFF_3_n11), .C2(
        keyFF_outputPar[38]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_9_SFF_3_n12) );
  INV_X1 keyFF_keystate_gff_9_SFF_3_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_9_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_9_SFF_3_U2 ( .A(keyFF_keystate_gff_9_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_9_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_9_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_9_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[35]), 
        .QN(keyFF_keystate_gff_9_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_10_SFF_0_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_10_SFF_0_n8), .A(keyFF_keystate_gff_10_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_10_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_10_SFF_0_U4 ( .B1(
        keyFF_keystate_gff_10_SFF_0_n10), .B2(keyFF_outputPar[32]), .C1(
        keyFF_keystate_gff_10_SFF_0_n11), .C2(keyFF_outputPar[39]), .A(
        keyFF_keystate_n10), .ZN(keyFF_keystate_gff_10_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_10_SFF_0_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_10_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_10_SFF_0_U2 ( .A(keyFF_keystate_gff_10_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_10_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_10_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_10_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[36]), 
        .QN(keyFF_keystate_gff_10_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_10_SFF_1_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_10_SFF_1_n8), .A(keyFF_keystate_gff_10_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_10_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_10_SFF_1_U4 ( .B1(
        keyFF_keystate_gff_10_SFF_1_n10), .B2(keyFF_outputPar[33]), .C1(
        keyFF_keystate_gff_10_SFF_1_n11), .C2(keyFF_outputPar[40]), .A(
        keyFF_keystate_n10), .ZN(keyFF_keystate_gff_10_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_10_SFF_1_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_10_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_10_SFF_1_U2 ( .A(keyFF_keystate_gff_10_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_10_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_10_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_10_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[37]), 
        .QN(keyFF_keystate_gff_10_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_10_SFF_2_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_10_SFF_2_n8), .A(keyFF_keystate_gff_10_SFF_2_n12), 
        .ZN(keyFF_keystate_gff_10_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_10_SFF_2_U4 ( .B1(
        keyFF_keystate_gff_10_SFF_2_n10), .B2(keyFF_outputPar[34]), .C1(
        keyFF_keystate_gff_10_SFF_2_n11), .C2(keyFF_outputPar[41]), .A(
        keyFF_keystate_n10), .ZN(keyFF_keystate_gff_10_SFF_2_n12) );
  INV_X1 keyFF_keystate_gff_10_SFF_2_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_10_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_10_SFF_2_U2 ( .A(keyFF_keystate_gff_10_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_10_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_10_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_10_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[38]), 
        .QN(keyFF_keystate_gff_10_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_10_SFF_3_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_10_SFF_3_n8), .A(keyFF_keystate_gff_10_SFF_3_n12), 
        .ZN(keyFF_keystate_gff_10_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_10_SFF_3_U4 ( .B1(
        keyFF_keystate_gff_10_SFF_3_n10), .B2(keyFF_outputPar[35]), .C1(
        keyFF_keystate_gff_10_SFF_3_n11), .C2(keyFF_outputPar[42]), .A(
        keyFF_keystate_n10), .ZN(keyFF_keystate_gff_10_SFF_3_n12) );
  INV_X1 keyFF_keystate_gff_10_SFF_3_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_10_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_10_SFF_3_U2 ( .A(keyFF_keystate_gff_10_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_10_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_10_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_10_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[39]), 
        .QN(keyFF_keystate_gff_10_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_11_SFF_0_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_11_SFF_0_n8), .A(keyFF_keystate_gff_11_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_11_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_11_SFF_0_U3 ( .B1(keyFF_keystate_n17), .B2(
        keyFF_outputPar[36]), .C1(keyFF_keystate_gff_11_SFF_0_n10), .C2(
        keyFF_outputPar[43]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_11_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_11_SFF_0_U2 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_11_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_11_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_11_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[40]), 
        .QN(keyFF_keystate_gff_11_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_11_SFF_1_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_11_SFF_1_n8), .A(keyFF_keystate_gff_11_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_11_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_11_SFF_1_U3 ( .B1(keyFF_keystate_n17), .B2(
        keyFF_outputPar[37]), .C1(keyFF_keystate_gff_11_SFF_1_n10), .C2(
        keyFF_outputPar[44]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_11_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_11_SFF_1_U2 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_11_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_11_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_11_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[41]), 
        .QN(keyFF_keystate_gff_11_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_11_SFF_2_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_11_SFF_2_n7), .A(keyFF_keystate_gff_11_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_11_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_11_SFF_2_U4 ( .B1(
        keyFF_keystate_gff_11_SFF_2_n9), .B2(keyFF_outputPar[38]), .C1(
        keyFF_keystate_gff_11_SFF_2_n10), .C2(keyFF_outputPar[45]), .A(
        keyFF_keystate_n12), .ZN(keyFF_keystate_gff_11_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_11_SFF_2_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_11_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_11_SFF_2_U2 ( .A(keyFF_keystate_gff_11_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_11_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_11_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_11_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[42]), 
        .QN(keyFF_keystate_gff_11_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_11_SFF_3_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_11_SFF_3_n7), .A(keyFF_keystate_gff_11_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_11_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_11_SFF_3_U4 ( .B1(
        keyFF_keystate_gff_11_SFF_3_n9), .B2(keyFF_outputPar[39]), .C1(
        keyFF_keystate_gff_11_SFF_3_n10), .C2(keyFF_outputPar[46]), .A(
        keyFF_keystate_n12), .ZN(keyFF_keystate_gff_11_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_11_SFF_3_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_11_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_11_SFF_3_U2 ( .A(keyFF_keystate_gff_11_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_11_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_11_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_11_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[43]), 
        .QN(keyFF_keystate_gff_11_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_12_SFF_0_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_12_SFF_0_n7), .A(keyFF_keystate_gff_12_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_12_SFF_0_n6) );
  OAI221_X1 keyFF_keystate_gff_12_SFF_0_U4 ( .B1(
        keyFF_keystate_gff_12_SFF_0_n9), .B2(keyFF_outputPar[40]), .C1(
        keyFF_keystate_gff_12_SFF_0_n10), .C2(keyFF_outputPar[47]), .A(
        keyFF_keystate_n13), .ZN(keyFF_keystate_gff_12_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_12_SFF_0_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_12_SFF_0_n10) );
  INV_X1 keyFF_keystate_gff_12_SFF_0_U2 ( .A(keyFF_keystate_gff_12_SFF_0_n10), 
        .ZN(keyFF_keystate_gff_12_SFF_0_n9) );
  DFF_X1 keyFF_keystate_gff_12_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_12_SFF_0_n6), .CK(clk), .Q(keyFF_outputPar[44]), 
        .QN(keyFF_keystate_gff_12_SFF_0_n7) );
  OAI21_X1 keyFF_keystate_gff_12_SFF_1_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_12_SFF_1_n7), .A(keyFF_keystate_gff_12_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_12_SFF_1_n6) );
  OAI221_X1 keyFF_keystate_gff_12_SFF_1_U4 ( .B1(
        keyFF_keystate_gff_12_SFF_1_n9), .B2(keyFF_outputPar[41]), .C1(
        keyFF_keystate_gff_12_SFF_1_n10), .C2(keyFF_outputPar[48]), .A(
        keyFF_keystate_n13), .ZN(keyFF_keystate_gff_12_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_12_SFF_1_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_12_SFF_1_n10) );
  INV_X1 keyFF_keystate_gff_12_SFF_1_U2 ( .A(keyFF_keystate_gff_12_SFF_1_n10), 
        .ZN(keyFF_keystate_gff_12_SFF_1_n9) );
  DFF_X1 keyFF_keystate_gff_12_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_12_SFF_1_n6), .CK(clk), .Q(keyFF_outputPar[45]), 
        .QN(keyFF_keystate_gff_12_SFF_1_n7) );
  OAI21_X1 keyFF_keystate_gff_12_SFF_2_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_12_SFF_2_n7), .A(keyFF_keystate_gff_12_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_12_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_12_SFF_2_U4 ( .B1(
        keyFF_keystate_gff_12_SFF_2_n9), .B2(keyFF_outputPar[42]), .C1(
        keyFF_keystate_gff_12_SFF_2_n10), .C2(keyFF_outputPar[49]), .A(
        keyFF_keystate_n13), .ZN(keyFF_keystate_gff_12_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_12_SFF_2_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_12_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_12_SFF_2_U2 ( .A(keyFF_keystate_gff_12_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_12_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_12_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_12_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[46]), 
        .QN(keyFF_keystate_gff_12_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_12_SFF_3_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_12_SFF_3_n7), .A(keyFF_keystate_gff_12_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_12_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_12_SFF_3_U4 ( .B1(
        keyFF_keystate_gff_12_SFF_3_n9), .B2(keyFF_outputPar[43]), .C1(
        keyFF_keystate_gff_12_SFF_3_n10), .C2(keyFF_outputPar[50]), .A(
        keyFF_keystate_n13), .ZN(keyFF_keystate_gff_12_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_12_SFF_3_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_12_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_12_SFF_3_U2 ( .A(keyFF_keystate_gff_12_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_12_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_12_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_12_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[47]), 
        .QN(keyFF_keystate_gff_12_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_13_SFF_0_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_13_SFF_0_n8), .A(keyFF_keystate_gff_13_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_13_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_13_SFF_0_U4 ( .B1(
        keyFF_keystate_gff_13_SFF_0_n10), .B2(keyFF_outputPar[44]), .C1(
        keyFF_keystate_gff_13_SFF_0_n11), .C2(keyFF_outputPar[51]), .A(
        keyFF_keystate_n10), .ZN(keyFF_keystate_gff_13_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_13_SFF_0_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_13_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_13_SFF_0_U2 ( .A(keyFF_keystate_gff_13_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_13_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_13_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_13_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[48]), 
        .QN(keyFF_keystate_gff_13_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_13_SFF_1_U5 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_13_SFF_1_n8), .A(keyFF_keystate_gff_13_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_13_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_13_SFF_1_U4 ( .B1(
        keyFF_keystate_gff_13_SFF_1_n10), .B2(keyFF_outputPar[45]), .C1(
        keyFF_keystate_gff_13_SFF_1_n11), .C2(keyFF_outputPar[52]), .A(
        keyFF_keystate_n10), .ZN(keyFF_keystate_gff_13_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_13_SFF_1_U3 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_13_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_13_SFF_1_U2 ( .A(keyFF_keystate_gff_13_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_13_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_13_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_13_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[49]), 
        .QN(keyFF_keystate_gff_13_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_13_SFF_2_U4 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_13_SFF_2_n8), .A(keyFF_keystate_gff_13_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_13_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_13_SFF_2_U3 ( .B1(keyFF_keystate_n15), .B2(
        keyFF_outputPar[46]), .C1(keyFF_keystate_gff_13_SFF_2_n10), .C2(
        keyFF_outputPar[53]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_13_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_13_SFF_2_U2 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_13_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_13_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_13_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[50]), 
        .QN(keyFF_keystate_gff_13_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_13_SFF_3_U4 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_13_SFF_3_n8), .A(keyFF_keystate_gff_13_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_13_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_13_SFF_3_U3 ( .B1(keyFF_keystate_n15), .B2(
        keyFF_outputPar[47]), .C1(keyFF_keystate_gff_13_SFF_3_n10), .C2(
        keyFF_outputPar[54]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_13_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_13_SFF_3_U2 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_13_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_13_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_13_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[51]), 
        .QN(keyFF_keystate_gff_13_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_14_SFF_0_U4 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_14_SFF_0_n8), .A(keyFF_keystate_gff_14_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_14_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_14_SFF_0_U3 ( .B1(keyFF_keystate_n15), .B2(
        keyFF_outputPar[48]), .C1(keyFF_keystate_gff_14_SFF_0_n10), .C2(
        keyFF_outputPar[55]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_14_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_14_SFF_0_U2 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_14_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_14_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_14_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[52]), 
        .QN(keyFF_keystate_gff_14_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_14_SFF_1_U4 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_14_SFF_1_n8), .A(keyFF_keystate_gff_14_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_14_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_14_SFF_1_U3 ( .B1(keyFF_keystate_n15), .B2(
        keyFF_outputPar[49]), .C1(keyFF_keystate_gff_14_SFF_1_n10), .C2(
        keyFF_outputPar[56]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_14_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_14_SFF_1_U2 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_14_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_14_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_14_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[53]), 
        .QN(keyFF_keystate_gff_14_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_14_SFF_2_U4 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_14_SFF_2_n8), .A(keyFF_keystate_gff_14_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_14_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_14_SFF_2_U3 ( .B1(keyFF_keystate_n15), .B2(
        keyFF_outputPar[50]), .C1(keyFF_keystate_gff_14_SFF_2_n10), .C2(
        keyFF_outputPar[57]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_14_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_14_SFF_2_U2 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_14_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_14_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_14_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[54]), 
        .QN(keyFF_keystate_gff_14_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_14_SFF_3_U4 ( .B1(keyFF_keystate_n10), .B2(
        keyFF_keystate_gff_14_SFF_3_n8), .A(keyFF_keystate_gff_14_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_14_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_14_SFF_3_U3 ( .B1(keyFF_keystate_n15), .B2(
        keyFF_outputPar[51]), .C1(keyFF_keystate_gff_14_SFF_3_n10), .C2(
        keyFF_outputPar[58]), .A(keyFF_keystate_n10), .ZN(
        keyFF_keystate_gff_14_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_14_SFF_3_U2 ( .A(keyFF_keystate_n15), .ZN(
        keyFF_keystate_gff_14_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_14_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_14_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[55]), 
        .QN(keyFF_keystate_gff_14_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_15_SFF_0_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_15_SFF_0_n8), .A(keyFF_keystate_gff_15_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_15_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_15_SFF_0_U3 ( .B1(keyFF_keystate_n17), .B2(
        keyFF_outputPar[52]), .C1(keyFF_keystate_gff_15_SFF_0_n10), .C2(
        keyFF_outputPar[59]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_15_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_15_SFF_0_U2 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_15_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_15_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_15_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[56]), 
        .QN(keyFF_keystate_gff_15_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_15_SFF_1_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_15_SFF_1_n8), .A(keyFF_keystate_gff_15_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_15_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_15_SFF_1_U3 ( .B1(keyFF_keystate_n17), .B2(
        keyFF_outputPar[53]), .C1(keyFF_keystate_gff_15_SFF_1_n10), .C2(
        keyFF_outputPar[60]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_15_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_15_SFF_1_U2 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_15_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_15_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_15_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[57]), 
        .QN(keyFF_keystate_gff_15_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_15_SFF_2_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_15_SFF_2_n7), .A(keyFF_keystate_gff_15_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_15_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_15_SFF_2_U4 ( .B1(
        keyFF_keystate_gff_15_SFF_2_n9), .B2(keyFF_outputPar[54]), .C1(
        keyFF_keystate_gff_15_SFF_2_n10), .C2(keyFF_outputPar[61]), .A(
        keyFF_keystate_n12), .ZN(keyFF_keystate_gff_15_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_15_SFF_2_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_15_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_15_SFF_2_U2 ( .A(keyFF_keystate_gff_15_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_15_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_15_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_15_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[58]), 
        .QN(keyFF_keystate_gff_15_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_15_SFF_3_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_15_SFF_3_n7), .A(keyFF_keystate_gff_15_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_15_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_15_SFF_3_U4 ( .B1(
        keyFF_keystate_gff_15_SFF_3_n9), .B2(keyFF_outputPar[55]), .C1(
        keyFF_keystate_gff_15_SFF_3_n10), .C2(keyFF_outputPar[62]), .A(
        keyFF_keystate_n12), .ZN(keyFF_keystate_gff_15_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_15_SFF_3_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_15_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_15_SFF_3_U2 ( .A(keyFF_keystate_gff_15_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_15_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_15_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_15_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[59]), 
        .QN(keyFF_keystate_gff_15_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_16_SFF_0_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_16_SFF_0_n7), .A(keyFF_keystate_gff_16_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_16_SFF_0_n6) );
  OAI221_X1 keyFF_keystate_gff_16_SFF_0_U4 ( .B1(
        keyFF_keystate_gff_16_SFF_0_n9), .B2(keyFF_outputPar[56]), .C1(
        keyFF_keystate_gff_16_SFF_0_n10), .C2(keyFF_outputPar[63]), .A(
        keyFF_keystate_n13), .ZN(keyFF_keystate_gff_16_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_16_SFF_0_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_16_SFF_0_n10) );
  INV_X1 keyFF_keystate_gff_16_SFF_0_U2 ( .A(keyFF_keystate_gff_16_SFF_0_n10), 
        .ZN(keyFF_keystate_gff_16_SFF_0_n9) );
  DFF_X1 keyFF_keystate_gff_16_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_16_SFF_0_n6), .CK(clk), .Q(keyFF_outputPar[60]), 
        .QN(keyFF_keystate_gff_16_SFF_0_n7) );
  OAI21_X1 keyFF_keystate_gff_16_SFF_1_U5 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_16_SFF_1_n7), .A(keyFF_keystate_gff_16_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_16_SFF_1_n6) );
  OAI221_X1 keyFF_keystate_gff_16_SFF_1_U4 ( .B1(
        keyFF_keystate_gff_16_SFF_1_n9), .B2(keyFF_outputPar[57]), .C1(
        keyFF_keystate_gff_16_SFF_1_n10), .C2(keyFF_outputPar[64]), .A(
        keyFF_keystate_n13), .ZN(keyFF_keystate_gff_16_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_16_SFF_1_U3 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_16_SFF_1_n10) );
  INV_X1 keyFF_keystate_gff_16_SFF_1_U2 ( .A(keyFF_keystate_gff_16_SFF_1_n10), 
        .ZN(keyFF_keystate_gff_16_SFF_1_n9) );
  DFF_X1 keyFF_keystate_gff_16_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_16_SFF_1_n6), .CK(clk), .Q(keyFF_outputPar[61]), 
        .QN(keyFF_keystate_gff_16_SFF_1_n7) );
  OAI21_X1 keyFF_keystate_gff_16_SFF_2_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_16_SFF_2_n7), .A(keyFF_keystate_gff_16_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_16_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_16_SFF_2_U3 ( .B1(keyFF_keystate_n18), .B2(
        keyFF_outputPar[58]), .C1(keyFF_keystate_gff_16_SFF_2_n9), .C2(
        keyFF_outputPar[65]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_16_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_16_SFF_2_U2 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_16_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_16_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_16_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[62]), 
        .QN(keyFF_keystate_gff_16_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_16_SFF_3_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_16_SFF_3_n7), .A(keyFF_keystate_gff_16_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_16_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_16_SFF_3_U3 ( .B1(keyFF_keystate_n18), .B2(
        keyFF_outputPar[59]), .C1(keyFF_keystate_gff_16_SFF_3_n9), .C2(
        keyFF_outputPar[66]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_16_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_16_SFF_3_U2 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_16_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_16_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_16_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[63]), 
        .QN(keyFF_keystate_gff_16_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_17_SFF_0_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_17_SFF_0_n8), .A(keyFF_keystate_gff_17_SFF_0_n12), 
        .ZN(keyFF_keystate_gff_17_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_17_SFF_0_U4 ( .B1(
        keyFF_keystate_gff_17_SFF_0_n10), .B2(keyFF_outputPar[60]), .C1(
        keyFF_keystate_gff_17_SFF_0_n11), .C2(keyFF_outputPar[67]), .A(
        keyFF_keystate_n11), .ZN(keyFF_keystate_gff_17_SFF_0_n12) );
  INV_X1 keyFF_keystate_gff_17_SFF_0_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_17_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_17_SFF_0_U2 ( .A(keyFF_keystate_gff_17_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_17_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_17_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_17_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[64]), 
        .QN(keyFF_keystate_gff_17_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_17_SFF_1_U5 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_17_SFF_1_n8), .A(keyFF_keystate_gff_17_SFF_1_n12), 
        .ZN(keyFF_keystate_gff_17_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_17_SFF_1_U4 ( .B1(
        keyFF_keystate_gff_17_SFF_1_n10), .B2(keyFF_outputPar[61]), .C1(
        keyFF_keystate_gff_17_SFF_1_n11), .C2(keyFF_outputPar[68]), .A(
        keyFF_keystate_n11), .ZN(keyFF_keystate_gff_17_SFF_1_n12) );
  INV_X1 keyFF_keystate_gff_17_SFF_1_U3 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_17_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_17_SFF_1_U2 ( .A(keyFF_keystate_gff_17_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_17_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_17_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_17_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[65]), 
        .QN(keyFF_keystate_gff_17_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_17_SFF_2_U4 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_17_SFF_2_n8), .A(keyFF_keystate_gff_17_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_17_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_17_SFF_2_U3 ( .B1(keyFF_keystate_n16), .B2(
        keyFF_outputPar[62]), .C1(keyFF_keystate_gff_17_SFF_2_n10), .C2(
        keyFF_outputPar[69]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_17_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_17_SFF_2_U2 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_17_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_17_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_17_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[66]), 
        .QN(keyFF_keystate_gff_17_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_17_SFF_3_U4 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_17_SFF_3_n8), .A(keyFF_keystate_gff_17_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_17_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_17_SFF_3_U3 ( .B1(keyFF_keystate_n16), .B2(
        keyFF_outputPar[63]), .C1(keyFF_keystate_gff_17_SFF_3_n10), .C2(
        keyFF_outputPar[70]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_17_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_17_SFF_3_U2 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_17_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_17_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_17_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[67]), 
        .QN(keyFF_keystate_gff_17_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_18_SFF_0_U4 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_18_SFF_0_n8), .A(keyFF_keystate_gff_18_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_18_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_18_SFF_0_U3 ( .B1(keyFF_keystate_n16), .B2(
        keyFF_outputPar[64]), .C1(keyFF_keystate_gff_18_SFF_0_n10), .C2(
        keyFF_outputPar[71]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_18_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_18_SFF_0_U2 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_18_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_18_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_18_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[68]), 
        .QN(keyFF_keystate_gff_18_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_18_SFF_1_U4 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_18_SFF_1_n8), .A(keyFF_keystate_gff_18_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_18_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_18_SFF_1_U3 ( .B1(keyFF_keystate_n16), .B2(
        keyFF_outputPar[65]), .C1(keyFF_keystate_gff_18_SFF_1_n10), .C2(
        keyFF_outputPar[72]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_18_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_18_SFF_1_U2 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_18_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_18_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_18_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[69]), 
        .QN(keyFF_keystate_gff_18_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_18_SFF_2_U4 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_18_SFF_2_n8), .A(keyFF_keystate_gff_18_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_18_SFF_2_n7) );
  OAI221_X1 keyFF_keystate_gff_18_SFF_2_U3 ( .B1(keyFF_keystate_n16), .B2(
        keyFF_outputPar[66]), .C1(keyFF_keystate_gff_18_SFF_2_n10), .C2(
        keyFF_outputPar[73]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_18_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_18_SFF_2_U2 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_18_SFF_2_n10) );
  DFF_X1 keyFF_keystate_gff_18_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_18_SFF_2_n7), .CK(clk), .Q(keyFF_outputPar[70]), 
        .QN(keyFF_keystate_gff_18_SFF_2_n8) );
  OAI21_X1 keyFF_keystate_gff_18_SFF_3_U4 ( .B1(keyFF_keystate_n11), .B2(
        keyFF_keystate_gff_18_SFF_3_n8), .A(keyFF_keystate_gff_18_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_18_SFF_3_n7) );
  OAI221_X1 keyFF_keystate_gff_18_SFF_3_U3 ( .B1(keyFF_keystate_n16), .B2(
        keyFF_outputPar[67]), .C1(keyFF_keystate_gff_18_SFF_3_n10), .C2(
        keyFF_outputPar[74]), .A(keyFF_keystate_n11), .ZN(
        keyFF_keystate_gff_18_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_18_SFF_3_U2 ( .A(keyFF_keystate_n16), .ZN(
        keyFF_keystate_gff_18_SFF_3_n10) );
  DFF_X1 keyFF_keystate_gff_18_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_18_SFF_3_n7), .CK(clk), .Q(keyFF_outputPar[71]), 
        .QN(keyFF_keystate_gff_18_SFF_3_n8) );
  OAI21_X1 keyFF_keystate_gff_19_SFF_0_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_19_SFF_0_n8), .A(keyFF_keystate_gff_19_SFF_0_n11), 
        .ZN(keyFF_keystate_gff_19_SFF_0_n7) );
  OAI221_X1 keyFF_keystate_gff_19_SFF_0_U3 ( .B1(keyFF_keystate_n17), .B2(
        keyFF_outputPar[68]), .C1(keyFF_keystate_gff_19_SFF_0_n10), .C2(
        keyFF_outputPar[75]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_19_SFF_0_n11) );
  INV_X1 keyFF_keystate_gff_19_SFF_0_U2 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_19_SFF_0_n10) );
  DFF_X1 keyFF_keystate_gff_19_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_19_SFF_0_n7), .CK(clk), .Q(keyFF_outputPar[72]), 
        .QN(keyFF_keystate_gff_19_SFF_0_n8) );
  OAI21_X1 keyFF_keystate_gff_19_SFF_1_U4 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_19_SFF_1_n8), .A(keyFF_keystate_gff_19_SFF_1_n11), 
        .ZN(keyFF_keystate_gff_19_SFF_1_n7) );
  OAI221_X1 keyFF_keystate_gff_19_SFF_1_U3 ( .B1(keyFF_keystate_n17), .B2(
        keyFF_outputPar[69]), .C1(keyFF_keystate_gff_19_SFF_1_n10), .C2(
        roundkey[0]), .A(keyFF_keystate_n12), .ZN(
        keyFF_keystate_gff_19_SFF_1_n11) );
  INV_X1 keyFF_keystate_gff_19_SFF_1_U2 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_19_SFF_1_n10) );
  DFF_X1 keyFF_keystate_gff_19_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_19_SFF_1_n7), .CK(clk), .Q(keyFF_outputPar[73]), 
        .QN(keyFF_keystate_gff_19_SFF_1_n8) );
  OAI21_X1 keyFF_keystate_gff_19_SFF_2_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_19_SFF_2_n7), .A(keyFF_keystate_gff_19_SFF_2_n11), 
        .ZN(keyFF_keystate_gff_19_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_19_SFF_2_U4 ( .B1(
        keyFF_keystate_gff_19_SFF_2_n9), .B2(keyFF_outputPar[70]), .C1(
        keyFF_keystate_gff_19_SFF_2_n10), .C2(roundkey[1]), .A(
        keyFF_keystate_n12), .ZN(keyFF_keystate_gff_19_SFF_2_n11) );
  INV_X1 keyFF_keystate_gff_19_SFF_2_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_19_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_19_SFF_2_U2 ( .A(keyFF_keystate_gff_19_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_19_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_19_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_19_SFF_2_n6), .CK(clk), .Q(keyFF_outputPar[74]), 
        .QN(keyFF_keystate_gff_19_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_19_SFF_3_U5 ( .B1(keyFF_keystate_n12), .B2(
        keyFF_keystate_gff_19_SFF_3_n7), .A(keyFF_keystate_gff_19_SFF_3_n11), 
        .ZN(keyFF_keystate_gff_19_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_19_SFF_3_U4 ( .B1(
        keyFF_keystate_gff_19_SFF_3_n9), .B2(keyFF_outputPar[71]), .C1(
        keyFF_keystate_gff_19_SFF_3_n10), .C2(roundkey[2]), .A(
        keyFF_keystate_n12), .ZN(keyFF_keystate_gff_19_SFF_3_n11) );
  INV_X1 keyFF_keystate_gff_19_SFF_3_U3 ( .A(keyFF_keystate_n17), .ZN(
        keyFF_keystate_gff_19_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_19_SFF_3_U2 ( .A(keyFF_keystate_gff_19_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_19_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_19_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_19_SFF_3_n6), .CK(clk), .Q(keyFF_outputPar[75]), 
        .QN(keyFF_keystate_gff_19_SFF_3_n7) );
  OAI21_X1 keyFF_keystate_gff_20_SFF_0_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_20_SFF_0_n7), .A(keyFF_keystate_gff_20_SFF_0_n10), 
        .ZN(keyFF_keystate_gff_20_SFF_0_n6) );
  OAI221_X1 keyFF_keystate_gff_20_SFF_0_U3 ( .B1(keyFF_keystate_n18), .B2(
        keyFF_outputPar[72]), .C1(keyFF_keystate_gff_20_SFF_0_n9), .C2(
        sboxKS[0]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_20_SFF_0_n10) );
  INV_X1 keyFF_keystate_gff_20_SFF_0_U2 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_20_SFF_0_n9) );
  DFF_X1 keyFF_keystate_gff_20_SFF_0_Cell_reg ( .D(
        keyFF_keystate_gff_20_SFF_0_n6), .CK(clk), .Q(roundkey[0]), .QN(
        keyFF_keystate_gff_20_SFF_0_n7) );
  OAI21_X1 keyFF_keystate_gff_20_SFF_1_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_20_SFF_1_n7), .A(keyFF_keystate_gff_20_SFF_1_n10), 
        .ZN(keyFF_keystate_gff_20_SFF_1_n6) );
  OAI221_X1 keyFF_keystate_gff_20_SFF_1_U3 ( .B1(keyFF_keystate_n18), .B2(
        keyFF_outputPar[73]), .C1(keyFF_keystate_gff_20_SFF_1_n9), .C2(
        sboxKS[1]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_20_SFF_1_n10) );
  INV_X1 keyFF_keystate_gff_20_SFF_1_U2 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_20_SFF_1_n9) );
  DFF_X1 keyFF_keystate_gff_20_SFF_1_Cell_reg ( .D(
        keyFF_keystate_gff_20_SFF_1_n6), .CK(clk), .Q(roundkey[1]), .QN(
        keyFF_keystate_gff_20_SFF_1_n7) );
  OAI21_X1 keyFF_keystate_gff_20_SFF_2_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_20_SFF_2_n7), .A(keyFF_keystate_gff_20_SFF_2_n10), 
        .ZN(keyFF_keystate_gff_20_SFF_2_n6) );
  OAI221_X1 keyFF_keystate_gff_20_SFF_2_U3 ( .B1(keyFF_keystate_n18), .B2(
        keyFF_outputPar[74]), .C1(keyFF_keystate_gff_20_SFF_2_n9), .C2(
        sboxKS[2]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_20_SFF_2_n10) );
  INV_X1 keyFF_keystate_gff_20_SFF_2_U2 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_20_SFF_2_n9) );
  DFF_X1 keyFF_keystate_gff_20_SFF_2_Cell_reg ( .D(
        keyFF_keystate_gff_20_SFF_2_n6), .CK(clk), .Q(roundkey[2]), .QN(
        keyFF_keystate_gff_20_SFF_2_n7) );
  OAI21_X1 keyFF_keystate_gff_20_SFF_3_U4 ( .B1(keyFF_keystate_n13), .B2(
        keyFF_keystate_gff_20_SFF_3_n7), .A(keyFF_keystate_gff_20_SFF_3_n10), 
        .ZN(keyFF_keystate_gff_20_SFF_3_n6) );
  OAI221_X1 keyFF_keystate_gff_20_SFF_3_U3 ( .B1(keyFF_keystate_n18), .B2(
        keyFF_outputPar[75]), .C1(keyFF_keystate_gff_20_SFF_3_n9), .C2(
        sboxKS[3]), .A(keyFF_keystate_n13), .ZN(
        keyFF_keystate_gff_20_SFF_3_n10) );
  INV_X1 keyFF_keystate_gff_20_SFF_3_U2 ( .A(keyFF_keystate_n18), .ZN(
        keyFF_keystate_gff_20_SFF_3_n9) );
  DFF_X1 keyFF_keystate_gff_20_SFF_3_Cell_reg ( .D(
        keyFF_keystate_gff_20_SFF_3_n6), .CK(clk), .Q(roundkey[3]), .QN(
        keyFF_keystate_gff_20_SFF_3_n7) );
  INV_X1 sbox_Inst_N_F1_U10 ( .A(sbox_Inst_N_F1_n10), .ZN(sbox_g[1]) );
  AOI211_X1 sbox_Inst_N_F1_U9 ( .C1(dataOut1[1]), .C2(dataOut1[2]), .A(
        sbox_Inst_N_F1_n9), .B(dataOut1[3]), .ZN(sbox_Inst_N_F1_n10) );
  INV_X1 sbox_Inst_N_F1_U8 ( .A(sbox_f[1]), .ZN(sbox_h[1]) );
  AOI221_X1 sbox_Inst_N_F1_U7 ( .B1(sbox_Inst_N_F1_n8), .B2(dataOut1[2]), .C1(
        dataOut1[3]), .C2(dataOut1[1]), .A(sbox_Inst_N_F1_n9), .ZN(sbox_f[1])
         );
  OAI21_X1 sbox_Inst_N_F1_U6 ( .B1(dataOut1[1]), .B2(dataOut1[2]), .A(
        dataOut2[0]), .ZN(sbox_Inst_N_F1_n9) );
  XNOR2_X1 sbox_Inst_N_F1_U5 ( .A(sbox_Inst_N_F1_n7), .B(sbox_Inst_N_F1_n6), 
        .ZN(sbox_e[1]) );
  NAND2_X1 sbox_Inst_N_F1_U4 ( .A1(dataOut1[2]), .A2(sbox_Inst_N_F1_n5), .ZN(
        sbox_Inst_N_F1_n6) );
  INV_X1 sbox_Inst_N_F1_U3 ( .A(dataOut1[1]), .ZN(sbox_Inst_N_F1_n5) );
  XNOR2_X1 sbox_Inst_N_F1_U2 ( .A(dataOut2[0]), .B(sbox_Inst_N_F1_n8), .ZN(
        sbox_Inst_N_F1_n7) );
  INV_X1 sbox_Inst_N_F1_U1 ( .A(dataOut1[3]), .ZN(sbox_Inst_N_F1_n8) );
  AOI211_X1 sbox_Inst_N_F2_U8 ( .C1(sbox_Inst_N_F2_n9), .C2(dataOut1[1]), .A(
        dataOut2[3]), .B(sbox_Inst_N_F2_n8), .ZN(sbox_g[2]) );
  OAI21_X1 sbox_Inst_N_F2_U7 ( .B1(sbox_Inst_N_F2_n9), .B2(dataOut1[1]), .A(
        dataOut1[0]), .ZN(sbox_Inst_N_F2_n8) );
  NOR2_X1 sbox_Inst_N_F2_U6 ( .A1(sbox_Inst_N_F2_n7), .A2(sbox_Inst_N_F2_n6), 
        .ZN(sbox_f[2]) );
  INV_X1 sbox_Inst_N_F2_U5 ( .A(dataOut1[0]), .ZN(sbox_Inst_N_F2_n6) );
  NOR2_X1 sbox_Inst_N_F2_U4 ( .A1(dataOut1[0]), .A2(sbox_Inst_N_F2_n7), .ZN(
        sbox_h[2]) );
  OAI221_X1 sbox_Inst_N_F2_U3 ( .B1(dataOut2[3]), .B2(dataOut1[2]), .C1(
        dataOut1[1]), .C2(sbox_Inst_N_F2_n9), .A(sbox_Inst_N_F2_n5), .ZN(
        sbox_Inst_N_F2_n7) );
  NAND2_X1 sbox_Inst_N_F2_U2 ( .A1(dataOut2[3]), .A2(dataOut1[1]), .ZN(
        sbox_Inst_N_F2_n5) );
  INV_X1 sbox_Inst_N_F2_U1 ( .A(dataOut1[2]), .ZN(sbox_Inst_N_F2_n9) );
  AOI211_X1 sbox_Inst_N_F3_U10 ( .C1(sbox_Inst_N_F3_n10), .C2(
        sbox_Inst_N_F3_n9), .A(sbox_Inst_N_F3_n8), .B(sbox_Inst_N_F3_n7), .ZN(
        sbox_g[3]) );
  AOI21_X1 sbox_Inst_N_F3_U9 ( .B1(sbox_Inst_N_F3_n6), .B2(sbox_Inst_N_F3_n5), 
        .A(sbox_Inst_N_F3_n7), .ZN(sbox_f[3]) );
  OAI21_X1 sbox_Inst_N_F3_U8 ( .B1(sbox_Inst_N_F3_n10), .B2(sbox_Inst_N_F3_n9), 
        .A(sbox_Inst_N_F3_n4), .ZN(sbox_Inst_N_F3_n7) );
  INV_X1 sbox_Inst_N_F3_U7 ( .A(dataOut1[1]), .ZN(sbox_Inst_N_F3_n9) );
  AOI221_X1 sbox_Inst_N_F3_U6 ( .B1(dataOut1[1]), .B2(sbox_Inst_N_F3_n6), .C1(
        sbox_Inst_N_F3_n5), .C2(sbox_Inst_N_F3_n6), .A(sbox_Inst_N_F3_n4), 
        .ZN(sbox_h[3]) );
  INV_X1 sbox_Inst_N_F3_U5 ( .A(dataOut1[0]), .ZN(sbox_Inst_N_F3_n4) );
  NAND2_X1 sbox_Inst_N_F3_U4 ( .A1(dataOut2[2]), .A2(sbox_Inst_N_F3_n8), .ZN(
        sbox_Inst_N_F3_n5) );
  INV_X1 sbox_Inst_N_F3_U3 ( .A(dataOut1[3]), .ZN(sbox_Inst_N_F3_n8) );
  NAND3_X1 sbox_Inst_N_F3_U2 ( .A1(dataOut1[1]), .A2(dataOut1[3]), .A3(
        sbox_Inst_N_F3_n10), .ZN(sbox_Inst_N_F3_n6) );
  INV_X1 sbox_Inst_N_F3_U1 ( .A(dataOut2[2]), .ZN(sbox_Inst_N_F3_n10) );
  NAND2_X1 sbox_Inst_N_F4_U14 ( .A1(sbox_Inst_N_F4_n13), .A2(
        sbox_Inst_N_F4_n12), .ZN(sbox_g[4]) );
  OAI221_X1 sbox_Inst_N_F4_U13 ( .B1(dataOut2[3]), .B2(sbox_Inst_N_F4_n11), 
        .C1(sbox_Inst_N_F4_n10), .C2(dataOut2[2]), .A(dataOut2[0]), .ZN(
        sbox_Inst_N_F4_n12) );
  OAI221_X1 sbox_Inst_N_F4_U12 ( .B1(dataOut2[3]), .B2(dataOut2[2]), .C1(
        sbox_Inst_N_F4_n10), .C2(dataOut1[1]), .A(sbox_Inst_N_F4_n9), .ZN(
        sbox_Inst_N_F4_n13) );
  OAI221_X1 sbox_Inst_N_F4_U11 ( .B1(dataOut2[0]), .B2(sbox_Inst_N_F4_n8), 
        .C1(sbox_Inst_N_F4_n9), .C2(sbox_Inst_N_F4_n10), .A(sbox_Inst_N_F4_n7), 
        .ZN(sbox_f[4]) );
  OAI22_X1 sbox_Inst_N_F4_U10 ( .A1(sbox_Inst_N_F4_n9), .A2(sbox_Inst_N_F4_n6), 
        .B1(dataOut1[1]), .B2(sbox_Inst_N_F4_n5), .ZN(sbox_e[2]) );
  INV_X1 sbox_Inst_N_F4_U9 ( .A(sbox_Inst_N_F4_n4), .ZN(sbox_Inst_N_F4_n5) );
  NOR2_X1 sbox_Inst_N_F4_U8 ( .A1(sbox_Inst_N_F4_n11), .A2(dataOut1[1]), .ZN(
        sbox_Inst_N_F4_n6) );
  OAI211_X1 sbox_Inst_N_F4_U7 ( .C1(dataOut2[3]), .C2(sbox_Inst_N_F4_n9), .A(
        sbox_Inst_N_F4_n8), .B(sbox_Inst_N_F4_n7), .ZN(sbox_h[4]) );
  NAND2_X1 sbox_Inst_N_F4_U6 ( .A1(dataOut1[1]), .A2(sbox_Inst_N_F4_n4), .ZN(
        sbox_Inst_N_F4_n7) );
  NOR2_X1 sbox_Inst_N_F4_U5 ( .A1(dataOut2[0]), .A2(sbox_Inst_N_F4_n11), .ZN(
        sbox_Inst_N_F4_n4) );
  INV_X1 sbox_Inst_N_F4_U4 ( .A(dataOut2[2]), .ZN(sbox_Inst_N_F4_n11) );
  OAI21_X1 sbox_Inst_N_F4_U3 ( .B1(dataOut2[2]), .B2(dataOut1[1]), .A(
        sbox_Inst_N_F4_n10), .ZN(sbox_Inst_N_F4_n8) );
  INV_X1 sbox_Inst_N_F4_U2 ( .A(dataOut2[3]), .ZN(sbox_Inst_N_F4_n10) );
  INV_X1 sbox_Inst_N_F4_U1 ( .A(dataOut2[0]), .ZN(sbox_Inst_N_F4_n9) );
  NOR4_X1 sbox_Inst_N_F5_U11 ( .A1(dataOut1[3]), .A2(sbox_Inst_N_F5_n11), .A3(
        sbox_Inst_N_F5_n10), .A4(sbox_Inst_N_F5_n9), .ZN(sbox_g[5]) );
  INV_X1 sbox_Inst_N_F5_U10 ( .A(sbox_Inst_N_F5_n8), .ZN(sbox_Inst_N_F5_n10)
         );
  AOI22_X1 sbox_Inst_N_F5_U9 ( .A1(dataOut1[3]), .A2(dataOut1[0]), .B1(
        sbox_Inst_N_F5_n7), .B2(sbox_Inst_N_F5_n6), .ZN(sbox_f[5]) );
  AOI21_X1 sbox_Inst_N_F5_U8 ( .B1(dataOut1[3]), .B2(sbox_Inst_N_F5_n8), .A(
        dataOut1[0]), .ZN(sbox_Inst_N_F5_n6) );
  OAI21_X1 sbox_Inst_N_F5_U7 ( .B1(sbox_Inst_N_F5_n9), .B2(sbox_Inst_N_F5_n7), 
        .A(sbox_Inst_N_F5_n5), .ZN(sbox_h[5]) );
  OAI21_X1 sbox_Inst_N_F5_U6 ( .B1(sbox_Inst_N_F5_n9), .B2(sbox_Inst_N_F5_n8), 
        .A(dataOut1[3]), .ZN(sbox_Inst_N_F5_n5) );
  NAND2_X1 sbox_Inst_N_F5_U5 ( .A1(dataOut1[2]), .A2(sbox_Inst_N_F5_n4), .ZN(
        sbox_Inst_N_F5_n8) );
  INV_X1 sbox_Inst_N_F5_U4 ( .A(sbox_Inst_N_F5_n11), .ZN(sbox_Inst_N_F5_n7) );
  NOR2_X1 sbox_Inst_N_F5_U3 ( .A1(sbox_Inst_N_F5_n4), .A2(dataOut1[2]), .ZN(
        sbox_Inst_N_F5_n11) );
  INV_X1 sbox_Inst_N_F5_U2 ( .A(dataOut2[1]), .ZN(sbox_Inst_N_F5_n4) );
  INV_X1 sbox_Inst_N_F5_U1 ( .A(dataOut1[0]), .ZN(sbox_Inst_N_F5_n9) );
  NAND3_X1 sbox_Inst_N_F6_U10 ( .A1(sbox_Inst_N_F6_n9), .A2(sbox_Inst_N_F6_n8), 
        .A3(sbox_Inst_N_F6_n7), .ZN(sbox_g[6]) );
  OAI221_X1 sbox_Inst_N_F6_U9 ( .B1(dataOut2[3]), .B2(sbox_Inst_N_F6_n6), .C1(
        sbox_Inst_N_F6_n5), .C2(dataOut1[2]), .A(dataOut2[0]), .ZN(
        sbox_Inst_N_F6_n7) );
  AOI22_X1 sbox_Inst_N_F6_U8 ( .A1(dataOut2[1]), .A2(sbox_Inst_N_F6_n9), .B1(
        sbox_Inst_N_F6_n8), .B2(sbox_Inst_N_F6_n6), .ZN(sbox_f[6]) );
  INV_X1 sbox_Inst_N_F6_U7 ( .A(dataOut2[1]), .ZN(sbox_Inst_N_F6_n6) );
  OR3_X1 sbox_Inst_N_F6_U6 ( .A1(sbox_Inst_N_F6_n5), .A2(dataOut1[2]), .A3(
        dataOut2[0]), .ZN(sbox_Inst_N_F6_n8) );
  NAND3_X1 sbox_Inst_N_F6_U5 ( .A1(dataOut1[2]), .A2(sbox_Inst_N_F6_n5), .A3(
        sbox_Inst_N_F6_n4), .ZN(sbox_Inst_N_F6_n9) );
  INV_X1 sbox_Inst_N_F6_U4 ( .A(dataOut2[3]), .ZN(sbox_Inst_N_F6_n5) );
  XOR2_X1 sbox_Inst_N_F6_U3 ( .A(sbox_Inst_N_F6_n3), .B(sbox_Inst_N_F6_n4), 
        .Z(sbox_e[3]) );
  INV_X1 sbox_Inst_N_F6_U2 ( .A(dataOut2[0]), .ZN(sbox_Inst_N_F6_n4) );
  NAND2_X1 sbox_Inst_N_F6_U1 ( .A1(dataOut1[2]), .A2(dataOut2[1]), .ZN(
        sbox_Inst_N_F6_n3) );
  NOR3_X1 sbox_Inst_N_F7_U7 ( .A1(dataOut2[0]), .A2(sbox_Inst_N_F7_n6), .A3(
        sbox_Inst_N_F7_n5), .ZN(sbox_g[7]) );
  INV_X1 sbox_Inst_N_F7_U6 ( .A(sbox_Inst_N_F7_n4), .ZN(sbox_f[7]) );
  OAI211_X1 sbox_Inst_N_F7_U5 ( .C1(dataOut1[3]), .C2(sbox_Inst_N_F7_n6), .A(
        dataOut2[0]), .B(sbox_Inst_N_F7_n5), .ZN(sbox_Inst_N_F7_n4) );
  NAND2_X1 sbox_Inst_N_F7_U4 ( .A1(dataOut1[3]), .A2(sbox_Inst_N_F7_n3), .ZN(
        sbox_Inst_N_F7_n5) );
  NAND2_X1 sbox_Inst_N_F7_U3 ( .A1(dataOut2[1]), .A2(sbox_Inst_N_F7_n2), .ZN(
        sbox_Inst_N_F7_n3) );
  NOR2_X1 sbox_Inst_N_F7_U2 ( .A1(dataOut2[1]), .A2(sbox_Inst_N_F7_n2), .ZN(
        sbox_Inst_N_F7_n6) );
  INV_X1 sbox_Inst_N_F7_U1 ( .A(dataOut2[2]), .ZN(sbox_Inst_N_F7_n2) );
  AND3_X1 sbox_Inst_N_F8_U10 ( .A1(sbox_Inst_N_F8_n8), .A2(dataOut2[3]), .A3(
        sbox_Inst_N_F8_n7), .ZN(sbox_g[8]) );
  NOR3_X1 sbox_Inst_N_F8_U9 ( .A1(sbox_Inst_N_F8_n8), .A2(sbox_Inst_N_F8_n6), 
        .A3(sbox_Inst_N_F8_n7), .ZN(sbox_f[8]) );
  INV_X1 sbox_Inst_N_F8_U8 ( .A(dataOut1[0]), .ZN(sbox_Inst_N_F8_n7) );
  INV_X1 sbox_Inst_N_F8_U7 ( .A(sbox_Inst_N_F8_n5), .ZN(sbox_Inst_N_F8_n8) );
  AOI21_X1 sbox_Inst_N_F8_U6 ( .B1(sbox_Inst_N_F8_n6), .B2(dataOut1[0]), .A(
        sbox_Inst_N_F8_n4), .ZN(sbox_e[4]) );
  NAND2_X1 sbox_Inst_N_F8_U5 ( .A1(sbox_Inst_N_F8_n4), .A2(sbox_Inst_N_F8_n5), 
        .ZN(sbox_h[8]) );
  OAI21_X1 sbox_Inst_N_F8_U4 ( .B1(dataOut2[2]), .B2(dataOut2[1]), .A(
        sbox_Inst_N_F8_n3), .ZN(sbox_Inst_N_F8_n5) );
  NOR2_X1 sbox_Inst_N_F8_U3 ( .A1(dataOut1[0]), .A2(sbox_Inst_N_F8_n6), .ZN(
        sbox_Inst_N_F8_n4) );
  XNOR2_X1 sbox_Inst_N_F8_U2 ( .A(dataOut2[3]), .B(sbox_Inst_N_F8_n3), .ZN(
        sbox_Inst_N_F8_n6) );
  NAND2_X1 sbox_Inst_N_F8_U1 ( .A1(dataOut2[2]), .A2(dataOut2[1]), .ZN(
        sbox_Inst_N_F8_n3) );
  DFF_X1 sbox_Gen_reg_Q_reg_4_ ( .D(sbox_f[5]), .CK(clk), .Q(sbox_f_reg[5]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_24_ ( .D(sbox_h[5]), .CK(clk), .Q(sbox_h_reg[5]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_17_ ( .D(sbox_g[6]), .CK(clk), .Q(sbox_g_reg[6]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_15_ ( .D(sbox_g[4]), .CK(clk), .Q(sbox_g_reg[4]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_1_ ( .D(sbox_f[2]), .CK(clk), .Q(sbox_f_reg[2]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_22_ ( .D(sbox_h[3]), .CK(clk), .Q(sbox_h_reg[3]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_6_ ( .D(sbox_f[7]), .CK(clk), .Q(sbox_f_reg[7]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_26_ ( .D(sbox_f[7]), .CK(clk), .Q(sbox_h_reg[7]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_2_ ( .D(sbox_f[3]), .CK(clk), .Q(sbox_f_reg[3]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_0_ ( .D(sbox_f[1]), .CK(clk), .Q(sbox_f_reg[1]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_13_ ( .D(sbox_g[2]), .CK(clk), .Q(sbox_g_reg[2]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_20_ ( .D(sbox_h[1]), .CK(clk), .Q(sbox_h_reg[1]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_21_ ( .D(sbox_h[2]), .CK(clk), .Q(sbox_h_reg[2]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_8_ ( .D(sbox_e[1]), .CK(clk), .Q(sbox_e_reg[1]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_11_ ( .D(sbox_e[4]), .CK(clk), .Q(sbox_e_reg[4]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_5_ ( .D(sbox_f[6]), .CK(clk), .Q(sbox_f_reg[6]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_25_ ( .D(sbox_f[6]), .CK(clk), .Q(sbox_h_reg[6]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_12_ ( .D(sbox_g[1]), .CK(clk), .Q(sbox_g_reg[1]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_10_ ( .D(sbox_e[3]), .CK(clk), .Q(sbox_e_reg[3]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_3_ ( .D(sbox_f[4]), .CK(clk), .Q(sbox_f_reg[4]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_23_ ( .D(sbox_h[4]), .CK(clk), .Q(sbox_h_reg[4]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_14_ ( .D(sbox_g[3]), .CK(clk), .Q(sbox_g_reg[3]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_18_ ( .D(sbox_g[7]), .CK(clk), .Q(sbox_g_reg[7]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_9_ ( .D(sbox_e[2]), .CK(clk), .Q(sbox_e_reg[2]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_7_ ( .D(sbox_f[8]), .CK(clk), .Q(sbox_f_reg[8]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_16_ ( .D(sbox_g[5]), .CK(clk), .Q(sbox_g_reg[5]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_27_ ( .D(sbox_h[8]), .CK(clk), .Q(sbox_h_reg[8]), 
        .QN() );
  DFF_X1 sbox_Gen_reg_Q_reg_19_ ( .D(sbox_g[8]), .CK(clk), .Q(sbox_g_reg[8]), 
        .QN() );
  XNOR2_X1 sbox_Inst_L_XORInst1_U3 ( .A(sbox_Inst_L_XORInst1_n6), .B(
        sbox_Inst_L_XORInst1_n5), .ZN(share1[1]) );
  XNOR2_X1 sbox_Inst_L_XORInst1_U2 ( .A(sbox_f_reg[3]), .B(sbox_f_reg[4]), 
        .ZN(sbox_Inst_L_XORInst1_n5) );
  XOR2_X1 sbox_Inst_L_XORInst1_U1 ( .A(sbox_f_reg[1]), .B(sbox_f_reg[2]), .Z(
        sbox_Inst_L_XORInst1_n6) );
  XNOR2_X1 sbox_Inst_L_XORInst2_U3 ( .A(sbox_Inst_L_XORInst2_n6), .B(
        sbox_Inst_L_XORInst2_n5), .ZN(share2[1]) );
  XNOR2_X1 sbox_Inst_L_XORInst2_U2 ( .A(sbox_f_reg[7]), .B(sbox_f_reg[8]), 
        .ZN(sbox_Inst_L_XORInst2_n5) );
  XOR2_X1 sbox_Inst_L_XORInst2_U1 ( .A(sbox_f_reg[5]), .B(sbox_f_reg[6]), .Z(
        sbox_Inst_L_XORInst2_n6) );
  XOR2_X1 sbox_Inst_L_XORInst3_U1 ( .A(sbox_e_reg[1]), .B(sbox_e_reg[2]), .Z(
        share1[0]) );
  XOR2_X1 sbox_Inst_L_XORInst4_U1 ( .A(sbox_e_reg[3]), .B(sbox_e_reg[4]), .Z(
        share2[0]) );
  XNOR2_X1 sbox_Inst_L_XORInst5_U3 ( .A(sbox_Inst_L_XORInst5_n6), .B(
        sbox_Inst_L_XORInst5_n5), .ZN(share1[2]) );
  XNOR2_X1 sbox_Inst_L_XORInst5_U2 ( .A(sbox_g_reg[3]), .B(sbox_g_reg[4]), 
        .ZN(sbox_Inst_L_XORInst5_n5) );
  XOR2_X1 sbox_Inst_L_XORInst5_U1 ( .A(sbox_g_reg[1]), .B(sbox_g_reg[2]), .Z(
        sbox_Inst_L_XORInst5_n6) );
  XNOR2_X1 sbox_Inst_L_XORInst6_U3 ( .A(sbox_Inst_L_XORInst6_n6), .B(
        sbox_Inst_L_XORInst6_n5), .ZN(share2[2]) );
  XNOR2_X1 sbox_Inst_L_XORInst6_U2 ( .A(sbox_g_reg[7]), .B(sbox_g_reg[8]), 
        .ZN(sbox_Inst_L_XORInst6_n5) );
  XOR2_X1 sbox_Inst_L_XORInst6_U1 ( .A(sbox_g_reg[5]), .B(sbox_g_reg[6]), .Z(
        sbox_Inst_L_XORInst6_n6) );
  XNOR2_X1 sbox_Inst_L_XORInst7_U3 ( .A(sbox_Inst_L_XORInst7_n6), .B(
        sbox_Inst_L_XORInst7_n5), .ZN(share1[3]) );
  XNOR2_X1 sbox_Inst_L_XORInst7_U2 ( .A(sbox_h_reg[3]), .B(sbox_h_reg[4]), 
        .ZN(sbox_Inst_L_XORInst7_n5) );
  XOR2_X1 sbox_Inst_L_XORInst7_U1 ( .A(sbox_h_reg[1]), .B(sbox_h_reg[2]), .Z(
        sbox_Inst_L_XORInst7_n6) );
  XNOR2_X1 sbox_Inst_L_XORInst8_U3 ( .A(sbox_Inst_L_XORInst8_n6), .B(
        sbox_Inst_L_XORInst8_n5), .ZN(share2[3]) );
  XNOR2_X1 sbox_Inst_L_XORInst8_U2 ( .A(sbox_h_reg[7]), .B(sbox_h_reg[8]), 
        .ZN(sbox_Inst_L_XORInst8_n5) );
  XOR2_X1 sbox_Inst_L_XORInst8_U1 ( .A(sbox_h_reg[5]), .B(sbox_h_reg[6]), .Z(
        sbox_Inst_L_XORInst8_n6) );
  OAI22_X1 sbox_KS_U18 ( .A1(keyRegKS[3]), .A2(sbox_KS_n18), .B1(keyRegKS[2]), 
        .B2(sbox_KS_n17), .ZN(sboxKS[3]) );
  AOI21_X1 sbox_KS_U17 ( .B1(sbox_KS_n18), .B2(keyRegKS[3]), .A(sbox_KS_n16), 
        .ZN(sbox_KS_n17) );
  INV_X1 sbox_KS_U16 ( .A(sbox_KS_n15), .ZN(sbox_KS_n16) );
  OAI21_X1 sbox_KS_U15 ( .B1(sbox_KS_n14), .B2(sbox_KS_n13), .A(sbox_KS_n12), 
        .ZN(sboxKS[2]) );
  OAI211_X1 sbox_KS_U14 ( .C1(sbox_KS_n18), .C2(sbox_KS_n11), .A(sbox_KS_n10), 
        .B(sbox_KS_n15), .ZN(sbox_KS_n12) );
  INV_X1 sbox_KS_U13 ( .A(sbox_KS_n9), .ZN(sbox_KS_n18) );
  OAI21_X1 sbox_KS_U12 ( .B1(roundkey[3]), .B2(keyRegKS[1]), .A(sbox_KS_n15), 
        .ZN(sbox_KS_n9) );
  AOI22_X1 sbox_KS_U11 ( .A1(sbox_KS_n8), .A2(sbox_KS_n7), .B1(sbox_KS_n13), 
        .B2(sbox_KS_n14), .ZN(sboxKS[1]) );
  AOI22_X1 sbox_KS_U10 ( .A1(keyRegKS[3]), .A2(sbox_KS_n15), .B1(keyRegKS[1]), 
        .B2(sbox_KS_n11), .ZN(sbox_KS_n13) );
  INV_X1 sbox_KS_U9 ( .A(keyRegKS[3]), .ZN(sbox_KS_n11) );
  OAI21_X1 sbox_KS_U8 ( .B1(keyRegKS[2]), .B2(roundkey[3]), .A(keyRegKS[1]), 
        .ZN(sbox_KS_n15) );
  INV_X1 sbox_KS_U7 ( .A(sbox_KS_n14), .ZN(sbox_KS_n8) );
  OAI21_X1 sbox_KS_U6 ( .B1(roundkey[3]), .B2(keyRegKS[3]), .A(keyRegKS[2]), 
        .ZN(sbox_KS_n14) );
  XNOR2_X1 sbox_KS_U5 ( .A(sbox_KS_n6), .B(sbox_KS_n5), .ZN(sboxKS[0]) );
  OAI21_X1 sbox_KS_U4 ( .B1(roundkey[3]), .B2(keyRegKS[3]), .A(sbox_KS_n7), 
        .ZN(sbox_KS_n5) );
  NAND2_X1 sbox_KS_U3 ( .A1(roundkey[3]), .A2(keyRegKS[3]), .ZN(sbox_KS_n7) );
  NOR2_X1 sbox_KS_U2 ( .A1(sbox_KS_n10), .A2(keyRegKS[1]), .ZN(sbox_KS_n6) );
  INV_X1 sbox_KS_U1 ( .A(keyRegKS[2]), .ZN(sbox_KS_n10) );
endmodule

