module circuit ( clk, reset, r, input1, input2, input3, output1, output2, 
        output3, Key1, Key2, Key3, enc_dec, done );
  input [127:0] r;
  input [63:0] input1;
  input [63:0] input2;
  input [63:0] input3;
  output [63:0] output1;
  output [63:0] output2;
  output [63:0] output3;
  input [127:0] Key1;
  input [127:0] Key2;
  input [127:0] Key3;
  input clk, reset, enc_dec;
  output done;
  wire   EN, controller_roundCounter_n34, controller_roundCounter_n33,
         controller_roundCounter_n32, controller_roundCounter_n31,
         controller_roundCounter_n30, controller_roundCounter_n29,
         controller_roundCounter_n28, controller_roundCounter_n27,
         controller_roundCounter_n26, controller_roundCounter_n25,
         controller_roundCounter_n24, controller_roundCounter_n23,
         controller_roundCounter_n22, controller_roundCounter_n15,
         controller_roundCounter_n14, controller_roundCounter_n13,
         controller_roundCounter_n12, controller_roundCounter_n11,
         controller_roundCounter_n10, controller_roundCounter_q_0_,
         controller_roundCounter_q_1_, Midori_rounds_n2068,
         Midori_rounds_n2067, Midori_rounds_n2066, Midori_rounds_n2065,
         Midori_rounds_n2064, Midori_rounds_n2063, Midori_rounds_n2062,
         Midori_rounds_n2061, Midori_rounds_n2060, Midori_rounds_n2059,
         Midori_rounds_n2058, Midori_rounds_n2057, Midori_rounds_n2056,
         Midori_rounds_n2055, Midori_rounds_n2054, Midori_rounds_n2053,
         Midori_rounds_n2052, Midori_rounds_n2051, Midori_rounds_n2050,
         Midori_rounds_n2049, Midori_rounds_n2048, Midori_rounds_n2047,
         Midori_rounds_n2046, Midori_rounds_n2045, Midori_rounds_n2044,
         Midori_rounds_n2043, Midori_rounds_n2042, Midori_rounds_n2041,
         Midori_rounds_n2040, Midori_rounds_n2039, Midori_rounds_n2038,
         Midori_rounds_n2037, Midori_rounds_n2036, Midori_rounds_n2035,
         Midori_rounds_n2034, Midori_rounds_n2033, Midori_rounds_n2032,
         Midori_rounds_n2031, Midori_rounds_n2030, Midori_rounds_n2029,
         Midori_rounds_n2028, Midori_rounds_n2027, Midori_rounds_n2026,
         Midori_rounds_n2025, Midori_rounds_n2024, Midori_rounds_n2023,
         Midori_rounds_n2022, Midori_rounds_n2021, Midori_rounds_n2020,
         Midori_rounds_n2019, Midori_rounds_n2018, Midori_rounds_n2017,
         Midori_rounds_n2016, Midori_rounds_n2015, Midori_rounds_n2014,
         Midori_rounds_n2013, Midori_rounds_n2012, Midori_rounds_n2011,
         Midori_rounds_n2010, Midori_rounds_n2009, Midori_rounds_n2008,
         Midori_rounds_n2007, Midori_rounds_n2006, Midori_rounds_n2005,
         Midori_rounds_n2004, Midori_rounds_n2003, Midori_rounds_n2002,
         Midori_rounds_n2001, Midori_rounds_n2000, Midori_rounds_n1999,
         Midori_rounds_n1998, Midori_rounds_n1997, Midori_rounds_n1996,
         Midori_rounds_n1995, Midori_rounds_n1994, Midori_rounds_n1993,
         Midori_rounds_n1992, Midori_rounds_n1991, Midori_rounds_n1990,
         Midori_rounds_n1989, Midori_rounds_n1988, Midori_rounds_n1987,
         Midori_rounds_n1986, Midori_rounds_n1985, Midori_rounds_n1984,
         Midori_rounds_n1983, Midori_rounds_n1982, Midori_rounds_n1981,
         Midori_rounds_n1980, Midori_rounds_n1979, Midori_rounds_n1978,
         Midori_rounds_n1977, Midori_rounds_n1976, Midori_rounds_n1975,
         Midori_rounds_n1974, Midori_rounds_n1973, Midori_rounds_n1972,
         Midori_rounds_n1971, Midori_rounds_n1970, Midori_rounds_n1969,
         Midori_rounds_n1968, Midori_rounds_n1967, Midori_rounds_n1966,
         Midori_rounds_n1965, Midori_rounds_n1964, Midori_rounds_n1963,
         Midori_rounds_n1962, Midori_rounds_n1961, Midori_rounds_n1960,
         Midori_rounds_n1959, Midori_rounds_n1958, Midori_rounds_n1957,
         Midori_rounds_n1956, Midori_rounds_n1955, Midori_rounds_n1954,
         Midori_rounds_n1953, Midori_rounds_n1952, Midori_rounds_n1951,
         Midori_rounds_n1950, Midori_rounds_n1949, Midori_rounds_n1948,
         Midori_rounds_n1947, Midori_rounds_n1946, Midori_rounds_n1945,
         Midori_rounds_n1944, Midori_rounds_n1943, Midori_rounds_n1942,
         Midori_rounds_n1941, Midori_rounds_n1940, Midori_rounds_n1939,
         Midori_rounds_n1938, Midori_rounds_n1937, Midori_rounds_n1936,
         Midori_rounds_n1935, Midori_rounds_n1934, Midori_rounds_n1933,
         Midori_rounds_n1932, Midori_rounds_n1931, Midori_rounds_n1930,
         Midori_rounds_n1929, Midori_rounds_n1928, Midori_rounds_n1927,
         Midori_rounds_n1926, Midori_rounds_n1925, Midori_rounds_n1924,
         Midori_rounds_n1923, Midori_rounds_n1922, Midori_rounds_n1921,
         Midori_rounds_n1920, Midori_rounds_n1919, Midori_rounds_n1918,
         Midori_rounds_n1917, Midori_rounds_n1916, Midori_rounds_n1915,
         Midori_rounds_n1914, Midori_rounds_n1913, Midori_rounds_n1912,
         Midori_rounds_n1911, Midori_rounds_n1910, Midori_rounds_n1909,
         Midori_rounds_n1908, Midori_rounds_n1907, Midori_rounds_n1906,
         Midori_rounds_n1905, Midori_rounds_n1904, Midori_rounds_n1903,
         Midori_rounds_n1902, Midori_rounds_n1901, Midori_rounds_n1900,
         Midori_rounds_n1899, Midori_rounds_n1898, Midori_rounds_n1897,
         Midori_rounds_n1896, Midori_rounds_n1895, Midori_rounds_n1894,
         Midori_rounds_n1893, Midori_rounds_n1892, Midori_rounds_n1891,
         Midori_rounds_n1890, Midori_rounds_n1889, Midori_rounds_n1888,
         Midori_rounds_n1887, Midori_rounds_n1886, Midori_rounds_n1885,
         Midori_rounds_n1884, Midori_rounds_n1883, Midori_rounds_n1882,
         Midori_rounds_n1881, Midori_rounds_n1880, Midori_rounds_n1879,
         Midori_rounds_n1878, Midori_rounds_n1877, Midori_rounds_n1876,
         Midori_rounds_n1875, Midori_rounds_n1874, Midori_rounds_n1873,
         Midori_rounds_n1872, Midori_rounds_n1871, Midori_rounds_n1870,
         Midori_rounds_n1869, Midori_rounds_n1868, Midori_rounds_n1867,
         Midori_rounds_n1866, Midori_rounds_n1865, Midori_rounds_n1864,
         Midori_rounds_n1863, Midori_rounds_n1862, Midori_rounds_n1861,
         Midori_rounds_n1860, Midori_rounds_n1859, Midori_rounds_n1858,
         Midori_rounds_n1857, Midori_rounds_n1856, Midori_rounds_n1855,
         Midori_rounds_n1854, Midori_rounds_n1853, Midori_rounds_n1852,
         Midori_rounds_n1851, Midori_rounds_n1850, Midori_rounds_n1849,
         Midori_rounds_n1848, Midori_rounds_n1847, Midori_rounds_n1846,
         Midori_rounds_n1845, Midori_rounds_n1844, Midori_rounds_n1843,
         Midori_rounds_n1842, Midori_rounds_n1841, Midori_rounds_n1840,
         Midori_rounds_n1839, Midori_rounds_n1838, Midori_rounds_n1837,
         Midori_rounds_n1836, Midori_rounds_n1835, Midori_rounds_n1834,
         Midori_rounds_n1833, Midori_rounds_n1832, Midori_rounds_n1831,
         Midori_rounds_n1830, Midori_rounds_n1829, Midori_rounds_n1828,
         Midori_rounds_n1827, Midori_rounds_n1826, Midori_rounds_n1825,
         Midori_rounds_n1824, Midori_rounds_n1823, Midori_rounds_n1822,
         Midori_rounds_n1821, Midori_rounds_n1820, Midori_rounds_n1819,
         Midori_rounds_n1818, Midori_rounds_n1817, Midori_rounds_n1816,
         Midori_rounds_n1815, Midori_rounds_n1814, Midori_rounds_n1813,
         Midori_rounds_n1812, Midori_rounds_n1811, Midori_rounds_n1810,
         Midori_rounds_n1809, Midori_rounds_n1808, Midori_rounds_n1807,
         Midori_rounds_n1806, Midori_rounds_n1805, Midori_rounds_n1804,
         Midori_rounds_n1803, Midori_rounds_n1802, Midori_rounds_n1801,
         Midori_rounds_n1800, Midori_rounds_n1799, Midori_rounds_n1798,
         Midori_rounds_n1797, Midori_rounds_n1796, Midori_rounds_n1795,
         Midori_rounds_n1794, Midori_rounds_n1793, Midori_rounds_n1792,
         Midori_rounds_n1791, Midori_rounds_n1790, Midori_rounds_n1789,
         Midori_rounds_n1788, Midori_rounds_n1787, Midori_rounds_n1786,
         Midori_rounds_n1785, Midori_rounds_n1784, Midori_rounds_n1783,
         Midori_rounds_n1782, Midori_rounds_n1781, Midori_rounds_n1780,
         Midori_rounds_n1779, Midori_rounds_n1778, Midori_rounds_n1777,
         Midori_rounds_n1776, Midori_rounds_n1775, Midori_rounds_n1774,
         Midori_rounds_n1773, Midori_rounds_n1772, Midori_rounds_n1771,
         Midori_rounds_n1770, Midori_rounds_n1769, Midori_rounds_n1768,
         Midori_rounds_n1767, Midori_rounds_n1766, Midori_rounds_n1765,
         Midori_rounds_n1764, Midori_rounds_n1763, Midori_rounds_n1762,
         Midori_rounds_n1761, Midori_rounds_n1760, Midori_rounds_n1759,
         Midori_rounds_n1758, Midori_rounds_n1757, Midori_rounds_n1756,
         Midori_rounds_n1755, Midori_rounds_n1754, Midori_rounds_n1753,
         Midori_rounds_n1752, Midori_rounds_n1751, Midori_rounds_n1750,
         Midori_rounds_n1749, Midori_rounds_n1748, Midori_rounds_n1747,
         Midori_rounds_n1746, Midori_rounds_n1745, Midori_rounds_n1744,
         Midori_rounds_n1743, Midori_rounds_n1742, Midori_rounds_n1741,
         Midori_rounds_n1740, Midori_rounds_n1739, Midori_rounds_n1738,
         Midori_rounds_n1737, Midori_rounds_n1736, Midori_rounds_n1735,
         Midori_rounds_n1734, Midori_rounds_n1733, Midori_rounds_n1732,
         Midori_rounds_n1731, Midori_rounds_n1730, Midori_rounds_n1729,
         Midori_rounds_n1728, Midori_rounds_n1727, Midori_rounds_n1726,
         Midori_rounds_n1725, Midori_rounds_n1724, Midori_rounds_n1723,
         Midori_rounds_n1722, Midori_rounds_n1721, Midori_rounds_n1720,
         Midori_rounds_n1719, Midori_rounds_n1718, Midori_rounds_n1717,
         Midori_rounds_n1716, Midori_rounds_n1715, Midori_rounds_n1714,
         Midori_rounds_n1713, Midori_rounds_n1712, Midori_rounds_n1711,
         Midori_rounds_n1710, Midori_rounds_n1709, Midori_rounds_n1708,
         Midori_rounds_n1707, Midori_rounds_n1706, Midori_rounds_n1705,
         Midori_rounds_n1704, Midori_rounds_n1703, Midori_rounds_n1702,
         Midori_rounds_n1701, Midori_rounds_n1700, Midori_rounds_n1699,
         Midori_rounds_n1698, Midori_rounds_n1697, Midori_rounds_n1696,
         Midori_rounds_n1695, Midori_rounds_n1694, Midori_rounds_n1693,
         Midori_rounds_n1692, Midori_rounds_n1691, Midori_rounds_n1690,
         Midori_rounds_n1689, Midori_rounds_n1688, Midori_rounds_n1687,
         Midori_rounds_n1686, Midori_rounds_n1685, Midori_rounds_n1684,
         Midori_rounds_n1683, Midori_rounds_n1682, Midori_rounds_n1681,
         Midori_rounds_n1680, Midori_rounds_n1679, Midori_rounds_n1678,
         Midori_rounds_n1677, Midori_rounds_n1676, Midori_rounds_n1675,
         Midori_rounds_n1674, Midori_rounds_n1673, Midori_rounds_n1672,
         Midori_rounds_n1671, Midori_rounds_n1670, Midori_rounds_n1669,
         Midori_rounds_n1668, Midori_rounds_n1667, Midori_rounds_n1666,
         Midori_rounds_n1665, Midori_rounds_n1664, Midori_rounds_n1663,
         Midori_rounds_n1662, Midori_rounds_n1661, Midori_rounds_n1660,
         Midori_rounds_n1659, Midori_rounds_n1658, Midori_rounds_n1657,
         Midori_rounds_n1656, Midori_rounds_n1655, Midori_rounds_n1654,
         Midori_rounds_n1653, Midori_rounds_n1652, Midori_rounds_n1651,
         Midori_rounds_n1650, Midori_rounds_n1649, Midori_rounds_n1648,
         Midori_rounds_n1647, Midori_rounds_n1646, Midori_rounds_n1645,
         Midori_rounds_n1644, Midori_rounds_n1643, Midori_rounds_n1642,
         Midori_rounds_n1641, Midori_rounds_n1640, Midori_rounds_n1639,
         Midori_rounds_n1638, Midori_rounds_n1637, Midori_rounds_n1636,
         Midori_rounds_n1635, Midori_rounds_n1634, Midori_rounds_n1633,
         Midori_rounds_n1632, Midori_rounds_n1631, Midori_rounds_n1630,
         Midori_rounds_n1629, Midori_rounds_n1628, Midori_rounds_n1627,
         Midori_rounds_n1626, Midori_rounds_n1625, Midori_rounds_n1624,
         Midori_rounds_n1623, Midori_rounds_n1622, Midori_rounds_n1621,
         Midori_rounds_n1620, Midori_rounds_n1619, Midori_rounds_n1618,
         Midori_rounds_n1617, Midori_rounds_n1616, Midori_rounds_n1615,
         Midori_rounds_n1614, Midori_rounds_n1613, Midori_rounds_n1612,
         Midori_rounds_n1611, Midori_rounds_n1610, Midori_rounds_n1609,
         Midori_rounds_n1608, Midori_rounds_n1607, Midori_rounds_n1606,
         Midori_rounds_n1605, Midori_rounds_n1604, Midori_rounds_n1603,
         Midori_rounds_n1602, Midori_rounds_n1601, Midori_rounds_n1600,
         Midori_rounds_n1599, Midori_rounds_n1598, Midori_rounds_n1597,
         Midori_rounds_n1596, Midori_rounds_n1595, Midori_rounds_n1594,
         Midori_rounds_n1593, Midori_rounds_n1592, Midori_rounds_n1591,
         Midori_rounds_n1590, Midori_rounds_n1589, Midori_rounds_n1588,
         Midori_rounds_n1587, Midori_rounds_n1586, Midori_rounds_n1585,
         Midori_rounds_n1584, Midori_rounds_n1583, Midori_rounds_n1582,
         Midori_rounds_n1581, Midori_rounds_n1580, Midori_rounds_n1579,
         Midori_rounds_n1578, Midori_rounds_n1577, Midori_rounds_n1576,
         Midori_rounds_n1575, Midori_rounds_n1574, Midori_rounds_n1573,
         Midori_rounds_n1572, Midori_rounds_n1571, Midori_rounds_n1570,
         Midori_rounds_n1569, Midori_rounds_n1568, Midori_rounds_n1567,
         Midori_rounds_n1566, Midori_rounds_n1565, Midori_rounds_n1564,
         Midori_rounds_n1563, Midori_rounds_n1562, Midori_rounds_n1561,
         Midori_rounds_n1560, Midori_rounds_n1559, Midori_rounds_n1558,
         Midori_rounds_n1557, Midori_rounds_n1556, Midori_rounds_n1555,
         Midori_rounds_n1554, Midori_rounds_n1553, Midori_rounds_n1552,
         Midori_rounds_n1551, Midori_rounds_n1550, Midori_rounds_n1549,
         Midori_rounds_n1548, Midori_rounds_n1547, Midori_rounds_n1546,
         Midori_rounds_n1545, Midori_rounds_n1544, Midori_rounds_n1543,
         Midori_rounds_n1542, Midori_rounds_n1541, Midori_rounds_n1540,
         Midori_rounds_n1539, Midori_rounds_n1538, Midori_rounds_n1537,
         Midori_rounds_n1536, Midori_rounds_n1535, Midori_rounds_n1534,
         Midori_rounds_n1533, Midori_rounds_n1532, Midori_rounds_n1531,
         Midori_rounds_n1530, Midori_rounds_n1529, Midori_rounds_n1528,
         Midori_rounds_n1527, Midori_rounds_n1526, Midori_rounds_n1525,
         Midori_rounds_n1524, Midori_rounds_n1523, Midori_rounds_n1522,
         Midori_rounds_n1521, Midori_rounds_n1520, Midori_rounds_n1519,
         Midori_rounds_n1518, Midori_rounds_n1517, Midori_rounds_n1516,
         Midori_rounds_n1515, Midori_rounds_n1514, Midori_rounds_n1513,
         Midori_rounds_n1512, Midori_rounds_n1511, Midori_rounds_n1510,
         Midori_rounds_n1509, Midori_rounds_n1508, Midori_rounds_n1507,
         Midori_rounds_n1506, Midori_rounds_n1505, Midori_rounds_n1504,
         Midori_rounds_n1503, Midori_rounds_n1502, Midori_rounds_n1501,
         Midori_rounds_n1500, Midori_rounds_n1499, Midori_rounds_n1498,
         Midori_rounds_n1497, Midori_rounds_n1496, Midori_rounds_n1495,
         Midori_rounds_n1494, Midori_rounds_n1493, Midori_rounds_n1492,
         Midori_rounds_n1491, Midori_rounds_n1490, Midori_rounds_n1489,
         Midori_rounds_n1488, Midori_rounds_n1487, Midori_rounds_n1486,
         Midori_rounds_n1485, Midori_rounds_n1484, Midori_rounds_n1483,
         Midori_rounds_n1482, Midori_rounds_n1481, Midori_rounds_n1480,
         Midori_rounds_n1479, Midori_rounds_n1478, Midori_rounds_n1477,
         Midori_rounds_n1476, Midori_rounds_n1475, Midori_rounds_n1474,
         Midori_rounds_n1473, Midori_rounds_n1472, Midori_rounds_n1471,
         Midori_rounds_n1470, Midori_rounds_n1469, Midori_rounds_n1468,
         Midori_rounds_n1467, Midori_rounds_n1466, Midori_rounds_n1465,
         Midori_rounds_n1464, Midori_rounds_n1463, Midori_rounds_n1462,
         Midori_rounds_n1461, Midori_rounds_n1460, Midori_rounds_n1459,
         Midori_rounds_n1458, Midori_rounds_n1457, Midori_rounds_n1456,
         Midori_rounds_n1455, Midori_rounds_n1454, Midori_rounds_n1453,
         Midori_rounds_n1452, Midori_rounds_n1451, Midori_rounds_n1450,
         Midori_rounds_n1449, Midori_rounds_n1448, Midori_rounds_n1447,
         Midori_rounds_n1446, Midori_rounds_n1445, Midori_rounds_n1444,
         Midori_rounds_n1443, Midori_rounds_n1442, Midori_rounds_n1441,
         Midori_rounds_n1440, Midori_rounds_n1439, Midori_rounds_n1438,
         Midori_rounds_n1437, Midori_rounds_n1436, Midori_rounds_n1435,
         Midori_rounds_n1434, Midori_rounds_n1433, Midori_rounds_n1432,
         Midori_rounds_n1431, Midori_rounds_n1430, Midori_rounds_n1429,
         Midori_rounds_n1428, Midori_rounds_n1427, Midori_rounds_n1426,
         Midori_rounds_n1425, Midori_rounds_n1424, Midori_rounds_n1423,
         Midori_rounds_n1422, Midori_rounds_n1421, Midori_rounds_n1420,
         Midori_rounds_n1419, Midori_rounds_n1418, Midori_rounds_n1417,
         Midori_rounds_n1416, Midori_rounds_n1415, Midori_rounds_n1414,
         Midori_rounds_n1413, Midori_rounds_n1412, Midori_rounds_n1411,
         Midori_rounds_n1410, Midori_rounds_n1409, Midori_rounds_n1408,
         Midori_rounds_n1407, Midori_rounds_n1406, Midori_rounds_n1405,
         Midori_rounds_n1404, Midori_rounds_n1403, Midori_rounds_n1402,
         Midori_rounds_n1401, Midori_rounds_n1400, Midori_rounds_n1399,
         Midori_rounds_n1398, Midori_rounds_n1397, Midori_rounds_n1396,
         Midori_rounds_n1395, Midori_rounds_n1394, Midori_rounds_n1393,
         Midori_rounds_n1392, Midori_rounds_n1391, Midori_rounds_n1390,
         Midori_rounds_n1389, Midori_rounds_n1388, Midori_rounds_n1387,
         Midori_rounds_n1386, Midori_rounds_n1385, Midori_rounds_n1384,
         Midori_rounds_n1383, Midori_rounds_n1382, Midori_rounds_n1381,
         Midori_rounds_n1380, Midori_rounds_n1379, Midori_rounds_n1378,
         Midori_rounds_n1377, Midori_rounds_n1376, Midori_rounds_n1375,
         Midori_rounds_n1374, Midori_rounds_n1373, Midori_rounds_n1372,
         Midori_rounds_n1371, Midori_rounds_n1370, Midori_rounds_n1369,
         Midori_rounds_n1368, Midori_rounds_n1367, Midori_rounds_n1366,
         Midori_rounds_n1365, Midori_rounds_n1364, Midori_rounds_n1363,
         Midori_rounds_n1362, Midori_rounds_n1361, Midori_rounds_n1360,
         Midori_rounds_n1359, Midori_rounds_n1358, Midori_rounds_n1357,
         Midori_rounds_n1356, Midori_rounds_n1355, Midori_rounds_n1354,
         Midori_rounds_n1353, Midori_rounds_n1352, Midori_rounds_n1351,
         Midori_rounds_n1350, Midori_rounds_n1349, Midori_rounds_n1348,
         Midori_rounds_n1347, Midori_rounds_n1346, Midori_rounds_n1345,
         Midori_rounds_n1344, Midori_rounds_n1343, Midori_rounds_n1342,
         Midori_rounds_n1341, Midori_rounds_n1340, Midori_rounds_n1339,
         Midori_rounds_n1338, Midori_rounds_n1337, Midori_rounds_n1336,
         Midori_rounds_n1335, Midori_rounds_n1334, Midori_rounds_n1333,
         Midori_rounds_n1332, Midori_rounds_n1331, Midori_rounds_n1330,
         Midori_rounds_n1329, Midori_rounds_n1328, Midori_rounds_n1327,
         Midori_rounds_n1326, Midori_rounds_n1325, Midori_rounds_n1324,
         Midori_rounds_n1323, Midori_rounds_n1322, Midori_rounds_n1321,
         Midori_rounds_n1320, Midori_rounds_n1319, Midori_rounds_n1318,
         Midori_rounds_n1317, Midori_rounds_n1316, Midori_rounds_n1315,
         Midori_rounds_n1314, Midori_rounds_n1313, Midori_rounds_n1312,
         Midori_rounds_n1311, Midori_rounds_n1310, Midori_rounds_n1309,
         Midori_rounds_n1308, Midori_rounds_n1307, Midori_rounds_n1306,
         Midori_rounds_n1305, Midori_rounds_n1304, Midori_rounds_n1303,
         Midori_rounds_n1302, Midori_rounds_n1301, Midori_rounds_n1300,
         Midori_rounds_n1299, Midori_rounds_n1298, Midori_rounds_n1297,
         Midori_rounds_n1296, Midori_rounds_n1295, Midori_rounds_n1294,
         Midori_rounds_n1293, Midori_rounds_n1292, Midori_rounds_n1291,
         Midori_rounds_n1290, Midori_rounds_n1289, Midori_rounds_n1288,
         Midori_rounds_n1287, Midori_rounds_n1286, Midori_rounds_n1285,
         Midori_rounds_n1284, Midori_rounds_n1283, Midori_rounds_n1282,
         Midori_rounds_n1281, Midori_rounds_n1280, Midori_rounds_n1279,
         Midori_rounds_n1278, Midori_rounds_n1277, Midori_rounds_n1276,
         Midori_rounds_n1275, Midori_rounds_n1274, Midori_rounds_n1273,
         Midori_rounds_n1272, Midori_rounds_n1271, Midori_rounds_n1270,
         Midori_rounds_n1269, Midori_rounds_n1268, Midori_rounds_n1267,
         Midori_rounds_n1266, Midori_rounds_n1265, Midori_rounds_n1264,
         Midori_rounds_n1263, Midori_rounds_n1262, Midori_rounds_n1261,
         Midori_rounds_n1260, Midori_rounds_n1259, Midori_rounds_n1258,
         Midori_rounds_n1257, Midori_rounds_n1256, Midori_rounds_n1255,
         Midori_rounds_n1254, Midori_rounds_n1253, Midori_rounds_n1252,
         Midori_rounds_n1251, Midori_rounds_n1250, Midori_rounds_n1249,
         Midori_rounds_n1248, Midori_rounds_n1247, Midori_rounds_n1246,
         Midori_rounds_n1245, Midori_rounds_n1244, Midori_rounds_n1243,
         Midori_rounds_n1242, Midori_rounds_n1241, Midori_rounds_n979,
         Midori_rounds_n977, Midori_rounds_n975, Midori_rounds_n973,
         Midori_rounds_n971, Midori_rounds_n969, Midori_rounds_n967,
         Midori_rounds_n965, Midori_rounds_n963, Midori_rounds_n961,
         Midori_rounds_n959, Midori_rounds_n957, Midori_rounds_n955,
         Midori_rounds_n953, Midori_rounds_n951, Midori_rounds_n949,
         Midori_rounds_n947, Midori_rounds_n945, Midori_rounds_n943,
         Midori_rounds_n941, Midori_rounds_n939, Midori_rounds_n937,
         Midori_rounds_n935, Midori_rounds_n933, Midori_rounds_n931,
         Midori_rounds_n929, Midori_rounds_n927, Midori_rounds_n925,
         Midori_rounds_n923, Midori_rounds_n921, Midori_rounds_n919,
         Midori_rounds_n917, Midori_rounds_n915, Midori_rounds_n913,
         Midori_rounds_n911, Midori_rounds_n909, Midori_rounds_n907,
         Midori_rounds_n905, Midori_rounds_n903, Midori_rounds_n901,
         Midori_rounds_n899, Midori_rounds_n897, Midori_rounds_n895,
         Midori_rounds_n893, Midori_rounds_n891, Midori_rounds_n889,
         Midori_rounds_n887, Midori_rounds_n885, Midori_rounds_n883,
         Midori_rounds_n881, Midori_rounds_n879, Midori_rounds_n877,
         Midori_rounds_n875, Midori_rounds_n873, Midori_rounds_n871,
         Midori_rounds_n869, Midori_rounds_n867, Midori_rounds_n865,
         Midori_rounds_n863, Midori_rounds_n861, Midori_rounds_n859,
         Midori_rounds_n857, Midori_rounds_n855, Midori_rounds_n853,
         Midori_rounds_n851, Midori_rounds_n850, Midori_rounds_n848,
         Midori_rounds_n847, Midori_rounds_n845, Midori_rounds_n844,
         Midori_rounds_n842, Midori_rounds_n841, Midori_rounds_n839,
         Midori_rounds_n838, Midori_rounds_n836, Midori_rounds_n835,
         Midori_rounds_n833, Midori_rounds_n832, Midori_rounds_n830,
         Midori_rounds_n829, Midori_rounds_n827, Midori_rounds_n826,
         Midori_rounds_n824, Midori_rounds_n823, Midori_rounds_n821,
         Midori_rounds_n820, Midori_rounds_n818, Midori_rounds_n817,
         Midori_rounds_n815, Midori_rounds_n814, Midori_rounds_n812,
         Midori_rounds_n811, Midori_rounds_n809, Midori_rounds_n808,
         Midori_rounds_n806, Midori_rounds_n805, Midori_rounds_n804,
         Midori_rounds_n803, Midori_rounds_n802, Midori_rounds_n801,
         Midori_rounds_n800, Midori_rounds_n799, Midori_rounds_n798,
         Midori_rounds_n797, Midori_rounds_n796, Midori_rounds_n795,
         Midori_rounds_n794, Midori_rounds_n793, Midori_rounds_n792,
         Midori_rounds_n791, Midori_rounds_n790, Midori_rounds_n789,
         Midori_rounds_constant_MUX_n70, Midori_rounds_constant_MUX_n69,
         Midori_rounds_constant_MUX_n68, Midori_rounds_constant_MUX_n67,
         Midori_rounds_constant_MUX_n66, Midori_rounds_constant_MUX_n65,
         Midori_rounds_constant_MUX_n64, Midori_rounds_constant_MUX_n63,
         Midori_rounds_constant_MUX_n62, Midori_rounds_constant_MUX_n61,
         Midori_rounds_constant_MUX_n60, Midori_rounds_constant_MUX_n59,
         Midori_rounds_constant_MUX_n58, Midori_rounds_constant_MUX_n57,
         Midori_rounds_constant_MUX_n56, Midori_rounds_constant_MUX_n55,
         Midori_rounds_constant_MUX_n54, Midori_rounds_constant_MUX_n53,
         Midori_rounds_constant_MUX_n52, Midori_rounds_constant_MUX_n51,
         Midori_rounds_constant_MUX_n50, Midori_rounds_constant_MUX_n49,
         Midori_rounds_constant_MUX_n48, Midori_rounds_constant_MUX_n47,
         Midori_rounds_constant_MUX_n46, Midori_rounds_constant_MUX_n45,
         Midori_rounds_constant_MUX_n44, Midori_rounds_constant_MUX_n43,
         Midori_rounds_constant_MUX_n42, Midori_rounds_constant_MUX_n41,
         Midori_rounds_constant_MUX_n40, Midori_rounds_constant_MUX_n39,
         Midori_rounds_constant_MUX_n38, Midori_rounds_constant_MUX_n37,
         Midori_rounds_constant_MUX_n36, Midori_rounds_constant_MUX_n35,
         Midori_rounds_constant_MUX_n34, Midori_rounds_constant_MUX_n33,
         Midori_rounds_constant_MUX_n32, Midori_rounds_constant_MUX_n31,
         Midori_rounds_constant_MUX_n30, Midori_rounds_constant_MUX_n29,
         Midori_rounds_constant_MUX_n28, Midori_rounds_constant_MUX_n27,
         Midori_rounds_constant_MUX_n26, Midori_rounds_constant_MUX_n25,
         Midori_rounds_constant_MUX_n24, Midori_rounds_constant_MUX_n23,
         Midori_rounds_constant_MUX_n22, Midori_rounds_constant_MUX_n21,
         Midori_rounds_constant_MUX_n20, Midori_rounds_constant_MUX_n19,
         Midori_rounds_constant_MUX_n18, Midori_rounds_constant_MUX_n17,
         Midori_rounds_constant_MUX_n16, Midori_rounds_constant_MUX_n15,
         Midori_rounds_constant_MUX_n14, Midori_rounds_constant_MUX_n13,
         Midori_rounds_constant_MUX_n12, Midori_rounds_constant_MUX_n11,
         Midori_rounds_constant_MUX_n10, Midori_rounds_sub_Sub_0_F_n4,
         Midori_rounds_sub_Sub_0_F_n3, Midori_rounds_sub_Sub_0_F_n2,
         Midori_rounds_sub_Sub_0_F_n1,
         Midori_rounds_sub_Sub_0_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_0_G_n1,
         Midori_rounds_sub_Sub_0_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_0_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_1_F_n12, Midori_rounds_sub_Sub_1_F_n11,
         Midori_rounds_sub_Sub_1_F_n10, Midori_rounds_sub_Sub_1_F_n9,
         Midori_rounds_sub_Sub_1_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_1_G_n1,
         Midori_rounds_sub_Sub_1_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_1_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_2_F_n12, Midori_rounds_sub_Sub_2_F_n11,
         Midori_rounds_sub_Sub_2_F_n10, Midori_rounds_sub_Sub_2_F_n9,
         Midori_rounds_sub_Sub_2_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_2_G_n1,
         Midori_rounds_sub_Sub_2_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_2_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_3_F_n12, Midori_rounds_sub_Sub_3_F_n11,
         Midori_rounds_sub_Sub_3_F_n10, Midori_rounds_sub_Sub_3_F_n9,
         Midori_rounds_sub_Sub_3_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_3_G_n1,
         Midori_rounds_sub_Sub_3_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_3_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_4_F_n12, Midori_rounds_sub_Sub_4_F_n11,
         Midori_rounds_sub_Sub_4_F_n10, Midori_rounds_sub_Sub_4_F_n9,
         Midori_rounds_sub_Sub_4_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_4_G_n1,
         Midori_rounds_sub_Sub_4_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_4_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_5_F_n12, Midori_rounds_sub_Sub_5_F_n11,
         Midori_rounds_sub_Sub_5_F_n10, Midori_rounds_sub_Sub_5_F_n9,
         Midori_rounds_sub_Sub_5_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_5_G_n1,
         Midori_rounds_sub_Sub_5_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_5_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_6_F_n12, Midori_rounds_sub_Sub_6_F_n11,
         Midori_rounds_sub_Sub_6_F_n10, Midori_rounds_sub_Sub_6_F_n9,
         Midori_rounds_sub_Sub_6_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_6_G_n1,
         Midori_rounds_sub_Sub_6_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_6_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_7_F_n12, Midori_rounds_sub_Sub_7_F_n11,
         Midori_rounds_sub_Sub_7_F_n10, Midori_rounds_sub_Sub_7_F_n9,
         Midori_rounds_sub_Sub_7_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_7_G_n1,
         Midori_rounds_sub_Sub_7_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_7_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_8_F_n12, Midori_rounds_sub_Sub_8_F_n11,
         Midori_rounds_sub_Sub_8_F_n10, Midori_rounds_sub_Sub_8_F_n9,
         Midori_rounds_sub_Sub_8_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_8_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_8_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_8_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_8_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_8_G_n1,
         Midori_rounds_sub_Sub_8_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_8_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_8_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_8_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_9_F_n12, Midori_rounds_sub_Sub_9_F_n11,
         Midori_rounds_sub_Sub_9_F_n10, Midori_rounds_sub_Sub_9_F_n9,
         Midori_rounds_sub_Sub_9_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_9_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_9_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_9_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_9_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_9_G_n1,
         Midori_rounds_sub_Sub_9_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_9_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_9_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_9_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_10_F_n12, Midori_rounds_sub_Sub_10_F_n11,
         Midori_rounds_sub_Sub_10_F_n10, Midori_rounds_sub_Sub_10_F_n9,
         Midori_rounds_sub_Sub_10_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_10_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_10_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_10_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_10_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_10_G_n2,
         Midori_rounds_sub_Sub_10_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_10_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_10_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_10_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_11_F_n12, Midori_rounds_sub_Sub_11_F_n11,
         Midori_rounds_sub_Sub_11_F_n10, Midori_rounds_sub_Sub_11_F_n9,
         Midori_rounds_sub_Sub_11_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_11_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_11_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_11_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_11_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_11_G_n1,
         Midori_rounds_sub_Sub_11_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_11_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_11_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_11_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_12_F_n12, Midori_rounds_sub_Sub_12_F_n11,
         Midori_rounds_sub_Sub_12_F_n10, Midori_rounds_sub_Sub_12_F_n9,
         Midori_rounds_sub_Sub_12_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_12_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_12_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_12_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_12_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_12_G_n1,
         Midori_rounds_sub_Sub_12_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_12_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_12_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_12_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_13_F_n12, Midori_rounds_sub_Sub_13_F_n11,
         Midori_rounds_sub_Sub_13_F_n10, Midori_rounds_sub_Sub_13_F_n9,
         Midori_rounds_sub_Sub_13_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_13_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_13_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_13_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_13_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_13_G_n1,
         Midori_rounds_sub_Sub_13_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_13_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_13_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_13_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_14_F_n12, Midori_rounds_sub_Sub_14_F_n11,
         Midori_rounds_sub_Sub_14_F_n10, Midori_rounds_sub_Sub_14_F_n9,
         Midori_rounds_sub_Sub_14_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_14_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_14_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_14_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_14_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_14_G_n1,
         Midori_rounds_sub_Sub_14_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_14_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_14_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_14_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_sub_Sub_15_F_n12, Midori_rounds_sub_Sub_15_F_n11,
         Midori_rounds_sub_Sub_15_F_n10, Midori_rounds_sub_Sub_15_F_n9,
         Midori_rounds_sub_Sub_15_F_Inst_1__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_4__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_5__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_n6,
         Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_n5,
         Midori_rounds_sub_Sub_15_F_Inst_9__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_n5,
         Midori_rounds_sub_Sub_15_F_Inst_11__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_15_F_Inst_13__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_15__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_F_Inst_17__CF_Inst_n6,
         Midori_rounds_sub_Sub_15_F_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_n10,
         Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_F_Inst_22__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_26__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_n8,
         Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_n4,
         Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_n10,
         Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_n10,
         Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_F_Inst_31__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_32__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n11,
         Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n10,
         Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_n4,
         Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression1_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression2_n3,
         Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression3_n3,
         Midori_rounds_sub_Sub_15_G_n1,
         Midori_rounds_sub_Sub_15_G_Inst_0__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_G_Inst_1__CF_Inst_n6,
         Midori_rounds_sub_Sub_15_G_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_6__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_G_Inst_7__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_G_Inst_8__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_10__CF_Inst_n6,
         Midori_rounds_sub_Sub_15_G_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_14__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_G_Inst_16__CF_Inst_n2,
         Midori_rounds_sub_Sub_15_G_Inst_17__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_18__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_n4,
         Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_20__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_n4,
         Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_G_Inst_23__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_n4,
         Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_n3,
         Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_n10,
         Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_n9,
         Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression1_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression2_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression3_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression1_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression2_n3,
         Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression3_n3,
         Midori_rounds_mul1_MC1_n24, Midori_rounds_mul1_MC1_n23,
         Midori_rounds_mul1_MC1_n22, Midori_rounds_mul1_MC1_n21,
         Midori_rounds_mul1_MC1_n20, Midori_rounds_mul1_MC1_n19,
         Midori_rounds_mul1_MC1_n18, Midori_rounds_mul1_MC1_n17,
         Midori_rounds_mul1_MC2_n24, Midori_rounds_mul1_MC2_n23,
         Midori_rounds_mul1_MC2_n22, Midori_rounds_mul1_MC2_n21,
         Midori_rounds_mul1_MC2_n20, Midori_rounds_mul1_MC2_n19,
         Midori_rounds_mul1_MC2_n18, Midori_rounds_mul1_MC2_n17,
         Midori_rounds_mul1_MC3_n24, Midori_rounds_mul1_MC3_n23,
         Midori_rounds_mul1_MC3_n22, Midori_rounds_mul1_MC3_n21,
         Midori_rounds_mul1_MC3_n20, Midori_rounds_mul1_MC3_n19,
         Midori_rounds_mul1_MC3_n18, Midori_rounds_mul1_MC3_n17,
         Midori_rounds_mul1_MC4_n24, Midori_rounds_mul1_MC4_n23,
         Midori_rounds_mul1_MC4_n22, Midori_rounds_mul1_MC4_n21,
         Midori_rounds_mul1_MC4_n20, Midori_rounds_mul1_MC4_n19,
         Midori_rounds_mul1_MC4_n18, Midori_rounds_mul1_MC4_n17,
         Midori_rounds_mul2_MC1_n24, Midori_rounds_mul2_MC1_n23,
         Midori_rounds_mul2_MC1_n22, Midori_rounds_mul2_MC1_n21,
         Midori_rounds_mul2_MC1_n20, Midori_rounds_mul2_MC1_n19,
         Midori_rounds_mul2_MC1_n18, Midori_rounds_mul2_MC1_n17,
         Midori_rounds_mul2_MC2_n24, Midori_rounds_mul2_MC2_n23,
         Midori_rounds_mul2_MC2_n22, Midori_rounds_mul2_MC2_n21,
         Midori_rounds_mul2_MC2_n20, Midori_rounds_mul2_MC2_n19,
         Midori_rounds_mul2_MC2_n18, Midori_rounds_mul2_MC2_n17,
         Midori_rounds_mul2_MC3_n24, Midori_rounds_mul2_MC3_n23,
         Midori_rounds_mul2_MC3_n22, Midori_rounds_mul2_MC3_n21,
         Midori_rounds_mul2_MC3_n20, Midori_rounds_mul2_MC3_n19,
         Midori_rounds_mul2_MC3_n18, Midori_rounds_mul2_MC3_n17,
         Midori_rounds_mul2_MC4_n24, Midori_rounds_mul2_MC4_n23,
         Midori_rounds_mul2_MC4_n22, Midori_rounds_mul2_MC4_n21,
         Midori_rounds_mul2_MC4_n20, Midori_rounds_mul2_MC4_n19,
         Midori_rounds_mul2_MC4_n18, Midori_rounds_mul2_MC4_n17,
         Midori_rounds_mul3_MC1_n24, Midori_rounds_mul3_MC1_n23,
         Midori_rounds_mul3_MC1_n22, Midori_rounds_mul3_MC1_n21,
         Midori_rounds_mul3_MC1_n20, Midori_rounds_mul3_MC1_n19,
         Midori_rounds_mul3_MC1_n18, Midori_rounds_mul3_MC1_n17,
         Midori_rounds_mul3_MC2_n24, Midori_rounds_mul3_MC2_n23,
         Midori_rounds_mul3_MC2_n22, Midori_rounds_mul3_MC2_n21,
         Midori_rounds_mul3_MC2_n20, Midori_rounds_mul3_MC2_n19,
         Midori_rounds_mul3_MC2_n18, Midori_rounds_mul3_MC2_n17,
         Midori_rounds_mul3_MC3_n24, Midori_rounds_mul3_MC3_n23,
         Midori_rounds_mul3_MC3_n22, Midori_rounds_mul3_MC3_n21,
         Midori_rounds_mul3_MC3_n20, Midori_rounds_mul3_MC3_n19,
         Midori_rounds_mul3_MC3_n18, Midori_rounds_mul3_MC3_n17,
         Midori_rounds_mul3_MC4_n24, Midori_rounds_mul3_MC4_n23,
         Midori_rounds_mul3_MC4_n22, Midori_rounds_mul3_MC4_n21,
         Midori_rounds_mul3_MC4_n20, Midori_rounds_mul3_MC4_n19,
         Midori_rounds_mul3_MC4_n18, Midori_rounds_mul3_MC4_n17;
  wire   [63:0] wk_share1;
  wire   [63:0] wk_share2;
  wire   [63:0] wk_share3;
  wire   [3:0] round_Signal;
  wire   [63:0] Midori_add_Result_Start3;
  wire   [63:0] Midori_add_Result_Start2;
  wire   [63:0] Midori_add_Result_Start1;
  wire   [63:0] Midori_rounds_SR_Inv_Result3;
  wire   [63:0] Midori_rounds_SR_Inv_Result2;
  wire   [63:0] Midori_rounds_SR_Inv_Result1;
  wire   [63:0] Midori_rounds_mul_input3;
  wire   [63:0] Midori_rounds_mul_input2;
  wire   [63:0] Midori_rounds_mul_input1;
  wire   [63:0] Midori_rounds_SR_Result3;
  wire   [63:0] Midori_rounds_SR_Result2;
  wire   [63:0] Midori_rounds_SR_Result1;
  wire   [15:0] Midori_rounds_round_Constant;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_0_q3;
  wire   [3:0] Midori_rounds_sub_Sub_0_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_0_q2;
  wire   [3:0] Midori_rounds_sub_Sub_0_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_0_q1;
  wire   [3:0] Midori_rounds_sub_Sub_0_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_0_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_0_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_0_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_0_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_0_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_1_q3;
  wire   [3:0] Midori_rounds_sub_Sub_1_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_1_q2;
  wire   [3:0] Midori_rounds_sub_Sub_1_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_1_q1;
  wire   [3:0] Midori_rounds_sub_Sub_1_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_1_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_1_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_1_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_1_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_1_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_2_q3;
  wire   [3:0] Midori_rounds_sub_Sub_2_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_2_q2;
  wire   [3:0] Midori_rounds_sub_Sub_2_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_2_q1;
  wire   [3:0] Midori_rounds_sub_Sub_2_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_2_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_2_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_2_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_2_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_2_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_3_q3;
  wire   [3:0] Midori_rounds_sub_Sub_3_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_3_q2;
  wire   [3:0] Midori_rounds_sub_Sub_3_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_3_q1;
  wire   [3:0] Midori_rounds_sub_Sub_3_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_3_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_3_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_3_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_3_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_3_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_4_q3;
  wire   [3:0] Midori_rounds_sub_Sub_4_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_4_q2;
  wire   [3:0] Midori_rounds_sub_Sub_4_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_4_q1;
  wire   [3:0] Midori_rounds_sub_Sub_4_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_4_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_4_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_4_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_4_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_4_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_5_q3;
  wire   [3:0] Midori_rounds_sub_Sub_5_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_5_q2;
  wire   [3:0] Midori_rounds_sub_Sub_5_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_5_q1;
  wire   [3:0] Midori_rounds_sub_Sub_5_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_5_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_5_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_5_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_5_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_5_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_6_q3;
  wire   [3:0] Midori_rounds_sub_Sub_6_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_6_q2;
  wire   [3:0] Midori_rounds_sub_Sub_6_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_6_q1;
  wire   [3:0] Midori_rounds_sub_Sub_6_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_6_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_6_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_6_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_6_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_6_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_7_q3;
  wire   [3:0] Midori_rounds_sub_Sub_7_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_7_q2;
  wire   [3:0] Midori_rounds_sub_Sub_7_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_7_q1;
  wire   [3:0] Midori_rounds_sub_Sub_7_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_7_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_7_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_7_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_7_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_7_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_8_q3;
  wire   [3:0] Midori_rounds_sub_Sub_8_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_8_q2;
  wire   [3:0] Midori_rounds_sub_Sub_8_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_8_q1;
  wire   [3:0] Midori_rounds_sub_Sub_8_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_8_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_8_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_8_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_8_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_8_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_9_q3;
  wire   [3:0] Midori_rounds_sub_Sub_9_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_9_q2;
  wire   [3:0] Midori_rounds_sub_Sub_9_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_9_q1;
  wire   [3:0] Midori_rounds_sub_Sub_9_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_9_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_9_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_9_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_9_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_9_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_10_q3;
  wire   [3:0] Midori_rounds_sub_Sub_10_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_10_q2;
  wire   [3:0] Midori_rounds_sub_Sub_10_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_10_q1;
  wire   [3:0] Midori_rounds_sub_Sub_10_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_10_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_10_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_10_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_10_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_10_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_11_q3;
  wire   [3:0] Midori_rounds_sub_Sub_11_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_11_q2;
  wire   [3:0] Midori_rounds_sub_Sub_11_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_11_q1;
  wire   [3:0] Midori_rounds_sub_Sub_11_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_11_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_11_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_11_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_11_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_11_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_12_q3;
  wire   [3:0] Midori_rounds_sub_Sub_12_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_12_q2;
  wire   [3:0] Midori_rounds_sub_Sub_12_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_12_q1;
  wire   [3:0] Midori_rounds_sub_Sub_12_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_12_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_12_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_12_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_12_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_12_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_13_q3;
  wire   [3:0] Midori_rounds_sub_Sub_13_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_13_q2;
  wire   [3:0] Midori_rounds_sub_Sub_13_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_13_q1;
  wire   [3:0] Midori_rounds_sub_Sub_13_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_13_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_13_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_13_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_13_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_13_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_14_q3;
  wire   [3:0] Midori_rounds_sub_Sub_14_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_14_q2;
  wire   [3:0] Midori_rounds_sub_Sub_14_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_14_q1;
  wire   [3:0] Midori_rounds_sub_Sub_14_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_14_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_14_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_14_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_14_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_14_G_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_in3;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_in3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_in2;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_in2_reg;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_in1;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_in1_reg;
  wire   [3:0] Midori_rounds_sub_Sub_15_q3;
  wire   [3:0] Midori_rounds_sub_Sub_15_Rq3;
  wire   [3:0] Midori_rounds_sub_Sub_15_q2;
  wire   [3:0] Midori_rounds_sub_Sub_15_Rq2;
  wire   [3:0] Midori_rounds_sub_Sub_15_q1;
  wire   [3:0] Midori_rounds_sub_Sub_15_Rq1;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_q3;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_q2;
  wire   [3:0] Midori_rounds_sub_Sub_15_F_q1;
  wire   [35:0] Midori_rounds_sub_Sub_15_F_CF_Reg;
  wire   [35:0] Midori_rounds_sub_Sub_15_F_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_15_G_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_15_G_CF_Out;

  XOR2_X1 KeySchadule1_U64 ( .A(Key1[73]), .B(Key1[9]), .Z(wk_share1[9]) );
  XOR2_X1 KeySchadule1_U63 ( .A(Key1[72]), .B(Key1[8]), .Z(wk_share1[8]) );
  XOR2_X1 KeySchadule1_U62 ( .A(Key1[71]), .B(Key1[7]), .Z(wk_share1[7]) );
  XOR2_X1 KeySchadule1_U61 ( .A(Key1[6]), .B(Key1[70]), .Z(wk_share1[6]) );
  XOR2_X1 KeySchadule1_U60 ( .A(Key1[127]), .B(Key1[63]), .Z(wk_share1[63]) );
  XOR2_X1 KeySchadule1_U59 ( .A(Key1[126]), .B(Key1[62]), .Z(wk_share1[62]) );
  XOR2_X1 KeySchadule1_U58 ( .A(Key1[125]), .B(Key1[61]), .Z(wk_share1[61]) );
  XOR2_X1 KeySchadule1_U57 ( .A(Key1[124]), .B(Key1[60]), .Z(wk_share1[60]) );
  XOR2_X1 KeySchadule1_U56 ( .A(Key1[5]), .B(Key1[69]), .Z(wk_share1[5]) );
  XOR2_X1 KeySchadule1_U55 ( .A(Key1[123]), .B(Key1[59]), .Z(wk_share1[59]) );
  XOR2_X1 KeySchadule1_U54 ( .A(Key1[122]), .B(Key1[58]), .Z(wk_share1[58]) );
  XOR2_X1 KeySchadule1_U53 ( .A(Key1[121]), .B(Key1[57]), .Z(wk_share1[57]) );
  XOR2_X1 KeySchadule1_U52 ( .A(Key1[120]), .B(Key1[56]), .Z(wk_share1[56]) );
  XOR2_X1 KeySchadule1_U51 ( .A(Key1[119]), .B(Key1[55]), .Z(wk_share1[55]) );
  XOR2_X1 KeySchadule1_U50 ( .A(Key1[118]), .B(Key1[54]), .Z(wk_share1[54]) );
  XOR2_X1 KeySchadule1_U49 ( .A(Key1[117]), .B(Key1[53]), .Z(wk_share1[53]) );
  XOR2_X1 KeySchadule1_U48 ( .A(Key1[116]), .B(Key1[52]), .Z(wk_share1[52]) );
  XOR2_X1 KeySchadule1_U47 ( .A(Key1[115]), .B(Key1[51]), .Z(wk_share1[51]) );
  XOR2_X1 KeySchadule1_U46 ( .A(Key1[114]), .B(Key1[50]), .Z(wk_share1[50]) );
  XOR2_X1 KeySchadule1_U45 ( .A(Key1[4]), .B(Key1[68]), .Z(wk_share1[4]) );
  XOR2_X1 KeySchadule1_U44 ( .A(Key1[113]), .B(Key1[49]), .Z(wk_share1[49]) );
  XOR2_X1 KeySchadule1_U43 ( .A(Key1[112]), .B(Key1[48]), .Z(wk_share1[48]) );
  XOR2_X1 KeySchadule1_U42 ( .A(Key1[111]), .B(Key1[47]), .Z(wk_share1[47]) );
  XOR2_X1 KeySchadule1_U41 ( .A(Key1[110]), .B(Key1[46]), .Z(wk_share1[46]) );
  XOR2_X1 KeySchadule1_U40 ( .A(Key1[109]), .B(Key1[45]), .Z(wk_share1[45]) );
  XOR2_X1 KeySchadule1_U39 ( .A(Key1[108]), .B(Key1[44]), .Z(wk_share1[44]) );
  XOR2_X1 KeySchadule1_U38 ( .A(Key1[107]), .B(Key1[43]), .Z(wk_share1[43]) );
  XOR2_X1 KeySchadule1_U37 ( .A(Key1[106]), .B(Key1[42]), .Z(wk_share1[42]) );
  XOR2_X1 KeySchadule1_U36 ( .A(Key1[105]), .B(Key1[41]), .Z(wk_share1[41]) );
  XOR2_X1 KeySchadule1_U35 ( .A(Key1[104]), .B(Key1[40]), .Z(wk_share1[40]) );
  XOR2_X1 KeySchadule1_U34 ( .A(Key1[3]), .B(Key1[67]), .Z(wk_share1[3]) );
  XOR2_X1 KeySchadule1_U33 ( .A(Key1[103]), .B(Key1[39]), .Z(wk_share1[39]) );
  XOR2_X1 KeySchadule1_U32 ( .A(Key1[102]), .B(Key1[38]), .Z(wk_share1[38]) );
  XOR2_X1 KeySchadule1_U31 ( .A(Key1[101]), .B(Key1[37]), .Z(wk_share1[37]) );
  XOR2_X1 KeySchadule1_U30 ( .A(Key1[100]), .B(Key1[36]), .Z(wk_share1[36]) );
  XOR2_X1 KeySchadule1_U29 ( .A(Key1[35]), .B(Key1[99]), .Z(wk_share1[35]) );
  XOR2_X1 KeySchadule1_U28 ( .A(Key1[34]), .B(Key1[98]), .Z(wk_share1[34]) );
  XOR2_X1 KeySchadule1_U27 ( .A(Key1[33]), .B(Key1[97]), .Z(wk_share1[33]) );
  XOR2_X1 KeySchadule1_U26 ( .A(Key1[32]), .B(Key1[96]), .Z(wk_share1[32]) );
  XOR2_X1 KeySchadule1_U25 ( .A(Key1[31]), .B(Key1[95]), .Z(wk_share1[31]) );
  XOR2_X1 KeySchadule1_U24 ( .A(Key1[30]), .B(Key1[94]), .Z(wk_share1[30]) );
  XOR2_X1 KeySchadule1_U23 ( .A(Key1[2]), .B(Key1[66]), .Z(wk_share1[2]) );
  XOR2_X1 KeySchadule1_U22 ( .A(Key1[29]), .B(Key1[93]), .Z(wk_share1[29]) );
  XOR2_X1 KeySchadule1_U21 ( .A(Key1[28]), .B(Key1[92]), .Z(wk_share1[28]) );
  XOR2_X1 KeySchadule1_U20 ( .A(Key1[27]), .B(Key1[91]), .Z(wk_share1[27]) );
  XOR2_X1 KeySchadule1_U19 ( .A(Key1[26]), .B(Key1[90]), .Z(wk_share1[26]) );
  XOR2_X1 KeySchadule1_U18 ( .A(Key1[25]), .B(Key1[89]), .Z(wk_share1[25]) );
  XOR2_X1 KeySchadule1_U17 ( .A(Key1[24]), .B(Key1[88]), .Z(wk_share1[24]) );
  XOR2_X1 KeySchadule1_U16 ( .A(Key1[23]), .B(Key1[87]), .Z(wk_share1[23]) );
  XOR2_X1 KeySchadule1_U15 ( .A(Key1[22]), .B(Key1[86]), .Z(wk_share1[22]) );
  XOR2_X1 KeySchadule1_U14 ( .A(Key1[21]), .B(Key1[85]), .Z(wk_share1[21]) );
  XOR2_X1 KeySchadule1_U13 ( .A(Key1[20]), .B(Key1[84]), .Z(wk_share1[20]) );
  XOR2_X1 KeySchadule1_U12 ( .A(Key1[1]), .B(Key1[65]), .Z(wk_share1[1]) );
  XOR2_X1 KeySchadule1_U11 ( .A(Key1[19]), .B(Key1[83]), .Z(wk_share1[19]) );
  XOR2_X1 KeySchadule1_U10 ( .A(Key1[18]), .B(Key1[82]), .Z(wk_share1[18]) );
  XOR2_X1 KeySchadule1_U9 ( .A(Key1[17]), .B(Key1[81]), .Z(wk_share1[17]) );
  XOR2_X1 KeySchadule1_U8 ( .A(Key1[16]), .B(Key1[80]), .Z(wk_share1[16]) );
  XOR2_X1 KeySchadule1_U7 ( .A(Key1[15]), .B(Key1[79]), .Z(wk_share1[15]) );
  XOR2_X1 KeySchadule1_U6 ( .A(Key1[14]), .B(Key1[78]), .Z(wk_share1[14]) );
  XOR2_X1 KeySchadule1_U5 ( .A(Key1[13]), .B(Key1[77]), .Z(wk_share1[13]) );
  XOR2_X1 KeySchadule1_U4 ( .A(Key1[12]), .B(Key1[76]), .Z(wk_share1[12]) );
  XOR2_X1 KeySchadule1_U3 ( .A(Key1[11]), .B(Key1[75]), .Z(wk_share1[11]) );
  XOR2_X1 KeySchadule1_U2 ( .A(Key1[10]), .B(Key1[74]), .Z(wk_share1[10]) );
  XOR2_X1 KeySchadule1_U1 ( .A(Key1[0]), .B(Key1[64]), .Z(wk_share1[0]) );
  XOR2_X1 KeySchadule2_U64 ( .A(Key2[73]), .B(Key2[9]), .Z(wk_share2[9]) );
  XOR2_X1 KeySchadule2_U63 ( .A(Key2[72]), .B(Key2[8]), .Z(wk_share2[8]) );
  XOR2_X1 KeySchadule2_U62 ( .A(Key2[71]), .B(Key2[7]), .Z(wk_share2[7]) );
  XOR2_X1 KeySchadule2_U61 ( .A(Key2[6]), .B(Key2[70]), .Z(wk_share2[6]) );
  XOR2_X1 KeySchadule2_U60 ( .A(Key2[127]), .B(Key2[63]), .Z(wk_share2[63]) );
  XOR2_X1 KeySchadule2_U59 ( .A(Key2[126]), .B(Key2[62]), .Z(wk_share2[62]) );
  XOR2_X1 KeySchadule2_U58 ( .A(Key2[125]), .B(Key2[61]), .Z(wk_share2[61]) );
  XOR2_X1 KeySchadule2_U57 ( .A(Key2[124]), .B(Key2[60]), .Z(wk_share2[60]) );
  XOR2_X1 KeySchadule2_U56 ( .A(Key2[5]), .B(Key2[69]), .Z(wk_share2[5]) );
  XOR2_X1 KeySchadule2_U55 ( .A(Key2[123]), .B(Key2[59]), .Z(wk_share2[59]) );
  XOR2_X1 KeySchadule2_U54 ( .A(Key2[122]), .B(Key2[58]), .Z(wk_share2[58]) );
  XOR2_X1 KeySchadule2_U53 ( .A(Key2[121]), .B(Key2[57]), .Z(wk_share2[57]) );
  XOR2_X1 KeySchadule2_U52 ( .A(Key2[120]), .B(Key2[56]), .Z(wk_share2[56]) );
  XOR2_X1 KeySchadule2_U51 ( .A(Key2[119]), .B(Key2[55]), .Z(wk_share2[55]) );
  XOR2_X1 KeySchadule2_U50 ( .A(Key2[118]), .B(Key2[54]), .Z(wk_share2[54]) );
  XOR2_X1 KeySchadule2_U49 ( .A(Key2[117]), .B(Key2[53]), .Z(wk_share2[53]) );
  XOR2_X1 KeySchadule2_U48 ( .A(Key2[116]), .B(Key2[52]), .Z(wk_share2[52]) );
  XOR2_X1 KeySchadule2_U47 ( .A(Key2[115]), .B(Key2[51]), .Z(wk_share2[51]) );
  XOR2_X1 KeySchadule2_U46 ( .A(Key2[114]), .B(Key2[50]), .Z(wk_share2[50]) );
  XOR2_X1 KeySchadule2_U45 ( .A(Key2[4]), .B(Key2[68]), .Z(wk_share2[4]) );
  XOR2_X1 KeySchadule2_U44 ( .A(Key2[113]), .B(Key2[49]), .Z(wk_share2[49]) );
  XOR2_X1 KeySchadule2_U43 ( .A(Key2[112]), .B(Key2[48]), .Z(wk_share2[48]) );
  XOR2_X1 KeySchadule2_U42 ( .A(Key2[111]), .B(Key2[47]), .Z(wk_share2[47]) );
  XOR2_X1 KeySchadule2_U41 ( .A(Key2[110]), .B(Key2[46]), .Z(wk_share2[46]) );
  XOR2_X1 KeySchadule2_U40 ( .A(Key2[109]), .B(Key2[45]), .Z(wk_share2[45]) );
  XOR2_X1 KeySchadule2_U39 ( .A(Key2[108]), .B(Key2[44]), .Z(wk_share2[44]) );
  XOR2_X1 KeySchadule2_U38 ( .A(Key2[107]), .B(Key2[43]), .Z(wk_share2[43]) );
  XOR2_X1 KeySchadule2_U37 ( .A(Key2[106]), .B(Key2[42]), .Z(wk_share2[42]) );
  XOR2_X1 KeySchadule2_U36 ( .A(Key2[105]), .B(Key2[41]), .Z(wk_share2[41]) );
  XOR2_X1 KeySchadule2_U35 ( .A(Key2[104]), .B(Key2[40]), .Z(wk_share2[40]) );
  XOR2_X1 KeySchadule2_U34 ( .A(Key2[3]), .B(Key2[67]), .Z(wk_share2[3]) );
  XOR2_X1 KeySchadule2_U33 ( .A(Key2[103]), .B(Key2[39]), .Z(wk_share2[39]) );
  XOR2_X1 KeySchadule2_U32 ( .A(Key2[102]), .B(Key2[38]), .Z(wk_share2[38]) );
  XOR2_X1 KeySchadule2_U31 ( .A(Key2[101]), .B(Key2[37]), .Z(wk_share2[37]) );
  XOR2_X1 KeySchadule2_U30 ( .A(Key2[100]), .B(Key2[36]), .Z(wk_share2[36]) );
  XOR2_X1 KeySchadule2_U29 ( .A(Key2[35]), .B(Key2[99]), .Z(wk_share2[35]) );
  XOR2_X1 KeySchadule2_U28 ( .A(Key2[34]), .B(Key2[98]), .Z(wk_share2[34]) );
  XOR2_X1 KeySchadule2_U27 ( .A(Key2[33]), .B(Key2[97]), .Z(wk_share2[33]) );
  XOR2_X1 KeySchadule2_U26 ( .A(Key2[32]), .B(Key2[96]), .Z(wk_share2[32]) );
  XOR2_X1 KeySchadule2_U25 ( .A(Key2[31]), .B(Key2[95]), .Z(wk_share2[31]) );
  XOR2_X1 KeySchadule2_U24 ( .A(Key2[30]), .B(Key2[94]), .Z(wk_share2[30]) );
  XOR2_X1 KeySchadule2_U23 ( .A(Key2[2]), .B(Key2[66]), .Z(wk_share2[2]) );
  XOR2_X1 KeySchadule2_U22 ( .A(Key2[29]), .B(Key2[93]), .Z(wk_share2[29]) );
  XOR2_X1 KeySchadule2_U21 ( .A(Key2[28]), .B(Key2[92]), .Z(wk_share2[28]) );
  XOR2_X1 KeySchadule2_U20 ( .A(Key2[27]), .B(Key2[91]), .Z(wk_share2[27]) );
  XOR2_X1 KeySchadule2_U19 ( .A(Key2[26]), .B(Key2[90]), .Z(wk_share2[26]) );
  XOR2_X1 KeySchadule2_U18 ( .A(Key2[25]), .B(Key2[89]), .Z(wk_share2[25]) );
  XOR2_X1 KeySchadule2_U17 ( .A(Key2[24]), .B(Key2[88]), .Z(wk_share2[24]) );
  XOR2_X1 KeySchadule2_U16 ( .A(Key2[23]), .B(Key2[87]), .Z(wk_share2[23]) );
  XOR2_X1 KeySchadule2_U15 ( .A(Key2[22]), .B(Key2[86]), .Z(wk_share2[22]) );
  XOR2_X1 KeySchadule2_U14 ( .A(Key2[21]), .B(Key2[85]), .Z(wk_share2[21]) );
  XOR2_X1 KeySchadule2_U13 ( .A(Key2[20]), .B(Key2[84]), .Z(wk_share2[20]) );
  XOR2_X1 KeySchadule2_U12 ( .A(Key2[1]), .B(Key2[65]), .Z(wk_share2[1]) );
  XOR2_X1 KeySchadule2_U11 ( .A(Key2[19]), .B(Key2[83]), .Z(wk_share2[19]) );
  XOR2_X1 KeySchadule2_U10 ( .A(Key2[18]), .B(Key2[82]), .Z(wk_share2[18]) );
  XOR2_X1 KeySchadule2_U9 ( .A(Key2[17]), .B(Key2[81]), .Z(wk_share2[17]) );
  XOR2_X1 KeySchadule2_U8 ( .A(Key2[16]), .B(Key2[80]), .Z(wk_share2[16]) );
  XOR2_X1 KeySchadule2_U7 ( .A(Key2[15]), .B(Key2[79]), .Z(wk_share2[15]) );
  XOR2_X1 KeySchadule2_U6 ( .A(Key2[14]), .B(Key2[78]), .Z(wk_share2[14]) );
  XOR2_X1 KeySchadule2_U5 ( .A(Key2[13]), .B(Key2[77]), .Z(wk_share2[13]) );
  XOR2_X1 KeySchadule2_U4 ( .A(Key2[12]), .B(Key2[76]), .Z(wk_share2[12]) );
  XOR2_X1 KeySchadule2_U3 ( .A(Key2[11]), .B(Key2[75]), .Z(wk_share2[11]) );
  XOR2_X1 KeySchadule2_U2 ( .A(Key2[10]), .B(Key2[74]), .Z(wk_share2[10]) );
  XOR2_X1 KeySchadule2_U1 ( .A(Key2[0]), .B(Key2[64]), .Z(wk_share2[0]) );
  XOR2_X1 KeySchadule3_U64 ( .A(Key3[73]), .B(Key3[9]), .Z(wk_share3[9]) );
  XOR2_X1 KeySchadule3_U63 ( .A(Key3[72]), .B(Key3[8]), .Z(wk_share3[8]) );
  XOR2_X1 KeySchadule3_U62 ( .A(Key3[71]), .B(Key3[7]), .Z(wk_share3[7]) );
  XOR2_X1 KeySchadule3_U61 ( .A(Key3[6]), .B(Key3[70]), .Z(wk_share3[6]) );
  XOR2_X1 KeySchadule3_U60 ( .A(Key3[127]), .B(Key3[63]), .Z(wk_share3[63]) );
  XOR2_X1 KeySchadule3_U59 ( .A(Key3[126]), .B(Key3[62]), .Z(wk_share3[62]) );
  XOR2_X1 KeySchadule3_U58 ( .A(Key3[125]), .B(Key3[61]), .Z(wk_share3[61]) );
  XOR2_X1 KeySchadule3_U57 ( .A(Key3[124]), .B(Key3[60]), .Z(wk_share3[60]) );
  XOR2_X1 KeySchadule3_U56 ( .A(Key3[5]), .B(Key3[69]), .Z(wk_share3[5]) );
  XOR2_X1 KeySchadule3_U55 ( .A(Key3[123]), .B(Key3[59]), .Z(wk_share3[59]) );
  XOR2_X1 KeySchadule3_U54 ( .A(Key3[122]), .B(Key3[58]), .Z(wk_share3[58]) );
  XOR2_X1 KeySchadule3_U53 ( .A(Key3[121]), .B(Key3[57]), .Z(wk_share3[57]) );
  XOR2_X1 KeySchadule3_U52 ( .A(Key3[120]), .B(Key3[56]), .Z(wk_share3[56]) );
  XOR2_X1 KeySchadule3_U51 ( .A(Key3[119]), .B(Key3[55]), .Z(wk_share3[55]) );
  XOR2_X1 KeySchadule3_U50 ( .A(Key3[118]), .B(Key3[54]), .Z(wk_share3[54]) );
  XOR2_X1 KeySchadule3_U49 ( .A(Key3[117]), .B(Key3[53]), .Z(wk_share3[53]) );
  XOR2_X1 KeySchadule3_U48 ( .A(Key3[116]), .B(Key3[52]), .Z(wk_share3[52]) );
  XOR2_X1 KeySchadule3_U47 ( .A(Key3[115]), .B(Key3[51]), .Z(wk_share3[51]) );
  XOR2_X1 KeySchadule3_U46 ( .A(Key3[114]), .B(Key3[50]), .Z(wk_share3[50]) );
  XOR2_X1 KeySchadule3_U45 ( .A(Key3[4]), .B(Key3[68]), .Z(wk_share3[4]) );
  XOR2_X1 KeySchadule3_U44 ( .A(Key3[113]), .B(Key3[49]), .Z(wk_share3[49]) );
  XOR2_X1 KeySchadule3_U43 ( .A(Key3[112]), .B(Key3[48]), .Z(wk_share3[48]) );
  XOR2_X1 KeySchadule3_U42 ( .A(Key3[111]), .B(Key3[47]), .Z(wk_share3[47]) );
  XOR2_X1 KeySchadule3_U41 ( .A(Key3[110]), .B(Key3[46]), .Z(wk_share3[46]) );
  XOR2_X1 KeySchadule3_U40 ( .A(Key3[109]), .B(Key3[45]), .Z(wk_share3[45]) );
  XOR2_X1 KeySchadule3_U39 ( .A(Key3[108]), .B(Key3[44]), .Z(wk_share3[44]) );
  XOR2_X1 KeySchadule3_U38 ( .A(Key3[107]), .B(Key3[43]), .Z(wk_share3[43]) );
  XOR2_X1 KeySchadule3_U37 ( .A(Key3[106]), .B(Key3[42]), .Z(wk_share3[42]) );
  XOR2_X1 KeySchadule3_U36 ( .A(Key3[105]), .B(Key3[41]), .Z(wk_share3[41]) );
  XOR2_X1 KeySchadule3_U35 ( .A(Key3[104]), .B(Key3[40]), .Z(wk_share3[40]) );
  XOR2_X1 KeySchadule3_U34 ( .A(Key3[3]), .B(Key3[67]), .Z(wk_share3[3]) );
  XOR2_X1 KeySchadule3_U33 ( .A(Key3[103]), .B(Key3[39]), .Z(wk_share3[39]) );
  XOR2_X1 KeySchadule3_U32 ( .A(Key3[102]), .B(Key3[38]), .Z(wk_share3[38]) );
  XOR2_X1 KeySchadule3_U31 ( .A(Key3[101]), .B(Key3[37]), .Z(wk_share3[37]) );
  XOR2_X1 KeySchadule3_U30 ( .A(Key3[100]), .B(Key3[36]), .Z(wk_share3[36]) );
  XOR2_X1 KeySchadule3_U29 ( .A(Key3[35]), .B(Key3[99]), .Z(wk_share3[35]) );
  XOR2_X1 KeySchadule3_U28 ( .A(Key3[34]), .B(Key3[98]), .Z(wk_share3[34]) );
  XOR2_X1 KeySchadule3_U27 ( .A(Key3[33]), .B(Key3[97]), .Z(wk_share3[33]) );
  XOR2_X1 KeySchadule3_U26 ( .A(Key3[32]), .B(Key3[96]), .Z(wk_share3[32]) );
  XOR2_X1 KeySchadule3_U25 ( .A(Key3[31]), .B(Key3[95]), .Z(wk_share3[31]) );
  XOR2_X1 KeySchadule3_U24 ( .A(Key3[30]), .B(Key3[94]), .Z(wk_share3[30]) );
  XOR2_X1 KeySchadule3_U23 ( .A(Key3[2]), .B(Key3[66]), .Z(wk_share3[2]) );
  XOR2_X1 KeySchadule3_U22 ( .A(Key3[29]), .B(Key3[93]), .Z(wk_share3[29]) );
  XOR2_X1 KeySchadule3_U21 ( .A(Key3[28]), .B(Key3[92]), .Z(wk_share3[28]) );
  XOR2_X1 KeySchadule3_U20 ( .A(Key3[27]), .B(Key3[91]), .Z(wk_share3[27]) );
  XOR2_X1 KeySchadule3_U19 ( .A(Key3[26]), .B(Key3[90]), .Z(wk_share3[26]) );
  XOR2_X1 KeySchadule3_U18 ( .A(Key3[25]), .B(Key3[89]), .Z(wk_share3[25]) );
  XOR2_X1 KeySchadule3_U17 ( .A(Key3[24]), .B(Key3[88]), .Z(wk_share3[24]) );
  XOR2_X1 KeySchadule3_U16 ( .A(Key3[23]), .B(Key3[87]), .Z(wk_share3[23]) );
  XOR2_X1 KeySchadule3_U15 ( .A(Key3[22]), .B(Key3[86]), .Z(wk_share3[22]) );
  XOR2_X1 KeySchadule3_U14 ( .A(Key3[21]), .B(Key3[85]), .Z(wk_share3[21]) );
  XOR2_X1 KeySchadule3_U13 ( .A(Key3[20]), .B(Key3[84]), .Z(wk_share3[20]) );
  XOR2_X1 KeySchadule3_U12 ( .A(Key3[1]), .B(Key3[65]), .Z(wk_share3[1]) );
  XOR2_X1 KeySchadule3_U11 ( .A(Key3[19]), .B(Key3[83]), .Z(wk_share3[19]) );
  XOR2_X1 KeySchadule3_U10 ( .A(Key3[18]), .B(Key3[82]), .Z(wk_share3[18]) );
  XOR2_X1 KeySchadule3_U9 ( .A(Key3[17]), .B(Key3[81]), .Z(wk_share3[17]) );
  XOR2_X1 KeySchadule3_U8 ( .A(Key3[16]), .B(Key3[80]), .Z(wk_share3[16]) );
  XOR2_X1 KeySchadule3_U7 ( .A(Key3[15]), .B(Key3[79]), .Z(wk_share3[15]) );
  XOR2_X1 KeySchadule3_U6 ( .A(Key3[14]), .B(Key3[78]), .Z(wk_share3[14]) );
  XOR2_X1 KeySchadule3_U5 ( .A(Key3[13]), .B(Key3[77]), .Z(wk_share3[13]) );
  XOR2_X1 KeySchadule3_U4 ( .A(Key3[12]), .B(Key3[76]), .Z(wk_share3[12]) );
  XOR2_X1 KeySchadule3_U3 ( .A(Key3[11]), .B(Key3[75]), .Z(wk_share3[11]) );
  XOR2_X1 KeySchadule3_U2 ( .A(Key3[10]), .B(Key3[74]), .Z(wk_share3[10]) );
  XOR2_X1 KeySchadule3_U1 ( .A(Key3[0]), .B(Key3[64]), .Z(wk_share3[0]) );
  AND4_X1 controller_U1 ( .A1(round_Signal[2]), .A2(round_Signal[3]), .A3(
        round_Signal[0]), .A4(round_Signal[1]), .ZN(done) );
  AOI21_X1 controller_roundCounter_U20 ( .B1(controller_roundCounter_q_0_), 
        .B2(EN), .A(reset), .ZN(controller_roundCounter_n15) );
  AOI21_X1 controller_roundCounter_U19 ( .B1(controller_roundCounter_n34), 
        .B2(controller_roundCounter_n22), .A(reset), .ZN(
        controller_roundCounter_n14) );
  AOI21_X1 controller_roundCounter_U18 ( .B1(EN), .B2(
        controller_roundCounter_n33), .A(reset), .ZN(
        controller_roundCounter_n13) );
  OAI21_X1 controller_roundCounter_U17 ( .B1(controller_roundCounter_q_0_), 
        .B2(controller_roundCounter_q_1_), .A(controller_roundCounter_n32), 
        .ZN(controller_roundCounter_n33) );
  AOI21_X1 controller_roundCounter_U16 ( .B1(EN), .B2(
        controller_roundCounter_n31), .A(reset), .ZN(
        controller_roundCounter_n12) );
  OAI21_X1 controller_roundCounter_U15 ( .B1(controller_roundCounter_n30), 
        .B2(round_Signal[0]), .A(controller_roundCounter_n29), .ZN(
        controller_roundCounter_n31) );
  AOI21_X1 controller_roundCounter_U14 ( .B1(EN), .B2(
        controller_roundCounter_n28), .A(reset), .ZN(
        controller_roundCounter_n11) );
  OAI21_X1 controller_roundCounter_U13 ( .B1(controller_roundCounter_n27), 
        .B2(round_Signal[1]), .A(controller_roundCounter_n26), .ZN(
        controller_roundCounter_n28) );
  AOI211_X1 controller_roundCounter_U12 ( .C1(controller_roundCounter_n23), 
        .C2(controller_roundCounter_n26), .A(reset), .B(
        controller_roundCounter_n25), .ZN(controller_roundCounter_n10) );
  NOR2_X1 controller_roundCounter_U11 ( .A1(round_Signal[3]), .A2(
        controller_roundCounter_n34), .ZN(controller_roundCounter_n25) );
  INV_X1 controller_roundCounter_U10 ( .A(controller_roundCounter_n24), .ZN(
        controller_roundCounter_n34) );
  NAND2_X1 controller_roundCounter_U9 ( .A1(controller_roundCounter_n24), .A2(
        round_Signal[3]), .ZN(EN) );
  NOR2_X1 controller_roundCounter_U8 ( .A1(controller_roundCounter_n23), .A2(
        controller_roundCounter_n26), .ZN(controller_roundCounter_n24) );
  NAND2_X1 controller_roundCounter_U7 ( .A1(controller_roundCounter_n27), .A2(
        round_Signal[1]), .ZN(controller_roundCounter_n26) );
  INV_X1 controller_roundCounter_U6 ( .A(controller_roundCounter_n29), .ZN(
        controller_roundCounter_n27) );
  NAND2_X1 controller_roundCounter_U5 ( .A1(controller_roundCounter_n30), .A2(
        round_Signal[0]), .ZN(controller_roundCounter_n29) );
  INV_X1 controller_roundCounter_U4 ( .A(controller_roundCounter_n32), .ZN(
        controller_roundCounter_n30) );
  NAND2_X1 controller_roundCounter_U3 ( .A1(controller_roundCounter_q_0_), 
        .A2(controller_roundCounter_q_1_), .ZN(controller_roundCounter_n32) );
  DFF_X1 controller_roundCounter_count_reg_4_ ( .D(controller_roundCounter_n10), .CK(clk), .Q(round_Signal[2]), .QN(controller_roundCounter_n23) );
  DFF_X1 controller_roundCounter_count_reg_3_ ( .D(controller_roundCounter_n11), .CK(clk), .Q(round_Signal[1]), .QN() );
  DFF_X1 controller_roundCounter_count_reg_2_ ( .D(controller_roundCounter_n12), .CK(clk), .Q(round_Signal[0]), .QN() );
  DFF_X1 controller_roundCounter_count_reg_1_ ( .D(controller_roundCounter_n13), .CK(clk), .Q(controller_roundCounter_q_1_), .QN() );
  DFF_X1 controller_roundCounter_count_reg_5_ ( .D(controller_roundCounter_n14), .CK(clk), .Q(round_Signal[3]), .QN(controller_roundCounter_n22) );
  DFF_X1 controller_roundCounter_count_reg_0_ ( .D(controller_roundCounter_n15), .CK(clk), .Q(controller_roundCounter_q_0_), .QN() );
  XOR2_X1 Midori_U384 ( .A(wk_share3[9]), .B(Midori_rounds_SR_Result3[9]), .Z(
        output3[9]) );
  XOR2_X1 Midori_U383 ( .A(wk_share3[8]), .B(Midori_rounds_SR_Result3[8]), .Z(
        output3[8]) );
  XOR2_X1 Midori_U382 ( .A(wk_share3[7]), .B(Midori_rounds_SR_Result3[47]), 
        .Z(output3[7]) );
  XOR2_X1 Midori_U381 ( .A(wk_share3[6]), .B(Midori_rounds_SR_Result3[46]), 
        .Z(output3[6]) );
  XOR2_X1 Midori_U380 ( .A(wk_share3[63]), .B(Midori_rounds_SR_Result3[63]), 
        .Z(output3[63]) );
  XOR2_X1 Midori_U379 ( .A(wk_share3[62]), .B(Midori_rounds_SR_Result3[62]), 
        .Z(output3[62]) );
  XOR2_X1 Midori_U378 ( .A(wk_share3[61]), .B(Midori_rounds_SR_Result3[61]), 
        .Z(output3[61]) );
  XOR2_X1 Midori_U377 ( .A(wk_share3[60]), .B(Midori_rounds_SR_Result3[60]), 
        .Z(output3[60]) );
  XOR2_X1 Midori_U376 ( .A(wk_share3[5]), .B(Midori_rounds_SR_Result3[45]), 
        .Z(output3[5]) );
  XOR2_X1 Midori_U375 ( .A(wk_share3[59]), .B(Midori_rounds_SR_Result3[35]), 
        .Z(output3[59]) );
  XOR2_X1 Midori_U374 ( .A(wk_share3[58]), .B(Midori_rounds_SR_Result3[34]), 
        .Z(output3[58]) );
  XOR2_X1 Midori_U373 ( .A(wk_share3[57]), .B(Midori_rounds_SR_Result3[33]), 
        .Z(output3[57]) );
  XOR2_X1 Midori_U372 ( .A(wk_share3[56]), .B(Midori_rounds_SR_Result3[32]), 
        .Z(output3[56]) );
  XOR2_X1 Midori_U371 ( .A(wk_share3[55]), .B(Midori_rounds_SR_Result3[7]), 
        .Z(output3[55]) );
  XOR2_X1 Midori_U370 ( .A(wk_share3[54]), .B(Midori_rounds_SR_Result3[6]), 
        .Z(output3[54]) );
  XOR2_X1 Midori_U369 ( .A(wk_share3[53]), .B(Midori_rounds_SR_Result3[5]), 
        .Z(output3[53]) );
  XOR2_X1 Midori_U368 ( .A(wk_share3[52]), .B(Midori_rounds_SR_Result3[4]), 
        .Z(output3[52]) );
  XOR2_X1 Midori_U367 ( .A(wk_share3[51]), .B(Midori_rounds_SR_Result3[27]), 
        .Z(output3[51]) );
  XOR2_X1 Midori_U366 ( .A(wk_share3[50]), .B(Midori_rounds_SR_Result3[26]), 
        .Z(output3[50]) );
  XOR2_X1 Midori_U365 ( .A(wk_share3[4]), .B(Midori_rounds_SR_Result3[44]), 
        .Z(output3[4]) );
  XOR2_X1 Midori_U364 ( .A(wk_share3[49]), .B(Midori_rounds_SR_Result3[25]), 
        .Z(output3[49]) );
  XOR2_X1 Midori_U363 ( .A(wk_share3[48]), .B(Midori_rounds_SR_Result3[24]), 
        .Z(output3[48]) );
  XOR2_X1 Midori_U362 ( .A(wk_share3[47]), .B(Midori_rounds_SR_Result3[43]), 
        .Z(output3[47]) );
  XOR2_X1 Midori_U361 ( .A(wk_share3[46]), .B(Midori_rounds_SR_Result3[42]), 
        .Z(output3[46]) );
  XOR2_X1 Midori_U360 ( .A(wk_share3[45]), .B(Midori_rounds_SR_Result3[41]), 
        .Z(output3[45]) );
  XOR2_X1 Midori_U359 ( .A(wk_share3[44]), .B(Midori_rounds_SR_Result3[40]), 
        .Z(output3[44]) );
  XOR2_X1 Midori_U358 ( .A(wk_share3[43]), .B(Midori_rounds_SR_Result3[55]), 
        .Z(output3[43]) );
  XOR2_X1 Midori_U357 ( .A(wk_share3[42]), .B(Midori_rounds_SR_Result3[54]), 
        .Z(output3[42]) );
  XOR2_X1 Midori_U356 ( .A(wk_share3[41]), .B(Midori_rounds_SR_Result3[53]), 
        .Z(output3[41]) );
  XOR2_X1 Midori_U355 ( .A(wk_share3[40]), .B(Midori_rounds_SR_Result3[52]), 
        .Z(output3[40]) );
  XOR2_X1 Midori_U354 ( .A(wk_share3[3]), .B(Midori_rounds_SR_Result3[51]), 
        .Z(output3[3]) );
  XOR2_X1 Midori_U353 ( .A(wk_share3[39]), .B(Midori_rounds_SR_Result3[19]), 
        .Z(output3[39]) );
  XOR2_X1 Midori_U352 ( .A(wk_share3[38]), .B(Midori_rounds_SR_Result3[18]), 
        .Z(output3[38]) );
  XOR2_X1 Midori_U351 ( .A(wk_share3[37]), .B(Midori_rounds_SR_Result3[17]), 
        .Z(output3[37]) );
  XOR2_X1 Midori_U350 ( .A(wk_share3[36]), .B(Midori_rounds_SR_Result3[16]), 
        .Z(output3[36]) );
  XOR2_X1 Midori_U349 ( .A(wk_share3[35]), .B(Midori_rounds_SR_Result3[15]), 
        .Z(output3[35]) );
  XOR2_X1 Midori_U348 ( .A(wk_share3[34]), .B(Midori_rounds_SR_Result3[14]), 
        .Z(output3[34]) );
  XOR2_X1 Midori_U347 ( .A(wk_share3[33]), .B(Midori_rounds_SR_Result3[13]), 
        .Z(output3[33]) );
  XOR2_X1 Midori_U346 ( .A(wk_share3[32]), .B(Midori_rounds_SR_Result3[12]), 
        .Z(output3[32]) );
  XOR2_X1 Midori_U345 ( .A(wk_share3[31]), .B(Midori_rounds_SR_Result3[3]), 
        .Z(output3[31]) );
  XOR2_X1 Midori_U344 ( .A(wk_share3[30]), .B(Midori_rounds_SR_Result3[2]), 
        .Z(output3[30]) );
  XOR2_X1 Midori_U343 ( .A(wk_share3[2]), .B(Midori_rounds_SR_Result3[50]), 
        .Z(output3[2]) );
  XOR2_X1 Midori_U342 ( .A(wk_share3[29]), .B(Midori_rounds_SR_Result3[1]), 
        .Z(output3[29]) );
  XOR2_X1 Midori_U341 ( .A(wk_share3[28]), .B(Midori_rounds_SR_Result3[0]), 
        .Z(output3[28]) );
  XOR2_X1 Midori_U340 ( .A(wk_share3[27]), .B(Midori_rounds_SR_Result3[31]), 
        .Z(output3[27]) );
  XOR2_X1 Midori_U339 ( .A(wk_share3[26]), .B(Midori_rounds_SR_Result3[30]), 
        .Z(output3[26]) );
  XOR2_X1 Midori_U338 ( .A(wk_share3[25]), .B(Midori_rounds_SR_Result3[29]), 
        .Z(output3[25]) );
  XOR2_X1 Midori_U337 ( .A(wk_share3[24]), .B(Midori_rounds_SR_Result3[28]), 
        .Z(output3[24]) );
  XOR2_X1 Midori_U336 ( .A(wk_share3[23]), .B(Midori_rounds_SR_Result3[59]), 
        .Z(output3[23]) );
  XOR2_X1 Midori_U335 ( .A(wk_share3[22]), .B(Midori_rounds_SR_Result3[58]), 
        .Z(output3[22]) );
  XOR2_X1 Midori_U334 ( .A(wk_share3[21]), .B(Midori_rounds_SR_Result3[57]), 
        .Z(output3[21]) );
  XOR2_X1 Midori_U333 ( .A(wk_share3[20]), .B(Midori_rounds_SR_Result3[56]), 
        .Z(output3[20]) );
  XOR2_X1 Midori_U332 ( .A(wk_share3[1]), .B(Midori_rounds_SR_Result3[49]), 
        .Z(output3[1]) );
  XOR2_X1 Midori_U331 ( .A(wk_share3[19]), .B(Midori_rounds_SR_Result3[39]), 
        .Z(output3[19]) );
  XOR2_X1 Midori_U330 ( .A(wk_share3[18]), .B(Midori_rounds_SR_Result3[38]), 
        .Z(output3[18]) );
  XOR2_X1 Midori_U329 ( .A(wk_share3[17]), .B(Midori_rounds_SR_Result3[37]), 
        .Z(output3[17]) );
  XOR2_X1 Midori_U328 ( .A(wk_share3[16]), .B(Midori_rounds_SR_Result3[36]), 
        .Z(output3[16]) );
  XOR2_X1 Midori_U327 ( .A(wk_share3[15]), .B(Midori_rounds_SR_Result3[23]), 
        .Z(output3[15]) );
  XOR2_X1 Midori_U326 ( .A(wk_share3[14]), .B(Midori_rounds_SR_Result3[22]), 
        .Z(output3[14]) );
  XOR2_X1 Midori_U325 ( .A(wk_share3[13]), .B(Midori_rounds_SR_Result3[21]), 
        .Z(output3[13]) );
  XOR2_X1 Midori_U324 ( .A(wk_share3[12]), .B(Midori_rounds_SR_Result3[20]), 
        .Z(output3[12]) );
  XOR2_X1 Midori_U323 ( .A(wk_share3[11]), .B(Midori_rounds_SR_Result3[11]), 
        .Z(output3[11]) );
  XOR2_X1 Midori_U322 ( .A(wk_share3[10]), .B(Midori_rounds_SR_Result3[10]), 
        .Z(output3[10]) );
  XOR2_X1 Midori_U321 ( .A(wk_share3[0]), .B(Midori_rounds_SR_Result3[48]), 
        .Z(output3[0]) );
  XOR2_X1 Midori_U320 ( .A(wk_share2[9]), .B(Midori_rounds_SR_Result2[9]), .Z(
        output2[9]) );
  XOR2_X1 Midori_U319 ( .A(wk_share2[8]), .B(Midori_rounds_SR_Result2[8]), .Z(
        output2[8]) );
  XOR2_X1 Midori_U318 ( .A(wk_share2[7]), .B(Midori_rounds_SR_Result2[47]), 
        .Z(output2[7]) );
  XOR2_X1 Midori_U317 ( .A(wk_share2[6]), .B(Midori_rounds_SR_Result2[46]), 
        .Z(output2[6]) );
  XOR2_X1 Midori_U316 ( .A(wk_share2[63]), .B(Midori_rounds_SR_Result2[63]), 
        .Z(output2[63]) );
  XOR2_X1 Midori_U315 ( .A(wk_share2[62]), .B(Midori_rounds_SR_Result2[62]), 
        .Z(output2[62]) );
  XOR2_X1 Midori_U314 ( .A(wk_share2[61]), .B(Midori_rounds_SR_Result2[61]), 
        .Z(output2[61]) );
  XOR2_X1 Midori_U313 ( .A(wk_share2[60]), .B(Midori_rounds_SR_Result2[60]), 
        .Z(output2[60]) );
  XOR2_X1 Midori_U312 ( .A(wk_share2[5]), .B(Midori_rounds_SR_Result2[45]), 
        .Z(output2[5]) );
  XOR2_X1 Midori_U311 ( .A(wk_share2[59]), .B(Midori_rounds_SR_Result2[35]), 
        .Z(output2[59]) );
  XOR2_X1 Midori_U310 ( .A(wk_share2[58]), .B(Midori_rounds_SR_Result2[34]), 
        .Z(output2[58]) );
  XOR2_X1 Midori_U309 ( .A(wk_share2[57]), .B(Midori_rounds_SR_Result2[33]), 
        .Z(output2[57]) );
  XOR2_X1 Midori_U308 ( .A(wk_share2[56]), .B(Midori_rounds_SR_Result2[32]), 
        .Z(output2[56]) );
  XOR2_X1 Midori_U307 ( .A(wk_share2[55]), .B(Midori_rounds_SR_Result2[7]), 
        .Z(output2[55]) );
  XOR2_X1 Midori_U306 ( .A(wk_share2[54]), .B(Midori_rounds_SR_Result2[6]), 
        .Z(output2[54]) );
  XOR2_X1 Midori_U305 ( .A(wk_share2[53]), .B(Midori_rounds_SR_Result2[5]), 
        .Z(output2[53]) );
  XOR2_X1 Midori_U304 ( .A(wk_share2[52]), .B(Midori_rounds_SR_Result2[4]), 
        .Z(output2[52]) );
  XOR2_X1 Midori_U303 ( .A(wk_share2[51]), .B(Midori_rounds_SR_Result2[27]), 
        .Z(output2[51]) );
  XOR2_X1 Midori_U302 ( .A(wk_share2[50]), .B(Midori_rounds_SR_Result2[26]), 
        .Z(output2[50]) );
  XOR2_X1 Midori_U301 ( .A(wk_share2[4]), .B(Midori_rounds_SR_Result2[44]), 
        .Z(output2[4]) );
  XOR2_X1 Midori_U300 ( .A(wk_share2[49]), .B(Midori_rounds_SR_Result2[25]), 
        .Z(output2[49]) );
  XOR2_X1 Midori_U299 ( .A(wk_share2[48]), .B(Midori_rounds_SR_Result2[24]), 
        .Z(output2[48]) );
  XOR2_X1 Midori_U298 ( .A(wk_share2[47]), .B(Midori_rounds_SR_Result2[43]), 
        .Z(output2[47]) );
  XOR2_X1 Midori_U297 ( .A(wk_share2[46]), .B(Midori_rounds_SR_Result2[42]), 
        .Z(output2[46]) );
  XOR2_X1 Midori_U296 ( .A(wk_share2[45]), .B(Midori_rounds_SR_Result2[41]), 
        .Z(output2[45]) );
  XOR2_X1 Midori_U295 ( .A(wk_share2[44]), .B(Midori_rounds_SR_Result2[40]), 
        .Z(output2[44]) );
  XOR2_X1 Midori_U294 ( .A(wk_share2[43]), .B(Midori_rounds_SR_Result2[55]), 
        .Z(output2[43]) );
  XOR2_X1 Midori_U293 ( .A(wk_share2[42]), .B(Midori_rounds_SR_Result2[54]), 
        .Z(output2[42]) );
  XOR2_X1 Midori_U292 ( .A(wk_share2[41]), .B(Midori_rounds_SR_Result2[53]), 
        .Z(output2[41]) );
  XOR2_X1 Midori_U291 ( .A(wk_share2[40]), .B(Midori_rounds_SR_Result2[52]), 
        .Z(output2[40]) );
  XOR2_X1 Midori_U290 ( .A(wk_share2[3]), .B(Midori_rounds_SR_Result2[51]), 
        .Z(output2[3]) );
  XOR2_X1 Midori_U289 ( .A(wk_share2[39]), .B(Midori_rounds_SR_Result2[19]), 
        .Z(output2[39]) );
  XOR2_X1 Midori_U288 ( .A(wk_share2[38]), .B(Midori_rounds_SR_Result2[18]), 
        .Z(output2[38]) );
  XOR2_X1 Midori_U287 ( .A(wk_share2[37]), .B(Midori_rounds_SR_Result2[17]), 
        .Z(output2[37]) );
  XOR2_X1 Midori_U286 ( .A(wk_share2[36]), .B(Midori_rounds_SR_Result2[16]), 
        .Z(output2[36]) );
  XOR2_X1 Midori_U285 ( .A(wk_share2[35]), .B(Midori_rounds_SR_Result2[15]), 
        .Z(output2[35]) );
  XOR2_X1 Midori_U284 ( .A(wk_share2[34]), .B(Midori_rounds_SR_Result2[14]), 
        .Z(output2[34]) );
  XOR2_X1 Midori_U283 ( .A(wk_share2[33]), .B(Midori_rounds_SR_Result2[13]), 
        .Z(output2[33]) );
  XOR2_X1 Midori_U282 ( .A(wk_share2[32]), .B(Midori_rounds_SR_Result2[12]), 
        .Z(output2[32]) );
  XOR2_X1 Midori_U281 ( .A(wk_share2[31]), .B(Midori_rounds_SR_Result2[3]), 
        .Z(output2[31]) );
  XOR2_X1 Midori_U280 ( .A(wk_share2[30]), .B(Midori_rounds_SR_Result2[2]), 
        .Z(output2[30]) );
  XOR2_X1 Midori_U279 ( .A(wk_share2[2]), .B(Midori_rounds_SR_Result2[50]), 
        .Z(output2[2]) );
  XOR2_X1 Midori_U278 ( .A(wk_share2[29]), .B(Midori_rounds_SR_Result2[1]), 
        .Z(output2[29]) );
  XOR2_X1 Midori_U277 ( .A(wk_share2[28]), .B(Midori_rounds_SR_Result2[0]), 
        .Z(output2[28]) );
  XOR2_X1 Midori_U276 ( .A(wk_share2[27]), .B(Midori_rounds_SR_Result2[31]), 
        .Z(output2[27]) );
  XOR2_X1 Midori_U275 ( .A(wk_share2[26]), .B(Midori_rounds_SR_Result2[30]), 
        .Z(output2[26]) );
  XOR2_X1 Midori_U274 ( .A(wk_share2[25]), .B(Midori_rounds_SR_Result2[29]), 
        .Z(output2[25]) );
  XOR2_X1 Midori_U273 ( .A(wk_share2[24]), .B(Midori_rounds_SR_Result2[28]), 
        .Z(output2[24]) );
  XOR2_X1 Midori_U272 ( .A(wk_share2[23]), .B(Midori_rounds_SR_Result2[59]), 
        .Z(output2[23]) );
  XOR2_X1 Midori_U271 ( .A(wk_share2[22]), .B(Midori_rounds_SR_Result2[58]), 
        .Z(output2[22]) );
  XOR2_X1 Midori_U270 ( .A(wk_share2[21]), .B(Midori_rounds_SR_Result2[57]), 
        .Z(output2[21]) );
  XOR2_X1 Midori_U269 ( .A(wk_share2[20]), .B(Midori_rounds_SR_Result2[56]), 
        .Z(output2[20]) );
  XOR2_X1 Midori_U268 ( .A(wk_share2[1]), .B(Midori_rounds_SR_Result2[49]), 
        .Z(output2[1]) );
  XOR2_X1 Midori_U267 ( .A(wk_share2[19]), .B(Midori_rounds_SR_Result2[39]), 
        .Z(output2[19]) );
  XOR2_X1 Midori_U266 ( .A(wk_share2[18]), .B(Midori_rounds_SR_Result2[38]), 
        .Z(output2[18]) );
  XOR2_X1 Midori_U265 ( .A(wk_share2[17]), .B(Midori_rounds_SR_Result2[37]), 
        .Z(output2[17]) );
  XOR2_X1 Midori_U264 ( .A(wk_share2[16]), .B(Midori_rounds_SR_Result2[36]), 
        .Z(output2[16]) );
  XOR2_X1 Midori_U263 ( .A(wk_share2[15]), .B(Midori_rounds_SR_Result2[23]), 
        .Z(output2[15]) );
  XOR2_X1 Midori_U262 ( .A(wk_share2[14]), .B(Midori_rounds_SR_Result2[22]), 
        .Z(output2[14]) );
  XOR2_X1 Midori_U261 ( .A(wk_share2[13]), .B(Midori_rounds_SR_Result2[21]), 
        .Z(output2[13]) );
  XOR2_X1 Midori_U260 ( .A(wk_share2[12]), .B(Midori_rounds_SR_Result2[20]), 
        .Z(output2[12]) );
  XOR2_X1 Midori_U259 ( .A(wk_share2[11]), .B(Midori_rounds_SR_Result2[11]), 
        .Z(output2[11]) );
  XOR2_X1 Midori_U258 ( .A(wk_share2[10]), .B(Midori_rounds_SR_Result2[10]), 
        .Z(output2[10]) );
  XOR2_X1 Midori_U257 ( .A(wk_share2[0]), .B(Midori_rounds_SR_Result2[48]), 
        .Z(output2[0]) );
  XOR2_X1 Midori_U256 ( .A(wk_share1[9]), .B(Midori_rounds_SR_Result1[9]), .Z(
        output1[9]) );
  XOR2_X1 Midori_U255 ( .A(wk_share1[8]), .B(Midori_rounds_SR_Result1[8]), .Z(
        output1[8]) );
  XOR2_X1 Midori_U254 ( .A(wk_share1[7]), .B(Midori_rounds_SR_Result1[47]), 
        .Z(output1[7]) );
  XOR2_X1 Midori_U253 ( .A(wk_share1[6]), .B(Midori_rounds_SR_Result1[46]), 
        .Z(output1[6]) );
  XOR2_X1 Midori_U252 ( .A(wk_share1[63]), .B(Midori_rounds_SR_Result1[63]), 
        .Z(output1[63]) );
  XOR2_X1 Midori_U251 ( .A(wk_share1[62]), .B(Midori_rounds_SR_Result1[62]), 
        .Z(output1[62]) );
  XOR2_X1 Midori_U250 ( .A(wk_share1[61]), .B(Midori_rounds_SR_Result1[61]), 
        .Z(output1[61]) );
  XOR2_X1 Midori_U249 ( .A(wk_share1[60]), .B(Midori_rounds_SR_Result1[60]), 
        .Z(output1[60]) );
  XOR2_X1 Midori_U248 ( .A(wk_share1[5]), .B(Midori_rounds_SR_Result1[45]), 
        .Z(output1[5]) );
  XOR2_X1 Midori_U247 ( .A(wk_share1[59]), .B(Midori_rounds_SR_Result1[35]), 
        .Z(output1[59]) );
  XOR2_X1 Midori_U246 ( .A(wk_share1[58]), .B(Midori_rounds_SR_Result1[34]), 
        .Z(output1[58]) );
  XOR2_X1 Midori_U245 ( .A(wk_share1[57]), .B(Midori_rounds_SR_Result1[33]), 
        .Z(output1[57]) );
  XOR2_X1 Midori_U244 ( .A(wk_share1[56]), .B(Midori_rounds_SR_Result1[32]), 
        .Z(output1[56]) );
  XOR2_X1 Midori_U243 ( .A(wk_share1[55]), .B(Midori_rounds_SR_Result1[7]), 
        .Z(output1[55]) );
  XOR2_X1 Midori_U242 ( .A(wk_share1[54]), .B(Midori_rounds_SR_Result1[6]), 
        .Z(output1[54]) );
  XOR2_X1 Midori_U241 ( .A(wk_share1[53]), .B(Midori_rounds_SR_Result1[5]), 
        .Z(output1[53]) );
  XOR2_X1 Midori_U240 ( .A(wk_share1[52]), .B(Midori_rounds_SR_Result1[4]), 
        .Z(output1[52]) );
  XOR2_X1 Midori_U239 ( .A(wk_share1[51]), .B(Midori_rounds_SR_Result1[27]), 
        .Z(output1[51]) );
  XOR2_X1 Midori_U238 ( .A(wk_share1[50]), .B(Midori_rounds_SR_Result1[26]), 
        .Z(output1[50]) );
  XOR2_X1 Midori_U237 ( .A(wk_share1[4]), .B(Midori_rounds_SR_Result1[44]), 
        .Z(output1[4]) );
  XOR2_X1 Midori_U236 ( .A(wk_share1[49]), .B(Midori_rounds_SR_Result1[25]), 
        .Z(output1[49]) );
  XOR2_X1 Midori_U235 ( .A(wk_share1[48]), .B(Midori_rounds_SR_Result1[24]), 
        .Z(output1[48]) );
  XOR2_X1 Midori_U234 ( .A(wk_share1[47]), .B(Midori_rounds_SR_Result1[43]), 
        .Z(output1[47]) );
  XOR2_X1 Midori_U233 ( .A(wk_share1[46]), .B(Midori_rounds_SR_Result1[42]), 
        .Z(output1[46]) );
  XOR2_X1 Midori_U232 ( .A(wk_share1[45]), .B(Midori_rounds_SR_Result1[41]), 
        .Z(output1[45]) );
  XOR2_X1 Midori_U231 ( .A(wk_share1[44]), .B(Midori_rounds_SR_Result1[40]), 
        .Z(output1[44]) );
  XOR2_X1 Midori_U230 ( .A(wk_share1[43]), .B(Midori_rounds_SR_Result1[55]), 
        .Z(output1[43]) );
  XOR2_X1 Midori_U229 ( .A(wk_share1[42]), .B(Midori_rounds_SR_Result1[54]), 
        .Z(output1[42]) );
  XOR2_X1 Midori_U228 ( .A(wk_share1[41]), .B(Midori_rounds_SR_Result1[53]), 
        .Z(output1[41]) );
  XOR2_X1 Midori_U227 ( .A(wk_share1[40]), .B(Midori_rounds_SR_Result1[52]), 
        .Z(output1[40]) );
  XOR2_X1 Midori_U226 ( .A(wk_share1[3]), .B(Midori_rounds_SR_Result1[51]), 
        .Z(output1[3]) );
  XOR2_X1 Midori_U225 ( .A(wk_share1[39]), .B(Midori_rounds_SR_Result1[19]), 
        .Z(output1[39]) );
  XOR2_X1 Midori_U224 ( .A(wk_share1[38]), .B(Midori_rounds_SR_Result1[18]), 
        .Z(output1[38]) );
  XOR2_X1 Midori_U223 ( .A(wk_share1[37]), .B(Midori_rounds_SR_Result1[17]), 
        .Z(output1[37]) );
  XOR2_X1 Midori_U222 ( .A(wk_share1[36]), .B(Midori_rounds_SR_Result1[16]), 
        .Z(output1[36]) );
  XOR2_X1 Midori_U221 ( .A(wk_share1[35]), .B(Midori_rounds_SR_Result1[15]), 
        .Z(output1[35]) );
  XOR2_X1 Midori_U220 ( .A(wk_share1[34]), .B(Midori_rounds_SR_Result1[14]), 
        .Z(output1[34]) );
  XOR2_X1 Midori_U219 ( .A(wk_share1[33]), .B(Midori_rounds_SR_Result1[13]), 
        .Z(output1[33]) );
  XOR2_X1 Midori_U218 ( .A(wk_share1[32]), .B(Midori_rounds_SR_Result1[12]), 
        .Z(output1[32]) );
  XOR2_X1 Midori_U217 ( .A(wk_share1[31]), .B(Midori_rounds_SR_Result1[3]), 
        .Z(output1[31]) );
  XOR2_X1 Midori_U216 ( .A(wk_share1[30]), .B(Midori_rounds_SR_Result1[2]), 
        .Z(output1[30]) );
  XOR2_X1 Midori_U215 ( .A(wk_share1[2]), .B(Midori_rounds_SR_Result1[50]), 
        .Z(output1[2]) );
  XOR2_X1 Midori_U214 ( .A(wk_share1[29]), .B(Midori_rounds_SR_Result1[1]), 
        .Z(output1[29]) );
  XOR2_X1 Midori_U213 ( .A(wk_share1[28]), .B(Midori_rounds_SR_Result1[0]), 
        .Z(output1[28]) );
  XOR2_X1 Midori_U212 ( .A(wk_share1[27]), .B(Midori_rounds_SR_Result1[31]), 
        .Z(output1[27]) );
  XOR2_X1 Midori_U211 ( .A(wk_share1[26]), .B(Midori_rounds_SR_Result1[30]), 
        .Z(output1[26]) );
  XOR2_X1 Midori_U210 ( .A(wk_share1[25]), .B(Midori_rounds_SR_Result1[29]), 
        .Z(output1[25]) );
  XOR2_X1 Midori_U209 ( .A(wk_share1[24]), .B(Midori_rounds_SR_Result1[28]), 
        .Z(output1[24]) );
  XOR2_X1 Midori_U208 ( .A(wk_share1[23]), .B(Midori_rounds_SR_Result1[59]), 
        .Z(output1[23]) );
  XOR2_X1 Midori_U207 ( .A(wk_share1[22]), .B(Midori_rounds_SR_Result1[58]), 
        .Z(output1[22]) );
  XOR2_X1 Midori_U206 ( .A(wk_share1[21]), .B(Midori_rounds_SR_Result1[57]), 
        .Z(output1[21]) );
  XOR2_X1 Midori_U205 ( .A(wk_share1[20]), .B(Midori_rounds_SR_Result1[56]), 
        .Z(output1[20]) );
  XOR2_X1 Midori_U204 ( .A(wk_share1[1]), .B(Midori_rounds_SR_Result1[49]), 
        .Z(output1[1]) );
  XOR2_X1 Midori_U203 ( .A(wk_share1[19]), .B(Midori_rounds_SR_Result1[39]), 
        .Z(output1[19]) );
  XOR2_X1 Midori_U202 ( .A(wk_share1[18]), .B(Midori_rounds_SR_Result1[38]), 
        .Z(output1[18]) );
  XOR2_X1 Midori_U201 ( .A(wk_share1[17]), .B(Midori_rounds_SR_Result1[37]), 
        .Z(output1[17]) );
  XOR2_X1 Midori_U200 ( .A(wk_share1[16]), .B(Midori_rounds_SR_Result1[36]), 
        .Z(output1[16]) );
  XOR2_X1 Midori_U199 ( .A(wk_share1[15]), .B(Midori_rounds_SR_Result1[23]), 
        .Z(output1[15]) );
  XOR2_X1 Midori_U198 ( .A(wk_share1[14]), .B(Midori_rounds_SR_Result1[22]), 
        .Z(output1[14]) );
  XOR2_X1 Midori_U197 ( .A(wk_share1[13]), .B(Midori_rounds_SR_Result1[21]), 
        .Z(output1[13]) );
  XOR2_X1 Midori_U196 ( .A(wk_share1[12]), .B(Midori_rounds_SR_Result1[20]), 
        .Z(output1[12]) );
  XOR2_X1 Midori_U195 ( .A(wk_share1[11]), .B(Midori_rounds_SR_Result1[11]), 
        .Z(output1[11]) );
  XOR2_X1 Midori_U194 ( .A(wk_share1[10]), .B(Midori_rounds_SR_Result1[10]), 
        .Z(output1[10]) );
  XOR2_X1 Midori_U193 ( .A(wk_share1[0]), .B(Midori_rounds_SR_Result1[48]), 
        .Z(output1[0]) );
  XOR2_X1 Midori_U192 ( .A(wk_share3[9]), .B(input3[9]), .Z(
        Midori_add_Result_Start3[9]) );
  XOR2_X1 Midori_U191 ( .A(wk_share3[8]), .B(input3[8]), .Z(
        Midori_add_Result_Start3[8]) );
  XOR2_X1 Midori_U190 ( .A(wk_share3[7]), .B(input3[7]), .Z(
        Midori_add_Result_Start3[7]) );
  XOR2_X1 Midori_U189 ( .A(wk_share3[6]), .B(input3[6]), .Z(
        Midori_add_Result_Start3[6]) );
  XOR2_X1 Midori_U188 ( .A(wk_share3[63]), .B(input3[63]), .Z(
        Midori_add_Result_Start3[63]) );
  XOR2_X1 Midori_U187 ( .A(wk_share3[62]), .B(input3[62]), .Z(
        Midori_add_Result_Start3[62]) );
  XOR2_X1 Midori_U186 ( .A(wk_share3[61]), .B(input3[61]), .Z(
        Midori_add_Result_Start3[61]) );
  XOR2_X1 Midori_U185 ( .A(wk_share3[60]), .B(input3[60]), .Z(
        Midori_add_Result_Start3[60]) );
  XOR2_X1 Midori_U184 ( .A(wk_share3[5]), .B(input3[5]), .Z(
        Midori_add_Result_Start3[5]) );
  XOR2_X1 Midori_U183 ( .A(wk_share3[59]), .B(input3[59]), .Z(
        Midori_add_Result_Start3[59]) );
  XOR2_X1 Midori_U182 ( .A(wk_share3[58]), .B(input3[58]), .Z(
        Midori_add_Result_Start3[58]) );
  XOR2_X1 Midori_U181 ( .A(wk_share3[57]), .B(input3[57]), .Z(
        Midori_add_Result_Start3[57]) );
  XOR2_X1 Midori_U180 ( .A(wk_share3[56]), .B(input3[56]), .Z(
        Midori_add_Result_Start3[56]) );
  XOR2_X1 Midori_U179 ( .A(wk_share3[55]), .B(input3[55]), .Z(
        Midori_add_Result_Start3[55]) );
  XOR2_X1 Midori_U178 ( .A(wk_share3[54]), .B(input3[54]), .Z(
        Midori_add_Result_Start3[54]) );
  XOR2_X1 Midori_U177 ( .A(wk_share3[53]), .B(input3[53]), .Z(
        Midori_add_Result_Start3[53]) );
  XOR2_X1 Midori_U176 ( .A(wk_share3[52]), .B(input3[52]), .Z(
        Midori_add_Result_Start3[52]) );
  XOR2_X1 Midori_U175 ( .A(wk_share3[51]), .B(input3[51]), .Z(
        Midori_add_Result_Start3[51]) );
  XOR2_X1 Midori_U174 ( .A(wk_share3[50]), .B(input3[50]), .Z(
        Midori_add_Result_Start3[50]) );
  XOR2_X1 Midori_U173 ( .A(wk_share3[4]), .B(input3[4]), .Z(
        Midori_add_Result_Start3[4]) );
  XOR2_X1 Midori_U172 ( .A(wk_share3[49]), .B(input3[49]), .Z(
        Midori_add_Result_Start3[49]) );
  XOR2_X1 Midori_U171 ( .A(wk_share3[48]), .B(input3[48]), .Z(
        Midori_add_Result_Start3[48]) );
  XOR2_X1 Midori_U170 ( .A(wk_share3[47]), .B(input3[47]), .Z(
        Midori_add_Result_Start3[47]) );
  XOR2_X1 Midori_U169 ( .A(wk_share3[46]), .B(input3[46]), .Z(
        Midori_add_Result_Start3[46]) );
  XOR2_X1 Midori_U168 ( .A(wk_share3[45]), .B(input3[45]), .Z(
        Midori_add_Result_Start3[45]) );
  XOR2_X1 Midori_U167 ( .A(wk_share3[44]), .B(input3[44]), .Z(
        Midori_add_Result_Start3[44]) );
  XOR2_X1 Midori_U166 ( .A(wk_share3[43]), .B(input3[43]), .Z(
        Midori_add_Result_Start3[43]) );
  XOR2_X1 Midori_U165 ( .A(wk_share3[42]), .B(input3[42]), .Z(
        Midori_add_Result_Start3[42]) );
  XOR2_X1 Midori_U164 ( .A(wk_share3[41]), .B(input3[41]), .Z(
        Midori_add_Result_Start3[41]) );
  XOR2_X1 Midori_U163 ( .A(wk_share3[40]), .B(input3[40]), .Z(
        Midori_add_Result_Start3[40]) );
  XOR2_X1 Midori_U162 ( .A(wk_share3[3]), .B(input3[3]), .Z(
        Midori_add_Result_Start3[3]) );
  XOR2_X1 Midori_U161 ( .A(wk_share3[39]), .B(input3[39]), .Z(
        Midori_add_Result_Start3[39]) );
  XOR2_X1 Midori_U160 ( .A(wk_share3[38]), .B(input3[38]), .Z(
        Midori_add_Result_Start3[38]) );
  XOR2_X1 Midori_U159 ( .A(wk_share3[37]), .B(input3[37]), .Z(
        Midori_add_Result_Start3[37]) );
  XOR2_X1 Midori_U158 ( .A(wk_share3[36]), .B(input3[36]), .Z(
        Midori_add_Result_Start3[36]) );
  XOR2_X1 Midori_U157 ( .A(wk_share3[35]), .B(input3[35]), .Z(
        Midori_add_Result_Start3[35]) );
  XOR2_X1 Midori_U156 ( .A(wk_share3[34]), .B(input3[34]), .Z(
        Midori_add_Result_Start3[34]) );
  XOR2_X1 Midori_U155 ( .A(wk_share3[33]), .B(input3[33]), .Z(
        Midori_add_Result_Start3[33]) );
  XOR2_X1 Midori_U154 ( .A(wk_share3[32]), .B(input3[32]), .Z(
        Midori_add_Result_Start3[32]) );
  XOR2_X1 Midori_U153 ( .A(wk_share3[31]), .B(input3[31]), .Z(
        Midori_add_Result_Start3[31]) );
  XOR2_X1 Midori_U152 ( .A(wk_share3[30]), .B(input3[30]), .Z(
        Midori_add_Result_Start3[30]) );
  XOR2_X1 Midori_U151 ( .A(wk_share3[2]), .B(input3[2]), .Z(
        Midori_add_Result_Start3[2]) );
  XOR2_X1 Midori_U150 ( .A(wk_share3[29]), .B(input3[29]), .Z(
        Midori_add_Result_Start3[29]) );
  XOR2_X1 Midori_U149 ( .A(wk_share3[28]), .B(input3[28]), .Z(
        Midori_add_Result_Start3[28]) );
  XOR2_X1 Midori_U148 ( .A(wk_share3[27]), .B(input3[27]), .Z(
        Midori_add_Result_Start3[27]) );
  XOR2_X1 Midori_U147 ( .A(wk_share3[26]), .B(input3[26]), .Z(
        Midori_add_Result_Start3[26]) );
  XOR2_X1 Midori_U146 ( .A(wk_share3[25]), .B(input3[25]), .Z(
        Midori_add_Result_Start3[25]) );
  XOR2_X1 Midori_U145 ( .A(wk_share3[24]), .B(input3[24]), .Z(
        Midori_add_Result_Start3[24]) );
  XOR2_X1 Midori_U144 ( .A(wk_share3[23]), .B(input3[23]), .Z(
        Midori_add_Result_Start3[23]) );
  XOR2_X1 Midori_U143 ( .A(wk_share3[22]), .B(input3[22]), .Z(
        Midori_add_Result_Start3[22]) );
  XOR2_X1 Midori_U142 ( .A(wk_share3[21]), .B(input3[21]), .Z(
        Midori_add_Result_Start3[21]) );
  XOR2_X1 Midori_U141 ( .A(wk_share3[20]), .B(input3[20]), .Z(
        Midori_add_Result_Start3[20]) );
  XOR2_X1 Midori_U140 ( .A(wk_share3[1]), .B(input3[1]), .Z(
        Midori_add_Result_Start3[1]) );
  XOR2_X1 Midori_U139 ( .A(wk_share3[19]), .B(input3[19]), .Z(
        Midori_add_Result_Start3[19]) );
  XOR2_X1 Midori_U138 ( .A(wk_share3[18]), .B(input3[18]), .Z(
        Midori_add_Result_Start3[18]) );
  XOR2_X1 Midori_U137 ( .A(wk_share3[17]), .B(input3[17]), .Z(
        Midori_add_Result_Start3[17]) );
  XOR2_X1 Midori_U136 ( .A(wk_share3[16]), .B(input3[16]), .Z(
        Midori_add_Result_Start3[16]) );
  XOR2_X1 Midori_U135 ( .A(wk_share3[15]), .B(input3[15]), .Z(
        Midori_add_Result_Start3[15]) );
  XOR2_X1 Midori_U134 ( .A(wk_share3[14]), .B(input3[14]), .Z(
        Midori_add_Result_Start3[14]) );
  XOR2_X1 Midori_U133 ( .A(wk_share3[13]), .B(input3[13]), .Z(
        Midori_add_Result_Start3[13]) );
  XOR2_X1 Midori_U132 ( .A(wk_share3[12]), .B(input3[12]), .Z(
        Midori_add_Result_Start3[12]) );
  XOR2_X1 Midori_U131 ( .A(wk_share3[11]), .B(input3[11]), .Z(
        Midori_add_Result_Start3[11]) );
  XOR2_X1 Midori_U130 ( .A(wk_share3[10]), .B(input3[10]), .Z(
        Midori_add_Result_Start3[10]) );
  XOR2_X1 Midori_U129 ( .A(wk_share3[0]), .B(input3[0]), .Z(
        Midori_add_Result_Start3[0]) );
  XOR2_X1 Midori_U128 ( .A(wk_share2[9]), .B(input2[9]), .Z(
        Midori_add_Result_Start2[9]) );
  XOR2_X1 Midori_U127 ( .A(wk_share2[8]), .B(input2[8]), .Z(
        Midori_add_Result_Start2[8]) );
  XOR2_X1 Midori_U126 ( .A(wk_share2[7]), .B(input2[7]), .Z(
        Midori_add_Result_Start2[7]) );
  XOR2_X1 Midori_U125 ( .A(wk_share2[6]), .B(input2[6]), .Z(
        Midori_add_Result_Start2[6]) );
  XOR2_X1 Midori_U124 ( .A(wk_share2[63]), .B(input2[63]), .Z(
        Midori_add_Result_Start2[63]) );
  XOR2_X1 Midori_U123 ( .A(wk_share2[62]), .B(input2[62]), .Z(
        Midori_add_Result_Start2[62]) );
  XOR2_X1 Midori_U122 ( .A(wk_share2[61]), .B(input2[61]), .Z(
        Midori_add_Result_Start2[61]) );
  XOR2_X1 Midori_U121 ( .A(wk_share2[60]), .B(input2[60]), .Z(
        Midori_add_Result_Start2[60]) );
  XOR2_X1 Midori_U120 ( .A(wk_share2[5]), .B(input2[5]), .Z(
        Midori_add_Result_Start2[5]) );
  XOR2_X1 Midori_U119 ( .A(wk_share2[59]), .B(input2[59]), .Z(
        Midori_add_Result_Start2[59]) );
  XOR2_X1 Midori_U118 ( .A(wk_share2[58]), .B(input2[58]), .Z(
        Midori_add_Result_Start2[58]) );
  XOR2_X1 Midori_U117 ( .A(wk_share2[57]), .B(input2[57]), .Z(
        Midori_add_Result_Start2[57]) );
  XOR2_X1 Midori_U116 ( .A(wk_share2[56]), .B(input2[56]), .Z(
        Midori_add_Result_Start2[56]) );
  XOR2_X1 Midori_U115 ( .A(wk_share2[55]), .B(input2[55]), .Z(
        Midori_add_Result_Start2[55]) );
  XOR2_X1 Midori_U114 ( .A(wk_share2[54]), .B(input2[54]), .Z(
        Midori_add_Result_Start2[54]) );
  XOR2_X1 Midori_U113 ( .A(wk_share2[53]), .B(input2[53]), .Z(
        Midori_add_Result_Start2[53]) );
  XOR2_X1 Midori_U112 ( .A(wk_share2[52]), .B(input2[52]), .Z(
        Midori_add_Result_Start2[52]) );
  XOR2_X1 Midori_U111 ( .A(wk_share2[51]), .B(input2[51]), .Z(
        Midori_add_Result_Start2[51]) );
  XOR2_X1 Midori_U110 ( .A(wk_share2[50]), .B(input2[50]), .Z(
        Midori_add_Result_Start2[50]) );
  XOR2_X1 Midori_U109 ( .A(wk_share2[4]), .B(input2[4]), .Z(
        Midori_add_Result_Start2[4]) );
  XOR2_X1 Midori_U108 ( .A(wk_share2[49]), .B(input2[49]), .Z(
        Midori_add_Result_Start2[49]) );
  XOR2_X1 Midori_U107 ( .A(wk_share2[48]), .B(input2[48]), .Z(
        Midori_add_Result_Start2[48]) );
  XOR2_X1 Midori_U106 ( .A(wk_share2[47]), .B(input2[47]), .Z(
        Midori_add_Result_Start2[47]) );
  XOR2_X1 Midori_U105 ( .A(wk_share2[46]), .B(input2[46]), .Z(
        Midori_add_Result_Start2[46]) );
  XOR2_X1 Midori_U104 ( .A(wk_share2[45]), .B(input2[45]), .Z(
        Midori_add_Result_Start2[45]) );
  XOR2_X1 Midori_U103 ( .A(wk_share2[44]), .B(input2[44]), .Z(
        Midori_add_Result_Start2[44]) );
  XOR2_X1 Midori_U102 ( .A(wk_share2[43]), .B(input2[43]), .Z(
        Midori_add_Result_Start2[43]) );
  XOR2_X1 Midori_U101 ( .A(wk_share2[42]), .B(input2[42]), .Z(
        Midori_add_Result_Start2[42]) );
  XOR2_X1 Midori_U100 ( .A(wk_share2[41]), .B(input2[41]), .Z(
        Midori_add_Result_Start2[41]) );
  XOR2_X1 Midori_U99 ( .A(wk_share2[40]), .B(input2[40]), .Z(
        Midori_add_Result_Start2[40]) );
  XOR2_X1 Midori_U98 ( .A(wk_share2[3]), .B(input2[3]), .Z(
        Midori_add_Result_Start2[3]) );
  XOR2_X1 Midori_U97 ( .A(wk_share2[39]), .B(input2[39]), .Z(
        Midori_add_Result_Start2[39]) );
  XOR2_X1 Midori_U96 ( .A(wk_share2[38]), .B(input2[38]), .Z(
        Midori_add_Result_Start2[38]) );
  XOR2_X1 Midori_U95 ( .A(wk_share2[37]), .B(input2[37]), .Z(
        Midori_add_Result_Start2[37]) );
  XOR2_X1 Midori_U94 ( .A(wk_share2[36]), .B(input2[36]), .Z(
        Midori_add_Result_Start2[36]) );
  XOR2_X1 Midori_U93 ( .A(wk_share2[35]), .B(input2[35]), .Z(
        Midori_add_Result_Start2[35]) );
  XOR2_X1 Midori_U92 ( .A(wk_share2[34]), .B(input2[34]), .Z(
        Midori_add_Result_Start2[34]) );
  XOR2_X1 Midori_U91 ( .A(wk_share2[33]), .B(input2[33]), .Z(
        Midori_add_Result_Start2[33]) );
  XOR2_X1 Midori_U90 ( .A(wk_share2[32]), .B(input2[32]), .Z(
        Midori_add_Result_Start2[32]) );
  XOR2_X1 Midori_U89 ( .A(wk_share2[31]), .B(input2[31]), .Z(
        Midori_add_Result_Start2[31]) );
  XOR2_X1 Midori_U88 ( .A(wk_share2[30]), .B(input2[30]), .Z(
        Midori_add_Result_Start2[30]) );
  XOR2_X1 Midori_U87 ( .A(wk_share2[2]), .B(input2[2]), .Z(
        Midori_add_Result_Start2[2]) );
  XOR2_X1 Midori_U86 ( .A(wk_share2[29]), .B(input2[29]), .Z(
        Midori_add_Result_Start2[29]) );
  XOR2_X1 Midori_U85 ( .A(wk_share2[28]), .B(input2[28]), .Z(
        Midori_add_Result_Start2[28]) );
  XOR2_X1 Midori_U84 ( .A(wk_share2[27]), .B(input2[27]), .Z(
        Midori_add_Result_Start2[27]) );
  XOR2_X1 Midori_U83 ( .A(wk_share2[26]), .B(input2[26]), .Z(
        Midori_add_Result_Start2[26]) );
  XOR2_X1 Midori_U82 ( .A(wk_share2[25]), .B(input2[25]), .Z(
        Midori_add_Result_Start2[25]) );
  XOR2_X1 Midori_U81 ( .A(wk_share2[24]), .B(input2[24]), .Z(
        Midori_add_Result_Start2[24]) );
  XOR2_X1 Midori_U80 ( .A(wk_share2[23]), .B(input2[23]), .Z(
        Midori_add_Result_Start2[23]) );
  XOR2_X1 Midori_U79 ( .A(wk_share2[22]), .B(input2[22]), .Z(
        Midori_add_Result_Start2[22]) );
  XOR2_X1 Midori_U78 ( .A(wk_share2[21]), .B(input2[21]), .Z(
        Midori_add_Result_Start2[21]) );
  XOR2_X1 Midori_U77 ( .A(wk_share2[20]), .B(input2[20]), .Z(
        Midori_add_Result_Start2[20]) );
  XOR2_X1 Midori_U76 ( .A(wk_share2[1]), .B(input2[1]), .Z(
        Midori_add_Result_Start2[1]) );
  XOR2_X1 Midori_U75 ( .A(wk_share2[19]), .B(input2[19]), .Z(
        Midori_add_Result_Start2[19]) );
  XOR2_X1 Midori_U74 ( .A(wk_share2[18]), .B(input2[18]), .Z(
        Midori_add_Result_Start2[18]) );
  XOR2_X1 Midori_U73 ( .A(wk_share2[17]), .B(input2[17]), .Z(
        Midori_add_Result_Start2[17]) );
  XOR2_X1 Midori_U72 ( .A(wk_share2[16]), .B(input2[16]), .Z(
        Midori_add_Result_Start2[16]) );
  XOR2_X1 Midori_U71 ( .A(wk_share2[15]), .B(input2[15]), .Z(
        Midori_add_Result_Start2[15]) );
  XOR2_X1 Midori_U70 ( .A(wk_share2[14]), .B(input2[14]), .Z(
        Midori_add_Result_Start2[14]) );
  XOR2_X1 Midori_U69 ( .A(wk_share2[13]), .B(input2[13]), .Z(
        Midori_add_Result_Start2[13]) );
  XOR2_X1 Midori_U68 ( .A(wk_share2[12]), .B(input2[12]), .Z(
        Midori_add_Result_Start2[12]) );
  XOR2_X1 Midori_U67 ( .A(wk_share2[11]), .B(input2[11]), .Z(
        Midori_add_Result_Start2[11]) );
  XOR2_X1 Midori_U66 ( .A(wk_share2[10]), .B(input2[10]), .Z(
        Midori_add_Result_Start2[10]) );
  XOR2_X1 Midori_U65 ( .A(wk_share2[0]), .B(input2[0]), .Z(
        Midori_add_Result_Start2[0]) );
  XOR2_X1 Midori_U64 ( .A(wk_share1[9]), .B(input1[9]), .Z(
        Midori_add_Result_Start1[9]) );
  XOR2_X1 Midori_U63 ( .A(wk_share1[8]), .B(input1[8]), .Z(
        Midori_add_Result_Start1[8]) );
  XOR2_X1 Midori_U62 ( .A(wk_share1[7]), .B(input1[7]), .Z(
        Midori_add_Result_Start1[7]) );
  XOR2_X1 Midori_U61 ( .A(wk_share1[6]), .B(input1[6]), .Z(
        Midori_add_Result_Start1[6]) );
  XOR2_X1 Midori_U60 ( .A(wk_share1[63]), .B(input1[63]), .Z(
        Midori_add_Result_Start1[63]) );
  XOR2_X1 Midori_U59 ( .A(wk_share1[62]), .B(input1[62]), .Z(
        Midori_add_Result_Start1[62]) );
  XOR2_X1 Midori_U58 ( .A(wk_share1[61]), .B(input1[61]), .Z(
        Midori_add_Result_Start1[61]) );
  XOR2_X1 Midori_U57 ( .A(wk_share1[60]), .B(input1[60]), .Z(
        Midori_add_Result_Start1[60]) );
  XOR2_X1 Midori_U56 ( .A(wk_share1[5]), .B(input1[5]), .Z(
        Midori_add_Result_Start1[5]) );
  XOR2_X1 Midori_U55 ( .A(wk_share1[59]), .B(input1[59]), .Z(
        Midori_add_Result_Start1[59]) );
  XOR2_X1 Midori_U54 ( .A(wk_share1[58]), .B(input1[58]), .Z(
        Midori_add_Result_Start1[58]) );
  XOR2_X1 Midori_U53 ( .A(wk_share1[57]), .B(input1[57]), .Z(
        Midori_add_Result_Start1[57]) );
  XOR2_X1 Midori_U52 ( .A(wk_share1[56]), .B(input1[56]), .Z(
        Midori_add_Result_Start1[56]) );
  XOR2_X1 Midori_U51 ( .A(wk_share1[55]), .B(input1[55]), .Z(
        Midori_add_Result_Start1[55]) );
  XOR2_X1 Midori_U50 ( .A(wk_share1[54]), .B(input1[54]), .Z(
        Midori_add_Result_Start1[54]) );
  XOR2_X1 Midori_U49 ( .A(wk_share1[53]), .B(input1[53]), .Z(
        Midori_add_Result_Start1[53]) );
  XOR2_X1 Midori_U48 ( .A(wk_share1[52]), .B(input1[52]), .Z(
        Midori_add_Result_Start1[52]) );
  XOR2_X1 Midori_U47 ( .A(wk_share1[51]), .B(input1[51]), .Z(
        Midori_add_Result_Start1[51]) );
  XOR2_X1 Midori_U46 ( .A(wk_share1[50]), .B(input1[50]), .Z(
        Midori_add_Result_Start1[50]) );
  XOR2_X1 Midori_U45 ( .A(wk_share1[4]), .B(input1[4]), .Z(
        Midori_add_Result_Start1[4]) );
  XOR2_X1 Midori_U44 ( .A(wk_share1[49]), .B(input1[49]), .Z(
        Midori_add_Result_Start1[49]) );
  XOR2_X1 Midori_U43 ( .A(wk_share1[48]), .B(input1[48]), .Z(
        Midori_add_Result_Start1[48]) );
  XOR2_X1 Midori_U42 ( .A(wk_share1[47]), .B(input1[47]), .Z(
        Midori_add_Result_Start1[47]) );
  XOR2_X1 Midori_U41 ( .A(wk_share1[46]), .B(input1[46]), .Z(
        Midori_add_Result_Start1[46]) );
  XOR2_X1 Midori_U40 ( .A(wk_share1[45]), .B(input1[45]), .Z(
        Midori_add_Result_Start1[45]) );
  XOR2_X1 Midori_U39 ( .A(wk_share1[44]), .B(input1[44]), .Z(
        Midori_add_Result_Start1[44]) );
  XOR2_X1 Midori_U38 ( .A(wk_share1[43]), .B(input1[43]), .Z(
        Midori_add_Result_Start1[43]) );
  XOR2_X1 Midori_U37 ( .A(wk_share1[42]), .B(input1[42]), .Z(
        Midori_add_Result_Start1[42]) );
  XOR2_X1 Midori_U36 ( .A(wk_share1[41]), .B(input1[41]), .Z(
        Midori_add_Result_Start1[41]) );
  XOR2_X1 Midori_U35 ( .A(wk_share1[40]), .B(input1[40]), .Z(
        Midori_add_Result_Start1[40]) );
  XOR2_X1 Midori_U34 ( .A(wk_share1[3]), .B(input1[3]), .Z(
        Midori_add_Result_Start1[3]) );
  XOR2_X1 Midori_U33 ( .A(wk_share1[39]), .B(input1[39]), .Z(
        Midori_add_Result_Start1[39]) );
  XOR2_X1 Midori_U32 ( .A(wk_share1[38]), .B(input1[38]), .Z(
        Midori_add_Result_Start1[38]) );
  XOR2_X1 Midori_U31 ( .A(wk_share1[37]), .B(input1[37]), .Z(
        Midori_add_Result_Start1[37]) );
  XOR2_X1 Midori_U30 ( .A(wk_share1[36]), .B(input1[36]), .Z(
        Midori_add_Result_Start1[36]) );
  XOR2_X1 Midori_U29 ( .A(wk_share1[35]), .B(input1[35]), .Z(
        Midori_add_Result_Start1[35]) );
  XOR2_X1 Midori_U28 ( .A(wk_share1[34]), .B(input1[34]), .Z(
        Midori_add_Result_Start1[34]) );
  XOR2_X1 Midori_U27 ( .A(wk_share1[33]), .B(input1[33]), .Z(
        Midori_add_Result_Start1[33]) );
  XOR2_X1 Midori_U26 ( .A(wk_share1[32]), .B(input1[32]), .Z(
        Midori_add_Result_Start1[32]) );
  XOR2_X1 Midori_U25 ( .A(wk_share1[31]), .B(input1[31]), .Z(
        Midori_add_Result_Start1[31]) );
  XOR2_X1 Midori_U24 ( .A(wk_share1[30]), .B(input1[30]), .Z(
        Midori_add_Result_Start1[30]) );
  XOR2_X1 Midori_U23 ( .A(wk_share1[2]), .B(input1[2]), .Z(
        Midori_add_Result_Start1[2]) );
  XOR2_X1 Midori_U22 ( .A(wk_share1[29]), .B(input1[29]), .Z(
        Midori_add_Result_Start1[29]) );
  XOR2_X1 Midori_U21 ( .A(wk_share1[28]), .B(input1[28]), .Z(
        Midori_add_Result_Start1[28]) );
  XOR2_X1 Midori_U20 ( .A(wk_share1[27]), .B(input1[27]), .Z(
        Midori_add_Result_Start1[27]) );
  XOR2_X1 Midori_U19 ( .A(wk_share1[26]), .B(input1[26]), .Z(
        Midori_add_Result_Start1[26]) );
  XOR2_X1 Midori_U18 ( .A(wk_share1[25]), .B(input1[25]), .Z(
        Midori_add_Result_Start1[25]) );
  XOR2_X1 Midori_U17 ( .A(wk_share1[24]), .B(input1[24]), .Z(
        Midori_add_Result_Start1[24]) );
  XOR2_X1 Midori_U16 ( .A(wk_share1[23]), .B(input1[23]), .Z(
        Midori_add_Result_Start1[23]) );
  XOR2_X1 Midori_U15 ( .A(wk_share1[22]), .B(input1[22]), .Z(
        Midori_add_Result_Start1[22]) );
  XOR2_X1 Midori_U14 ( .A(wk_share1[21]), .B(input1[21]), .Z(
        Midori_add_Result_Start1[21]) );
  XOR2_X1 Midori_U13 ( .A(wk_share1[20]), .B(input1[20]), .Z(
        Midori_add_Result_Start1[20]) );
  XOR2_X1 Midori_U12 ( .A(wk_share1[1]), .B(input1[1]), .Z(
        Midori_add_Result_Start1[1]) );
  XOR2_X1 Midori_U11 ( .A(wk_share1[19]), .B(input1[19]), .Z(
        Midori_add_Result_Start1[19]) );
  XOR2_X1 Midori_U10 ( .A(wk_share1[18]), .B(input1[18]), .Z(
        Midori_add_Result_Start1[18]) );
  XOR2_X1 Midori_U9 ( .A(wk_share1[17]), .B(input1[17]), .Z(
        Midori_add_Result_Start1[17]) );
  XOR2_X1 Midori_U8 ( .A(wk_share1[16]), .B(input1[16]), .Z(
        Midori_add_Result_Start1[16]) );
  XOR2_X1 Midori_U7 ( .A(wk_share1[15]), .B(input1[15]), .Z(
        Midori_add_Result_Start1[15]) );
  XOR2_X1 Midori_U6 ( .A(wk_share1[14]), .B(input1[14]), .Z(
        Midori_add_Result_Start1[14]) );
  XOR2_X1 Midori_U5 ( .A(wk_share1[13]), .B(input1[13]), .Z(
        Midori_add_Result_Start1[13]) );
  XOR2_X1 Midori_U4 ( .A(wk_share1[12]), .B(input1[12]), .Z(
        Midori_add_Result_Start1[12]) );
  XOR2_X1 Midori_U3 ( .A(wk_share1[11]), .B(input1[11]), .Z(
        Midori_add_Result_Start1[11]) );
  XOR2_X1 Midori_U2 ( .A(wk_share1[10]), .B(input1[10]), .Z(
        Midori_add_Result_Start1[10]) );
  XOR2_X1 Midori_U1 ( .A(wk_share1[0]), .B(input1[0]), .Z(
        Midori_add_Result_Start1[0]) );
  OAI21_X1 Midori_rounds_U1214 ( .B1(Midori_rounds_n2068), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2066), .ZN(Midori_rounds_n789)
         );
  AOI22_X1 Midori_rounds_U1213 ( .A1(reset), .A2(Midori_add_Result_Start1[0]), 
        .B1(Midori_rounds_n2065), .B2(Midori_rounds_SR_Inv_Result1[0]), .ZN(
        Midori_rounds_n2066) );
  XOR2_X1 Midori_rounds_U1212 ( .A(Midori_rounds_SR_Inv_Result1[28]), .B(
        Midori_rounds_n2064), .Z(Midori_rounds_n2068) );
  OAI21_X1 Midori_rounds_U1211 ( .B1(Midori_rounds_n2063), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2062), .ZN(Midori_rounds_n790)
         );
  AOI22_X1 Midori_rounds_U1210 ( .A1(reset), .A2(Midori_add_Result_Start1[4]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[4]), .ZN(
        Midori_rounds_n2062) );
  XOR2_X1 Midori_rounds_U1209 ( .A(Midori_rounds_SR_Inv_Result1[52]), .B(
        Midori_rounds_n2061), .Z(Midori_rounds_n2063) );
  OAI21_X1 Midori_rounds_U1208 ( .B1(Midori_rounds_n2060), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2059), .ZN(Midori_rounds_n791)
         );
  AOI22_X1 Midori_rounds_U1207 ( .A1(reset), .A2(Midori_add_Result_Start1[8]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[8]), .ZN(
        Midori_rounds_n2059) );
  XOR2_X1 Midori_rounds_U1206 ( .A(Midori_rounds_SR_Inv_Result1[8]), .B(
        Midori_rounds_n2058), .Z(Midori_rounds_n2060) );
  OAI21_X1 Midori_rounds_U1205 ( .B1(Midori_rounds_n2057), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2056), .ZN(Midori_rounds_n792)
         );
  AOI22_X1 Midori_rounds_U1204 ( .A1(reset), .A2(Midori_add_Result_Start1[12]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[12]), .ZN(
        Midori_rounds_n2056) );
  XOR2_X1 Midori_rounds_U1203 ( .A(Midori_rounds_SR_Inv_Result1[32]), .B(
        Midori_rounds_n2055), .Z(Midori_rounds_n2057) );
  OAI21_X1 Midori_rounds_U1202 ( .B1(Midori_rounds_n2054), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2053), .ZN(Midori_rounds_n793)
         );
  AOI22_X1 Midori_rounds_U1201 ( .A1(reset), .A2(Midori_add_Result_Start1[16]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[16]), .ZN(
        Midori_rounds_n2053) );
  XOR2_X1 Midori_rounds_U1200 ( .A(Midori_rounds_SR_Inv_Result1[36]), .B(
        Midori_rounds_n2052), .Z(Midori_rounds_n2054) );
  OAI21_X1 Midori_rounds_U1199 ( .B1(Midori_rounds_n2051), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2050), .ZN(Midori_rounds_n794)
         );
  AOI22_X1 Midori_rounds_U1198 ( .A1(reset), .A2(Midori_add_Result_Start1[20]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[20]), .ZN(
        Midori_rounds_n2050) );
  XOR2_X1 Midori_rounds_U1197 ( .A(Midori_rounds_SR_Inv_Result1[12]), .B(
        Midori_rounds_n2049), .Z(Midori_rounds_n2051) );
  OAI21_X1 Midori_rounds_U1196 ( .B1(Midori_rounds_n2048), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2047), .ZN(Midori_rounds_n795)
         );
  AOI22_X1 Midori_rounds_U1195 ( .A1(reset), .A2(Midori_add_Result_Start1[24]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[24]), .ZN(
        Midori_rounds_n2047) );
  XOR2_X1 Midori_rounds_U1194 ( .A(Midori_rounds_SR_Inv_Result1[48]), .B(
        Midori_rounds_n2046), .Z(Midori_rounds_n2048) );
  OAI21_X1 Midori_rounds_U1193 ( .B1(Midori_rounds_n2045), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2044), .ZN(Midori_rounds_n796)
         );
  AOI22_X1 Midori_rounds_U1192 ( .A1(reset), .A2(Midori_add_Result_Start1[28]), 
        .B1(Midori_rounds_n2065), .B2(Midori_rounds_SR_Inv_Result1[28]), .ZN(
        Midori_rounds_n2044) );
  XOR2_X1 Midori_rounds_U1191 ( .A(Midori_rounds_SR_Inv_Result1[24]), .B(
        Midori_rounds_n2043), .Z(Midori_rounds_n2045) );
  OAI21_X1 Midori_rounds_U1190 ( .B1(Midori_rounds_n2042), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2041), .ZN(Midori_rounds_n797)
         );
  AOI22_X1 Midori_rounds_U1189 ( .A1(reset), .A2(Midori_add_Result_Start1[32]), 
        .B1(Midori_rounds_n2065), .B2(Midori_rounds_SR_Inv_Result1[32]), .ZN(
        Midori_rounds_n2041) );
  XOR2_X1 Midori_rounds_U1188 ( .A(Midori_rounds_SR_Inv_Result1[56]), .B(
        Midori_rounds_n2040), .Z(Midori_rounds_n2042) );
  OAI21_X1 Midori_rounds_U1187 ( .B1(Midori_rounds_n2039), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2038), .ZN(Midori_rounds_n798)
         );
  AOI22_X1 Midori_rounds_U1186 ( .A1(reset), .A2(Midori_add_Result_Start1[36]), 
        .B1(Midori_rounds_n2065), .B2(Midori_rounds_SR_Inv_Result1[36]), .ZN(
        Midori_rounds_n2038) );
  XOR2_X1 Midori_rounds_U1185 ( .A(Midori_rounds_SR_Inv_Result1[16]), .B(
        Midori_rounds_n2037), .Z(Midori_rounds_n2039) );
  OAI21_X1 Midori_rounds_U1184 ( .B1(Midori_rounds_n2036), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2035), .ZN(Midori_rounds_n799)
         );
  AOI22_X1 Midori_rounds_U1183 ( .A1(reset), .A2(Midori_add_Result_Start1[40]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[40]), .ZN(
        Midori_rounds_n2035) );
  XOR2_X1 Midori_rounds_U1182 ( .A(Midori_rounds_SR_Inv_Result1[44]), .B(
        Midori_rounds_n2034), .Z(Midori_rounds_n2036) );
  OAI21_X1 Midori_rounds_U1181 ( .B1(Midori_rounds_n2033), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2032), .ZN(Midori_rounds_n800)
         );
  AOI22_X1 Midori_rounds_U1180 ( .A1(reset), .A2(Midori_add_Result_Start1[44]), 
        .B1(Midori_rounds_n2065), .B2(Midori_rounds_SR_Inv_Result1[44]), .ZN(
        Midori_rounds_n2032) );
  XOR2_X1 Midori_rounds_U1179 ( .A(Midori_rounds_SR_Inv_Result1[4]), .B(
        Midori_rounds_n2031), .Z(Midori_rounds_n2033) );
  OAI21_X1 Midori_rounds_U1178 ( .B1(Midori_rounds_n2030), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2029), .ZN(Midori_rounds_n801)
         );
  AOI22_X1 Midori_rounds_U1177 ( .A1(reset), .A2(Midori_add_Result_Start1[48]), 
        .B1(Midori_rounds_n2065), .B2(Midori_rounds_SR_Inv_Result1[48]), .ZN(
        Midori_rounds_n2029) );
  XOR2_X1 Midori_rounds_U1176 ( .A(Midori_rounds_SR_Inv_Result1[0]), .B(
        Midori_rounds_n2028), .Z(Midori_rounds_n2030) );
  OAI21_X1 Midori_rounds_U1175 ( .B1(Midori_rounds_n2027), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2026), .ZN(Midori_rounds_n802)
         );
  AOI22_X1 Midori_rounds_U1174 ( .A1(reset), .A2(Midori_add_Result_Start1[52]), 
        .B1(Midori_rounds_n2065), .B2(Midori_rounds_SR_Inv_Result1[52]), .ZN(
        Midori_rounds_n2026) );
  XOR2_X1 Midori_rounds_U1173 ( .A(Midori_rounds_SR_Inv_Result1[40]), .B(
        Midori_rounds_n2025), .Z(Midori_rounds_n2027) );
  OAI21_X1 Midori_rounds_U1172 ( .B1(Midori_rounds_n2024), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2023), .ZN(Midori_rounds_n803)
         );
  AOI22_X1 Midori_rounds_U1171 ( .A1(reset), .A2(Midori_add_Result_Start1[56]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[56]), .ZN(
        Midori_rounds_n2023) );
  XOR2_X1 Midori_rounds_U1170 ( .A(Midori_rounds_SR_Inv_Result1[20]), .B(
        Midori_rounds_n2022), .Z(Midori_rounds_n2024) );
  OAI21_X1 Midori_rounds_U1169 ( .B1(Midori_rounds_n2021), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2020), .ZN(Midori_rounds_n804)
         );
  AOI22_X1 Midori_rounds_U1168 ( .A1(reset), .A2(Midori_add_Result_Start1[60]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[60]), .ZN(
        Midori_rounds_n2020) );
  XOR2_X1 Midori_rounds_U1167 ( .A(Midori_rounds_SR_Inv_Result1[60]), .B(
        Midori_rounds_n2019), .Z(Midori_rounds_n2021) );
  OAI21_X1 Midori_rounds_U1166 ( .B1(Midori_rounds_n2018), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2017), .ZN(Midori_rounds_n805)
         );
  AOI22_X1 Midori_rounds_U1165 ( .A1(reset), .A2(Midori_add_Result_Start1[1]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[1]), .ZN(
        Midori_rounds_n2017) );
  XOR2_X1 Midori_rounds_U1164 ( .A(Midori_rounds_SR_Inv_Result1[29]), .B(
        Midori_rounds_n2016), .Z(Midori_rounds_n2018) );
  OAI21_X1 Midori_rounds_U1163 ( .B1(Midori_rounds_n2015), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2014), .ZN(Midori_rounds_n806)
         );
  AOI22_X1 Midori_rounds_U1162 ( .A1(reset), .A2(Midori_add_Result_Start1[2]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[2]), .ZN(
        Midori_rounds_n2014) );
  XOR2_X1 Midori_rounds_U1161 ( .A(Midori_rounds_SR_Inv_Result1[30]), .B(
        Midori_rounds_n2013), .Z(Midori_rounds_n2015) );
  OAI21_X1 Midori_rounds_U1160 ( .B1(Midori_rounds_n2012), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2011), .ZN(
        Midori_rounds_sub_Sub_0_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1159 ( .A1(reset), .A2(Midori_add_Result_Start1[3]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[3]), .ZN(
        Midori_rounds_n2011) );
  XOR2_X1 Midori_rounds_U1158 ( .A(Midori_rounds_SR_Inv_Result1[31]), .B(
        Midori_rounds_n2010), .Z(Midori_rounds_n2012) );
  OAI21_X1 Midori_rounds_U1157 ( .B1(Midori_rounds_n2009), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2008), .ZN(Midori_rounds_n808)
         );
  AOI22_X1 Midori_rounds_U1156 ( .A1(reset), .A2(Midori_add_Result_Start1[5]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[5]), .ZN(
        Midori_rounds_n2008) );
  XOR2_X1 Midori_rounds_U1155 ( .A(Midori_rounds_SR_Inv_Result1[53]), .B(
        Midori_rounds_n2007), .Z(Midori_rounds_n2009) );
  OAI21_X1 Midori_rounds_U1154 ( .B1(Midori_rounds_n2006), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2005), .ZN(Midori_rounds_n809)
         );
  AOI22_X1 Midori_rounds_U1153 ( .A1(reset), .A2(Midori_add_Result_Start1[6]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[6]), .ZN(
        Midori_rounds_n2005) );
  XOR2_X1 Midori_rounds_U1152 ( .A(Midori_rounds_SR_Inv_Result1[54]), .B(
        Midori_rounds_n2004), .Z(Midori_rounds_n2006) );
  OAI21_X1 Midori_rounds_U1151 ( .B1(Midori_rounds_n2003), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2002), .ZN(
        Midori_rounds_sub_Sub_1_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1150 ( .A1(reset), .A2(Midori_add_Result_Start1[7]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[7]), .ZN(
        Midori_rounds_n2002) );
  XOR2_X1 Midori_rounds_U1149 ( .A(Midori_rounds_SR_Inv_Result1[55]), .B(
        Midori_rounds_n2001), .Z(Midori_rounds_n2003) );
  OAI21_X1 Midori_rounds_U1148 ( .B1(Midori_rounds_n2000), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1999), .ZN(Midori_rounds_n811)
         );
  AOI22_X1 Midori_rounds_U1147 ( .A1(reset), .A2(Midori_add_Result_Start1[9]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[9]), .ZN(
        Midori_rounds_n1999) );
  XOR2_X1 Midori_rounds_U1146 ( .A(Midori_rounds_SR_Inv_Result1[9]), .B(
        Midori_rounds_n1998), .Z(Midori_rounds_n2000) );
  OAI21_X1 Midori_rounds_U1145 ( .B1(Midori_rounds_n1997), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1996), .ZN(Midori_rounds_n812)
         );
  AOI22_X1 Midori_rounds_U1144 ( .A1(reset), .A2(Midori_add_Result_Start1[10]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[10]), .ZN(
        Midori_rounds_n1996) );
  XOR2_X1 Midori_rounds_U1143 ( .A(Midori_rounds_SR_Inv_Result1[10]), .B(
        Midori_rounds_n1995), .Z(Midori_rounds_n1997) );
  OAI21_X1 Midori_rounds_U1142 ( .B1(Midori_rounds_n1994), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1993), .ZN(
        Midori_rounds_sub_Sub_2_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1141 ( .A1(reset), .A2(Midori_add_Result_Start1[11]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[11]), .ZN(
        Midori_rounds_n1993) );
  XOR2_X1 Midori_rounds_U1140 ( .A(Midori_rounds_SR_Inv_Result1[11]), .B(
        Midori_rounds_n1992), .Z(Midori_rounds_n1994) );
  OAI21_X1 Midori_rounds_U1139 ( .B1(Midori_rounds_n1991), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1990), .ZN(Midori_rounds_n814)
         );
  AOI22_X1 Midori_rounds_U1138 ( .A1(reset), .A2(Midori_add_Result_Start1[13]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[13]), .ZN(
        Midori_rounds_n1990) );
  XOR2_X1 Midori_rounds_U1137 ( .A(Midori_rounds_SR_Inv_Result1[33]), .B(
        Midori_rounds_n1989), .Z(Midori_rounds_n1991) );
  OAI21_X1 Midori_rounds_U1136 ( .B1(Midori_rounds_n1988), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1987), .ZN(Midori_rounds_n815)
         );
  AOI22_X1 Midori_rounds_U1135 ( .A1(reset), .A2(Midori_add_Result_Start1[14]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[14]), .ZN(
        Midori_rounds_n1987) );
  XOR2_X1 Midori_rounds_U1134 ( .A(Midori_rounds_SR_Inv_Result1[34]), .B(
        Midori_rounds_n1986), .Z(Midori_rounds_n1988) );
  OAI21_X1 Midori_rounds_U1133 ( .B1(Midori_rounds_n1985), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1984), .ZN(
        Midori_rounds_sub_Sub_3_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1132 ( .A1(reset), .A2(Midori_add_Result_Start1[15]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[15]), .ZN(
        Midori_rounds_n1984) );
  XOR2_X1 Midori_rounds_U1131 ( .A(Midori_rounds_SR_Inv_Result1[35]), .B(
        Midori_rounds_n1983), .Z(Midori_rounds_n1985) );
  OAI21_X1 Midori_rounds_U1130 ( .B1(Midori_rounds_n1982), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1981), .ZN(Midori_rounds_n817)
         );
  AOI22_X1 Midori_rounds_U1129 ( .A1(reset), .A2(Midori_add_Result_Start1[17]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[17]), .ZN(
        Midori_rounds_n1981) );
  XOR2_X1 Midori_rounds_U1128 ( .A(Midori_rounds_SR_Inv_Result1[37]), .B(
        Midori_rounds_n1980), .Z(Midori_rounds_n1982) );
  OAI21_X1 Midori_rounds_U1127 ( .B1(Midori_rounds_n1979), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1978), .ZN(Midori_rounds_n818)
         );
  AOI22_X1 Midori_rounds_U1126 ( .A1(reset), .A2(Midori_add_Result_Start1[18]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[18]), .ZN(
        Midori_rounds_n1978) );
  XOR2_X1 Midori_rounds_U1125 ( .A(Midori_rounds_SR_Inv_Result1[38]), .B(
        Midori_rounds_n1977), .Z(Midori_rounds_n1979) );
  OAI21_X1 Midori_rounds_U1124 ( .B1(Midori_rounds_n1976), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1975), .ZN(
        Midori_rounds_sub_Sub_4_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1123 ( .A1(reset), .A2(Midori_add_Result_Start1[19]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[19]), .ZN(
        Midori_rounds_n1975) );
  XOR2_X1 Midori_rounds_U1122 ( .A(Midori_rounds_SR_Inv_Result1[39]), .B(
        Midori_rounds_n1974), .Z(Midori_rounds_n1976) );
  OAI21_X1 Midori_rounds_U1121 ( .B1(Midori_rounds_n1973), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1972), .ZN(Midori_rounds_n820)
         );
  AOI22_X1 Midori_rounds_U1120 ( .A1(reset), .A2(Midori_add_Result_Start1[21]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[21]), .ZN(
        Midori_rounds_n1972) );
  XOR2_X1 Midori_rounds_U1119 ( .A(Midori_rounds_SR_Inv_Result1[13]), .B(
        Midori_rounds_n1971), .Z(Midori_rounds_n1973) );
  OAI21_X1 Midori_rounds_U1118 ( .B1(Midori_rounds_n1970), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1969), .ZN(Midori_rounds_n821)
         );
  AOI22_X1 Midori_rounds_U1117 ( .A1(reset), .A2(Midori_add_Result_Start1[22]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[22]), .ZN(
        Midori_rounds_n1969) );
  XOR2_X1 Midori_rounds_U1116 ( .A(Midori_rounds_SR_Inv_Result1[14]), .B(
        Midori_rounds_n1968), .Z(Midori_rounds_n1970) );
  OAI21_X1 Midori_rounds_U1115 ( .B1(Midori_rounds_n1967), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1966), .ZN(
        Midori_rounds_sub_Sub_5_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1114 ( .A1(reset), .A2(Midori_add_Result_Start1[23]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[23]), .ZN(
        Midori_rounds_n1966) );
  XOR2_X1 Midori_rounds_U1113 ( .A(Midori_rounds_SR_Inv_Result1[15]), .B(
        Midori_rounds_n1965), .Z(Midori_rounds_n1967) );
  OAI21_X1 Midori_rounds_U1112 ( .B1(Midori_rounds_n1964), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1963), .ZN(Midori_rounds_n823)
         );
  AOI22_X1 Midori_rounds_U1111 ( .A1(reset), .A2(Midori_add_Result_Start1[25]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[25]), .ZN(
        Midori_rounds_n1963) );
  XOR2_X1 Midori_rounds_U1110 ( .A(Midori_rounds_SR_Inv_Result1[49]), .B(
        Midori_rounds_n1962), .Z(Midori_rounds_n1964) );
  OAI21_X1 Midori_rounds_U1109 ( .B1(Midori_rounds_n1961), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1960), .ZN(Midori_rounds_n824)
         );
  AOI22_X1 Midori_rounds_U1108 ( .A1(reset), .A2(Midori_add_Result_Start1[26]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[26]), .ZN(
        Midori_rounds_n1960) );
  XOR2_X1 Midori_rounds_U1107 ( .A(Midori_rounds_SR_Inv_Result1[50]), .B(
        Midori_rounds_n1959), .Z(Midori_rounds_n1961) );
  OAI21_X1 Midori_rounds_U1106 ( .B1(Midori_rounds_n1958), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1957), .ZN(
        Midori_rounds_sub_Sub_6_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1105 ( .A1(reset), .A2(Midori_add_Result_Start1[27]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[27]), .ZN(
        Midori_rounds_n1957) );
  XOR2_X1 Midori_rounds_U1104 ( .A(Midori_rounds_SR_Inv_Result1[51]), .B(
        Midori_rounds_n1956), .Z(Midori_rounds_n1958) );
  OAI21_X1 Midori_rounds_U1103 ( .B1(Midori_rounds_n1955), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1954), .ZN(Midori_rounds_n826)
         );
  AOI22_X1 Midori_rounds_U1102 ( .A1(reset), .A2(Midori_add_Result_Start1[29]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[29]), .ZN(
        Midori_rounds_n1954) );
  XOR2_X1 Midori_rounds_U1101 ( .A(Midori_rounds_SR_Inv_Result1[25]), .B(
        Midori_rounds_n1953), .Z(Midori_rounds_n1955) );
  OAI21_X1 Midori_rounds_U1100 ( .B1(Midori_rounds_n1952), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1951), .ZN(Midori_rounds_n827)
         );
  AOI22_X1 Midori_rounds_U1099 ( .A1(reset), .A2(Midori_add_Result_Start1[30]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[30]), .ZN(
        Midori_rounds_n1951) );
  XOR2_X1 Midori_rounds_U1098 ( .A(Midori_rounds_SR_Inv_Result1[26]), .B(
        Midori_rounds_n1950), .Z(Midori_rounds_n1952) );
  OAI21_X1 Midori_rounds_U1097 ( .B1(Midori_rounds_n1949), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1948), .ZN(
        Midori_rounds_sub_Sub_7_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1096 ( .A1(reset), .A2(Midori_add_Result_Start1[31]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[31]), .ZN(
        Midori_rounds_n1948) );
  XOR2_X1 Midori_rounds_U1095 ( .A(Midori_rounds_SR_Inv_Result1[27]), .B(
        Midori_rounds_n1947), .Z(Midori_rounds_n1949) );
  OAI21_X1 Midori_rounds_U1094 ( .B1(Midori_rounds_n1946), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1945), .ZN(Midori_rounds_n829)
         );
  AOI22_X1 Midori_rounds_U1093 ( .A1(reset), .A2(Midori_add_Result_Start1[33]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[33]), .ZN(
        Midori_rounds_n1945) );
  XOR2_X1 Midori_rounds_U1092 ( .A(Midori_rounds_SR_Inv_Result1[57]), .B(
        Midori_rounds_n1944), .Z(Midori_rounds_n1946) );
  OAI21_X1 Midori_rounds_U1091 ( .B1(Midori_rounds_n1943), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1942), .ZN(Midori_rounds_n830)
         );
  AOI22_X1 Midori_rounds_U1090 ( .A1(reset), .A2(Midori_add_Result_Start1[34]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[34]), .ZN(
        Midori_rounds_n1942) );
  XOR2_X1 Midori_rounds_U1089 ( .A(Midori_rounds_SR_Inv_Result1[58]), .B(
        Midori_rounds_n1941), .Z(Midori_rounds_n1943) );
  OAI21_X1 Midori_rounds_U1088 ( .B1(Midori_rounds_n1940), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1939), .ZN(
        Midori_rounds_sub_Sub_8_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1087 ( .A1(reset), .A2(Midori_add_Result_Start1[35]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[35]), .ZN(
        Midori_rounds_n1939) );
  XOR2_X1 Midori_rounds_U1086 ( .A(Midori_rounds_SR_Inv_Result1[59]), .B(
        Midori_rounds_n1938), .Z(Midori_rounds_n1940) );
  OAI21_X1 Midori_rounds_U1085 ( .B1(Midori_rounds_n1937), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1936), .ZN(Midori_rounds_n832)
         );
  AOI22_X1 Midori_rounds_U1084 ( .A1(reset), .A2(Midori_add_Result_Start1[37]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[37]), .ZN(
        Midori_rounds_n1936) );
  XOR2_X1 Midori_rounds_U1083 ( .A(Midori_rounds_SR_Inv_Result1[17]), .B(
        Midori_rounds_n1935), .Z(Midori_rounds_n1937) );
  OAI21_X1 Midori_rounds_U1082 ( .B1(Midori_rounds_n1934), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1933), .ZN(Midori_rounds_n833)
         );
  AOI22_X1 Midori_rounds_U1081 ( .A1(reset), .A2(Midori_add_Result_Start1[38]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[38]), .ZN(
        Midori_rounds_n1933) );
  XOR2_X1 Midori_rounds_U1080 ( .A(Midori_rounds_SR_Inv_Result1[18]), .B(
        Midori_rounds_n1932), .Z(Midori_rounds_n1934) );
  OAI21_X1 Midori_rounds_U1079 ( .B1(Midori_rounds_n1931), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1930), .ZN(
        Midori_rounds_sub_Sub_9_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1078 ( .A1(reset), .A2(Midori_add_Result_Start1[39]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[39]), .ZN(
        Midori_rounds_n1930) );
  XOR2_X1 Midori_rounds_U1077 ( .A(Midori_rounds_SR_Inv_Result1[19]), .B(
        Midori_rounds_n1929), .Z(Midori_rounds_n1931) );
  OAI21_X1 Midori_rounds_U1076 ( .B1(Midori_rounds_n1928), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1927), .ZN(Midori_rounds_n835)
         );
  AOI22_X1 Midori_rounds_U1075 ( .A1(reset), .A2(Midori_add_Result_Start1[41]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[41]), .ZN(
        Midori_rounds_n1927) );
  XOR2_X1 Midori_rounds_U1074 ( .A(Midori_rounds_SR_Inv_Result1[45]), .B(
        Midori_rounds_n1926), .Z(Midori_rounds_n1928) );
  OAI21_X1 Midori_rounds_U1073 ( .B1(Midori_rounds_n1925), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1924), .ZN(Midori_rounds_n836)
         );
  AOI22_X1 Midori_rounds_U1072 ( .A1(reset), .A2(Midori_add_Result_Start1[42]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[42]), .ZN(
        Midori_rounds_n1924) );
  XOR2_X1 Midori_rounds_U1071 ( .A(Midori_rounds_SR_Inv_Result1[46]), .B(
        Midori_rounds_n1923), .Z(Midori_rounds_n1925) );
  OAI21_X1 Midori_rounds_U1070 ( .B1(Midori_rounds_n1922), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1921), .ZN(
        Midori_rounds_sub_Sub_10_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1069 ( .A1(reset), .A2(Midori_add_Result_Start1[43]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[43]), .ZN(
        Midori_rounds_n1921) );
  XOR2_X1 Midori_rounds_U1068 ( .A(Midori_rounds_SR_Inv_Result1[47]), .B(
        Midori_rounds_n1920), .Z(Midori_rounds_n1922) );
  OAI21_X1 Midori_rounds_U1067 ( .B1(Midori_rounds_n1919), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1918), .ZN(Midori_rounds_n838)
         );
  AOI22_X1 Midori_rounds_U1066 ( .A1(reset), .A2(Midori_add_Result_Start1[45]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[45]), .ZN(
        Midori_rounds_n1918) );
  XOR2_X1 Midori_rounds_U1065 ( .A(Midori_rounds_SR_Inv_Result1[5]), .B(
        Midori_rounds_n1917), .Z(Midori_rounds_n1919) );
  OAI21_X1 Midori_rounds_U1064 ( .B1(Midori_rounds_n1916), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1915), .ZN(Midori_rounds_n839)
         );
  AOI22_X1 Midori_rounds_U1063 ( .A1(reset), .A2(Midori_add_Result_Start1[46]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[46]), .ZN(
        Midori_rounds_n1915) );
  XOR2_X1 Midori_rounds_U1062 ( .A(Midori_rounds_SR_Inv_Result1[6]), .B(
        Midori_rounds_n1914), .Z(Midori_rounds_n1916) );
  OAI21_X1 Midori_rounds_U1061 ( .B1(Midori_rounds_n1913), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1912), .ZN(
        Midori_rounds_sub_Sub_11_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1060 ( .A1(reset), .A2(Midori_add_Result_Start1[47]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[47]), .ZN(
        Midori_rounds_n1912) );
  XOR2_X1 Midori_rounds_U1059 ( .A(Midori_rounds_SR_Inv_Result1[7]), .B(
        Midori_rounds_n1911), .Z(Midori_rounds_n1913) );
  OAI21_X1 Midori_rounds_U1058 ( .B1(Midori_rounds_n1910), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1909), .ZN(Midori_rounds_n841)
         );
  AOI22_X1 Midori_rounds_U1057 ( .A1(reset), .A2(Midori_add_Result_Start1[49]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[49]), .ZN(
        Midori_rounds_n1909) );
  XOR2_X1 Midori_rounds_U1056 ( .A(Midori_rounds_SR_Inv_Result1[1]), .B(
        Midori_rounds_n1908), .Z(Midori_rounds_n1910) );
  OAI21_X1 Midori_rounds_U1055 ( .B1(Midori_rounds_n1907), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1906), .ZN(Midori_rounds_n842)
         );
  AOI22_X1 Midori_rounds_U1054 ( .A1(reset), .A2(Midori_add_Result_Start1[50]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[50]), .ZN(
        Midori_rounds_n1906) );
  XOR2_X1 Midori_rounds_U1053 ( .A(Midori_rounds_SR_Inv_Result1[2]), .B(
        Midori_rounds_n1905), .Z(Midori_rounds_n1907) );
  OAI21_X1 Midori_rounds_U1052 ( .B1(Midori_rounds_n1904), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1903), .ZN(
        Midori_rounds_sub_Sub_12_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1051 ( .A1(reset), .A2(Midori_add_Result_Start1[51]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[51]), .ZN(
        Midori_rounds_n1903) );
  XOR2_X1 Midori_rounds_U1050 ( .A(Midori_rounds_SR_Inv_Result1[3]), .B(
        Midori_rounds_n1902), .Z(Midori_rounds_n1904) );
  OAI21_X1 Midori_rounds_U1049 ( .B1(Midori_rounds_n1901), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1900), .ZN(Midori_rounds_n844)
         );
  AOI22_X1 Midori_rounds_U1048 ( .A1(reset), .A2(Midori_add_Result_Start1[53]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[53]), .ZN(
        Midori_rounds_n1900) );
  XOR2_X1 Midori_rounds_U1047 ( .A(Midori_rounds_SR_Inv_Result1[41]), .B(
        Midori_rounds_n1899), .Z(Midori_rounds_n1901) );
  OAI21_X1 Midori_rounds_U1046 ( .B1(Midori_rounds_n1898), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1897), .ZN(Midori_rounds_n845)
         );
  AOI22_X1 Midori_rounds_U1045 ( .A1(reset), .A2(Midori_add_Result_Start1[54]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[54]), .ZN(
        Midori_rounds_n1897) );
  XOR2_X1 Midori_rounds_U1044 ( .A(Midori_rounds_SR_Inv_Result1[42]), .B(
        Midori_rounds_n1896), .Z(Midori_rounds_n1898) );
  OAI21_X1 Midori_rounds_U1043 ( .B1(Midori_rounds_n1895), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1894), .ZN(
        Midori_rounds_sub_Sub_13_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1042 ( .A1(reset), .A2(Midori_add_Result_Start1[55]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[55]), .ZN(
        Midori_rounds_n1894) );
  XOR2_X1 Midori_rounds_U1041 ( .A(Midori_rounds_SR_Inv_Result1[43]), .B(
        Midori_rounds_n1893), .Z(Midori_rounds_n1895) );
  OAI21_X1 Midori_rounds_U1040 ( .B1(Midori_rounds_n1892), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1891), .ZN(Midori_rounds_n847)
         );
  AOI22_X1 Midori_rounds_U1039 ( .A1(reset), .A2(Midori_add_Result_Start1[57]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[57]), .ZN(
        Midori_rounds_n1891) );
  XOR2_X1 Midori_rounds_U1038 ( .A(Midori_rounds_SR_Inv_Result1[21]), .B(
        Midori_rounds_n1890), .Z(Midori_rounds_n1892) );
  OAI21_X1 Midori_rounds_U1037 ( .B1(Midori_rounds_n1889), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1888), .ZN(Midori_rounds_n848)
         );
  AOI22_X1 Midori_rounds_U1036 ( .A1(reset), .A2(Midori_add_Result_Start1[58]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[58]), .ZN(
        Midori_rounds_n1888) );
  XOR2_X1 Midori_rounds_U1035 ( .A(Midori_rounds_SR_Inv_Result1[22]), .B(
        Midori_rounds_n1887), .Z(Midori_rounds_n1889) );
  OAI21_X1 Midori_rounds_U1034 ( .B1(Midori_rounds_n1886), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1885), .ZN(
        Midori_rounds_sub_Sub_14_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1033 ( .A1(reset), .A2(Midori_add_Result_Start1[59]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[59]), .ZN(
        Midori_rounds_n1885) );
  XOR2_X1 Midori_rounds_U1032 ( .A(Midori_rounds_SR_Inv_Result1[23]), .B(
        Midori_rounds_n1884), .Z(Midori_rounds_n1886) );
  OAI21_X1 Midori_rounds_U1031 ( .B1(Midori_rounds_n1883), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1882), .ZN(Midori_rounds_n850)
         );
  AOI22_X1 Midori_rounds_U1030 ( .A1(reset), .A2(Midori_add_Result_Start1[61]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[61]), .ZN(
        Midori_rounds_n1882) );
  XOR2_X1 Midori_rounds_U1029 ( .A(Midori_rounds_SR_Inv_Result1[61]), .B(
        Midori_rounds_n1881), .Z(Midori_rounds_n1883) );
  OAI21_X1 Midori_rounds_U1028 ( .B1(Midori_rounds_n1880), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1879), .ZN(Midori_rounds_n851)
         );
  AOI22_X1 Midori_rounds_U1027 ( .A1(reset), .A2(Midori_add_Result_Start1[62]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[62]), .ZN(
        Midori_rounds_n1879) );
  XOR2_X1 Midori_rounds_U1026 ( .A(Midori_rounds_SR_Inv_Result1[62]), .B(
        Midori_rounds_n1878), .Z(Midori_rounds_n1880) );
  OAI21_X1 Midori_rounds_U1025 ( .B1(Midori_rounds_n1877), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1876), .ZN(
        Midori_rounds_sub_Sub_15_F_in1[2]) );
  AOI22_X1 Midori_rounds_U1024 ( .A1(reset), .A2(Midori_add_Result_Start1[63]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[63]), .ZN(
        Midori_rounds_n1876) );
  XOR2_X1 Midori_rounds_U1023 ( .A(Midori_rounds_SR_Inv_Result1[63]), .B(
        Midori_rounds_n1875), .Z(Midori_rounds_n1877) );
  OAI21_X1 Midori_rounds_U1022 ( .B1(Midori_rounds_n1874), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1873), .ZN(Midori_rounds_n853)
         );
  AOI22_X1 Midori_rounds_U1021 ( .A1(reset), .A2(Midori_add_Result_Start2[0]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[0]), .ZN(
        Midori_rounds_n1873) );
  XOR2_X1 Midori_rounds_U1020 ( .A(Midori_rounds_SR_Inv_Result2[28]), .B(
        Midori_rounds_n1872), .Z(Midori_rounds_n1874) );
  OAI21_X1 Midori_rounds_U1019 ( .B1(Midori_rounds_n1871), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1870), .ZN(
        Midori_rounds_sub_Sub_0_F_in2[0]) );
  AOI22_X1 Midori_rounds_U1018 ( .A1(reset), .A2(Midori_add_Result_Start2[1]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[1]), .ZN(
        Midori_rounds_n1870) );
  XOR2_X1 Midori_rounds_U1017 ( .A(Midori_rounds_SR_Inv_Result2[29]), .B(
        Midori_rounds_n1869), .Z(Midori_rounds_n1871) );
  OAI21_X1 Midori_rounds_U1016 ( .B1(Midori_rounds_n1868), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1867), .ZN(Midori_rounds_n855)
         );
  AOI22_X1 Midori_rounds_U1015 ( .A1(reset), .A2(Midori_add_Result_Start2[2]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[2]), .ZN(
        Midori_rounds_n1867) );
  XOR2_X1 Midori_rounds_U1014 ( .A(Midori_rounds_SR_Inv_Result2[30]), .B(
        Midori_rounds_n1866), .Z(Midori_rounds_n1868) );
  OAI21_X1 Midori_rounds_U1013 ( .B1(Midori_rounds_n1865), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1864), .ZN(
        Midori_rounds_sub_Sub_0_F_in2[2]) );
  AOI22_X1 Midori_rounds_U1012 ( .A1(reset), .A2(Midori_add_Result_Start2[3]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result2[3]), .ZN(
        Midori_rounds_n1864) );
  XOR2_X1 Midori_rounds_U1011 ( .A(Midori_rounds_SR_Inv_Result2[31]), .B(
        Midori_rounds_n1863), .Z(Midori_rounds_n1865) );
  OAI21_X1 Midori_rounds_U1010 ( .B1(Midori_rounds_n1862), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1861), .ZN(Midori_rounds_n857)
         );
  AOI22_X1 Midori_rounds_U1009 ( .A1(reset), .A2(Midori_add_Result_Start2[4]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[4]), .ZN(
        Midori_rounds_n1861) );
  XOR2_X1 Midori_rounds_U1008 ( .A(Midori_rounds_SR_Inv_Result2[52]), .B(
        Midori_rounds_n1860), .Z(Midori_rounds_n1862) );
  OAI21_X1 Midori_rounds_U1007 ( .B1(Midori_rounds_n1859), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1858), .ZN(
        Midori_rounds_sub_Sub_1_F_in2[0]) );
  AOI22_X1 Midori_rounds_U1006 ( .A1(reset), .A2(Midori_add_Result_Start2[5]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[5]), .ZN(
        Midori_rounds_n1858) );
  XOR2_X1 Midori_rounds_U1005 ( .A(Midori_rounds_SR_Inv_Result2[53]), .B(
        Midori_rounds_n1857), .Z(Midori_rounds_n1859) );
  OAI21_X1 Midori_rounds_U1004 ( .B1(Midori_rounds_n1856), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1855), .ZN(Midori_rounds_n859)
         );
  AOI22_X1 Midori_rounds_U1003 ( .A1(reset), .A2(Midori_add_Result_Start2[6]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[6]), .ZN(
        Midori_rounds_n1855) );
  XOR2_X1 Midori_rounds_U1002 ( .A(Midori_rounds_SR_Inv_Result2[54]), .B(
        Midori_rounds_n1854), .Z(Midori_rounds_n1856) );
  OAI21_X1 Midori_rounds_U1001 ( .B1(Midori_rounds_n1853), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1852), .ZN(
        Midori_rounds_sub_Sub_1_F_in2[2]) );
  AOI22_X1 Midori_rounds_U1000 ( .A1(reset), .A2(Midori_add_Result_Start2[7]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[7]), .ZN(
        Midori_rounds_n1852) );
  XOR2_X1 Midori_rounds_U999 ( .A(Midori_rounds_SR_Inv_Result2[55]), .B(
        Midori_rounds_n1851), .Z(Midori_rounds_n1853) );
  OAI21_X1 Midori_rounds_U998 ( .B1(Midori_rounds_n1850), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1849), .ZN(Midori_rounds_n861)
         );
  AOI22_X1 Midori_rounds_U997 ( .A1(reset), .A2(Midori_add_Result_Start2[8]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[8]), .ZN(
        Midori_rounds_n1849) );
  XOR2_X1 Midori_rounds_U996 ( .A(Midori_rounds_SR_Inv_Result2[8]), .B(
        Midori_rounds_n1848), .Z(Midori_rounds_n1850) );
  OAI21_X1 Midori_rounds_U995 ( .B1(Midori_rounds_n1847), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1846), .ZN(
        Midori_rounds_sub_Sub_2_F_in2[0]) );
  AOI22_X1 Midori_rounds_U994 ( .A1(reset), .A2(Midori_add_Result_Start2[9]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result2[9]), .ZN(
        Midori_rounds_n1846) );
  XOR2_X1 Midori_rounds_U993 ( .A(Midori_rounds_SR_Inv_Result2[9]), .B(
        Midori_rounds_n1845), .Z(Midori_rounds_n1847) );
  OAI21_X1 Midori_rounds_U992 ( .B1(Midori_rounds_n1844), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1843), .ZN(Midori_rounds_n863)
         );
  AOI22_X1 Midori_rounds_U991 ( .A1(reset), .A2(Midori_add_Result_Start2[10]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[10]), .ZN(
        Midori_rounds_n1843) );
  XOR2_X1 Midori_rounds_U990 ( .A(Midori_rounds_SR_Inv_Result2[10]), .B(
        Midori_rounds_n1842), .Z(Midori_rounds_n1844) );
  OAI21_X1 Midori_rounds_U989 ( .B1(Midori_rounds_n1841), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1840), .ZN(
        Midori_rounds_sub_Sub_2_F_in2[2]) );
  AOI22_X1 Midori_rounds_U988 ( .A1(reset), .A2(Midori_add_Result_Start2[11]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[11]), .ZN(
        Midori_rounds_n1840) );
  XOR2_X1 Midori_rounds_U987 ( .A(Midori_rounds_SR_Inv_Result2[11]), .B(
        Midori_rounds_n1839), .Z(Midori_rounds_n1841) );
  OAI21_X1 Midori_rounds_U986 ( .B1(Midori_rounds_n1838), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1837), .ZN(Midori_rounds_n865)
         );
  AOI22_X1 Midori_rounds_U985 ( .A1(reset), .A2(Midori_add_Result_Start2[12]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[12]), .ZN(
        Midori_rounds_n1837) );
  XOR2_X1 Midori_rounds_U984 ( .A(Midori_rounds_SR_Inv_Result2[32]), .B(
        Midori_rounds_n1836), .Z(Midori_rounds_n1838) );
  OAI21_X1 Midori_rounds_U983 ( .B1(Midori_rounds_n1835), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1834), .ZN(
        Midori_rounds_sub_Sub_3_F_in2[0]) );
  AOI22_X1 Midori_rounds_U982 ( .A1(reset), .A2(Midori_add_Result_Start2[13]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result2[13]), .ZN(
        Midori_rounds_n1834) );
  XOR2_X1 Midori_rounds_U981 ( .A(Midori_rounds_SR_Inv_Result2[33]), .B(
        Midori_rounds_n1833), .Z(Midori_rounds_n1835) );
  OAI21_X1 Midori_rounds_U980 ( .B1(Midori_rounds_n1832), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1831), .ZN(Midori_rounds_n867)
         );
  AOI22_X1 Midori_rounds_U979 ( .A1(reset), .A2(Midori_add_Result_Start2[14]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result2[14]), .ZN(
        Midori_rounds_n1831) );
  XOR2_X1 Midori_rounds_U978 ( .A(Midori_rounds_SR_Inv_Result2[34]), .B(
        Midori_rounds_n1830), .Z(Midori_rounds_n1832) );
  OAI21_X1 Midori_rounds_U977 ( .B1(Midori_rounds_n1829), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1828), .ZN(
        Midori_rounds_sub_Sub_3_F_in2[2]) );
  AOI22_X1 Midori_rounds_U976 ( .A1(reset), .A2(Midori_add_Result_Start2[15]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result2[15]), .ZN(
        Midori_rounds_n1828) );
  XOR2_X1 Midori_rounds_U975 ( .A(Midori_rounds_SR_Inv_Result2[35]), .B(
        Midori_rounds_n1827), .Z(Midori_rounds_n1829) );
  OAI21_X1 Midori_rounds_U974 ( .B1(Midori_rounds_n1826), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1825), .ZN(Midori_rounds_n869)
         );
  AOI22_X1 Midori_rounds_U973 ( .A1(reset), .A2(Midori_add_Result_Start2[16]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[16]), .ZN(
        Midori_rounds_n1825) );
  XOR2_X1 Midori_rounds_U972 ( .A(Midori_rounds_SR_Inv_Result2[36]), .B(
        Midori_rounds_n1824), .Z(Midori_rounds_n1826) );
  OAI21_X1 Midori_rounds_U971 ( .B1(Midori_rounds_n1823), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1822), .ZN(
        Midori_rounds_sub_Sub_4_F_in2[0]) );
  AOI22_X1 Midori_rounds_U970 ( .A1(reset), .A2(Midori_add_Result_Start2[17]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[17]), .ZN(
        Midori_rounds_n1822) );
  XOR2_X1 Midori_rounds_U969 ( .A(Midori_rounds_SR_Inv_Result2[37]), .B(
        Midori_rounds_n1821), .Z(Midori_rounds_n1823) );
  OAI21_X1 Midori_rounds_U968 ( .B1(Midori_rounds_n1820), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1819), .ZN(Midori_rounds_n871)
         );
  AOI22_X1 Midori_rounds_U967 ( .A1(reset), .A2(Midori_add_Result_Start2[18]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[18]), .ZN(
        Midori_rounds_n1819) );
  XOR2_X1 Midori_rounds_U966 ( .A(Midori_rounds_SR_Inv_Result2[38]), .B(
        Midori_rounds_n1818), .Z(Midori_rounds_n1820) );
  OAI21_X1 Midori_rounds_U965 ( .B1(Midori_rounds_n1817), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1816), .ZN(
        Midori_rounds_sub_Sub_4_F_in2[2]) );
  AOI22_X1 Midori_rounds_U964 ( .A1(reset), .A2(Midori_add_Result_Start2[19]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result2[19]), .ZN(
        Midori_rounds_n1816) );
  XOR2_X1 Midori_rounds_U963 ( .A(Midori_rounds_SR_Inv_Result2[39]), .B(
        Midori_rounds_n1815), .Z(Midori_rounds_n1817) );
  OAI21_X1 Midori_rounds_U962 ( .B1(Midori_rounds_n1814), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1813), .ZN(Midori_rounds_n873)
         );
  AOI22_X1 Midori_rounds_U961 ( .A1(reset), .A2(Midori_add_Result_Start2[20]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[20]), .ZN(
        Midori_rounds_n1813) );
  XOR2_X1 Midori_rounds_U960 ( .A(Midori_rounds_SR_Inv_Result2[12]), .B(
        Midori_rounds_n1812), .Z(Midori_rounds_n1814) );
  OAI21_X1 Midori_rounds_U959 ( .B1(Midori_rounds_n1811), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1810), .ZN(
        Midori_rounds_sub_Sub_5_F_in2[0]) );
  AOI22_X1 Midori_rounds_U958 ( .A1(reset), .A2(Midori_add_Result_Start2[21]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[21]), .ZN(
        Midori_rounds_n1810) );
  XOR2_X1 Midori_rounds_U957 ( .A(Midori_rounds_SR_Inv_Result2[13]), .B(
        Midori_rounds_n1809), .Z(Midori_rounds_n1811) );
  OAI21_X1 Midori_rounds_U956 ( .B1(Midori_rounds_n1808), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1807), .ZN(Midori_rounds_n875)
         );
  AOI22_X1 Midori_rounds_U955 ( .A1(reset), .A2(Midori_add_Result_Start2[22]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[22]), .ZN(
        Midori_rounds_n1807) );
  XOR2_X1 Midori_rounds_U954 ( .A(Midori_rounds_SR_Inv_Result2[14]), .B(
        Midori_rounds_n1806), .Z(Midori_rounds_n1808) );
  OAI21_X1 Midori_rounds_U953 ( .B1(Midori_rounds_n1805), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1804), .ZN(
        Midori_rounds_sub_Sub_5_F_in2[2]) );
  AOI22_X1 Midori_rounds_U952 ( .A1(reset), .A2(Midori_add_Result_Start2[23]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[23]), .ZN(
        Midori_rounds_n1804) );
  XOR2_X1 Midori_rounds_U951 ( .A(Midori_rounds_SR_Inv_Result2[15]), .B(
        Midori_rounds_n1803), .Z(Midori_rounds_n1805) );
  OAI21_X1 Midori_rounds_U950 ( .B1(Midori_rounds_n1802), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1801), .ZN(Midori_rounds_n877)
         );
  AOI22_X1 Midori_rounds_U949 ( .A1(reset), .A2(Midori_add_Result_Start2[24]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[24]), .ZN(
        Midori_rounds_n1801) );
  XOR2_X1 Midori_rounds_U948 ( .A(Midori_rounds_SR_Inv_Result2[48]), .B(
        Midori_rounds_n1800), .Z(Midori_rounds_n1802) );
  OAI21_X1 Midori_rounds_U947 ( .B1(Midori_rounds_n1799), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1798), .ZN(
        Midori_rounds_sub_Sub_6_F_in2[0]) );
  AOI22_X1 Midori_rounds_U946 ( .A1(reset), .A2(Midori_add_Result_Start2[25]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[25]), .ZN(
        Midori_rounds_n1798) );
  XOR2_X1 Midori_rounds_U945 ( .A(Midori_rounds_SR_Inv_Result2[49]), .B(
        Midori_rounds_n1797), .Z(Midori_rounds_n1799) );
  OAI21_X1 Midori_rounds_U944 ( .B1(Midori_rounds_n1796), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1795), .ZN(Midori_rounds_n879)
         );
  AOI22_X1 Midori_rounds_U943 ( .A1(reset), .A2(Midori_add_Result_Start2[26]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result2[26]), .ZN(
        Midori_rounds_n1795) );
  XOR2_X1 Midori_rounds_U942 ( .A(Midori_rounds_SR_Inv_Result2[50]), .B(
        Midori_rounds_n1794), .Z(Midori_rounds_n1796) );
  OAI21_X1 Midori_rounds_U941 ( .B1(Midori_rounds_n1793), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1792), .ZN(
        Midori_rounds_sub_Sub_6_F_in2[2]) );
  AOI22_X1 Midori_rounds_U940 ( .A1(reset), .A2(Midori_add_Result_Start2[27]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result2[27]), .ZN(
        Midori_rounds_n1792) );
  XOR2_X1 Midori_rounds_U939 ( .A(Midori_rounds_SR_Inv_Result2[51]), .B(
        Midori_rounds_n1791), .Z(Midori_rounds_n1793) );
  OAI21_X1 Midori_rounds_U938 ( .B1(Midori_rounds_n1790), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1789), .ZN(Midori_rounds_n881)
         );
  AOI22_X1 Midori_rounds_U937 ( .A1(reset), .A2(Midori_add_Result_Start2[28]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[28]), .ZN(
        Midori_rounds_n1789) );
  XOR2_X1 Midori_rounds_U936 ( .A(Midori_rounds_SR_Inv_Result2[24]), .B(
        Midori_rounds_n1788), .Z(Midori_rounds_n1790) );
  OAI21_X1 Midori_rounds_U935 ( .B1(Midori_rounds_n1787), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1786), .ZN(
        Midori_rounds_sub_Sub_7_F_in2[0]) );
  AOI22_X1 Midori_rounds_U934 ( .A1(reset), .A2(Midori_add_Result_Start2[29]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[29]), .ZN(
        Midori_rounds_n1786) );
  XOR2_X1 Midori_rounds_U933 ( .A(Midori_rounds_SR_Inv_Result2[25]), .B(
        Midori_rounds_n1785), .Z(Midori_rounds_n1787) );
  OAI21_X1 Midori_rounds_U932 ( .B1(Midori_rounds_n1784), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1783), .ZN(Midori_rounds_n883)
         );
  AOI22_X1 Midori_rounds_U931 ( .A1(reset), .A2(Midori_add_Result_Start2[30]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[30]), .ZN(
        Midori_rounds_n1783) );
  XOR2_X1 Midori_rounds_U930 ( .A(Midori_rounds_SR_Inv_Result2[26]), .B(
        Midori_rounds_n1782), .Z(Midori_rounds_n1784) );
  OAI21_X1 Midori_rounds_U929 ( .B1(Midori_rounds_n1781), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1780), .ZN(
        Midori_rounds_sub_Sub_7_F_in2[2]) );
  AOI22_X1 Midori_rounds_U928 ( .A1(reset), .A2(Midori_add_Result_Start2[31]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[31]), .ZN(
        Midori_rounds_n1780) );
  XOR2_X1 Midori_rounds_U927 ( .A(Midori_rounds_SR_Inv_Result2[27]), .B(
        Midori_rounds_n1779), .Z(Midori_rounds_n1781) );
  OAI21_X1 Midori_rounds_U926 ( .B1(Midori_rounds_n1778), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1777), .ZN(Midori_rounds_n885)
         );
  AOI22_X1 Midori_rounds_U925 ( .A1(reset), .A2(Midori_add_Result_Start2[32]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[32]), .ZN(
        Midori_rounds_n1777) );
  XOR2_X1 Midori_rounds_U924 ( .A(Midori_rounds_SR_Inv_Result2[56]), .B(
        Midori_rounds_n1776), .Z(Midori_rounds_n1778) );
  OAI21_X1 Midori_rounds_U923 ( .B1(Midori_rounds_n1775), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1774), .ZN(
        Midori_rounds_sub_Sub_8_F_in2[0]) );
  AOI22_X1 Midori_rounds_U922 ( .A1(reset), .A2(Midori_add_Result_Start2[33]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[33]), .ZN(
        Midori_rounds_n1774) );
  XOR2_X1 Midori_rounds_U921 ( .A(Midori_rounds_SR_Inv_Result2[57]), .B(
        Midori_rounds_n1773), .Z(Midori_rounds_n1775) );
  OAI21_X1 Midori_rounds_U920 ( .B1(Midori_rounds_n1772), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1771), .ZN(Midori_rounds_n887)
         );
  AOI22_X1 Midori_rounds_U919 ( .A1(reset), .A2(Midori_add_Result_Start2[34]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[34]), .ZN(
        Midori_rounds_n1771) );
  XOR2_X1 Midori_rounds_U918 ( .A(Midori_rounds_SR_Inv_Result2[58]), .B(
        Midori_rounds_n1770), .Z(Midori_rounds_n1772) );
  OAI21_X1 Midori_rounds_U917 ( .B1(Midori_rounds_n1769), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1768), .ZN(
        Midori_rounds_sub_Sub_8_F_in2[2]) );
  AOI22_X1 Midori_rounds_U916 ( .A1(reset), .A2(Midori_add_Result_Start2[35]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[35]), .ZN(
        Midori_rounds_n1768) );
  XOR2_X1 Midori_rounds_U915 ( .A(Midori_rounds_SR_Inv_Result2[59]), .B(
        Midori_rounds_n1767), .Z(Midori_rounds_n1769) );
  OAI21_X1 Midori_rounds_U914 ( .B1(Midori_rounds_n1766), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1765), .ZN(Midori_rounds_n889)
         );
  AOI22_X1 Midori_rounds_U913 ( .A1(reset), .A2(Midori_add_Result_Start2[36]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[36]), .ZN(
        Midori_rounds_n1765) );
  XOR2_X1 Midori_rounds_U912 ( .A(Midori_rounds_SR_Inv_Result2[16]), .B(
        Midori_rounds_n1764), .Z(Midori_rounds_n1766) );
  OAI21_X1 Midori_rounds_U911 ( .B1(Midori_rounds_n1763), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1762), .ZN(
        Midori_rounds_sub_Sub_9_F_in2[0]) );
  AOI22_X1 Midori_rounds_U910 ( .A1(reset), .A2(Midori_add_Result_Start2[37]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[37]), .ZN(
        Midori_rounds_n1762) );
  XOR2_X1 Midori_rounds_U909 ( .A(Midori_rounds_SR_Inv_Result2[17]), .B(
        Midori_rounds_n1761), .Z(Midori_rounds_n1763) );
  OAI21_X1 Midori_rounds_U908 ( .B1(Midori_rounds_n1760), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1759), .ZN(Midori_rounds_n891)
         );
  AOI22_X1 Midori_rounds_U907 ( .A1(reset), .A2(Midori_add_Result_Start2[38]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[38]), .ZN(
        Midori_rounds_n1759) );
  XOR2_X1 Midori_rounds_U906 ( .A(Midori_rounds_SR_Inv_Result2[18]), .B(
        Midori_rounds_n1758), .Z(Midori_rounds_n1760) );
  OAI21_X1 Midori_rounds_U905 ( .B1(Midori_rounds_n1757), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1756), .ZN(
        Midori_rounds_sub_Sub_9_F_in2[2]) );
  AOI22_X1 Midori_rounds_U904 ( .A1(reset), .A2(Midori_add_Result_Start2[39]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[39]), .ZN(
        Midori_rounds_n1756) );
  XOR2_X1 Midori_rounds_U903 ( .A(Midori_rounds_SR_Inv_Result2[19]), .B(
        Midori_rounds_n1755), .Z(Midori_rounds_n1757) );
  OAI21_X1 Midori_rounds_U902 ( .B1(Midori_rounds_n1754), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1753), .ZN(Midori_rounds_n893)
         );
  AOI22_X1 Midori_rounds_U901 ( .A1(reset), .A2(Midori_add_Result_Start2[40]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[40]), .ZN(
        Midori_rounds_n1753) );
  XOR2_X1 Midori_rounds_U900 ( .A(Midori_rounds_SR_Inv_Result2[44]), .B(
        Midori_rounds_n1752), .Z(Midori_rounds_n1754) );
  OAI21_X1 Midori_rounds_U899 ( .B1(Midori_rounds_n1751), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1750), .ZN(
        Midori_rounds_sub_Sub_10_F_in2[0]) );
  AOI22_X1 Midori_rounds_U898 ( .A1(reset), .A2(Midori_add_Result_Start2[41]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[41]), .ZN(
        Midori_rounds_n1750) );
  XOR2_X1 Midori_rounds_U897 ( .A(Midori_rounds_SR_Inv_Result2[45]), .B(
        Midori_rounds_n1749), .Z(Midori_rounds_n1751) );
  OAI21_X1 Midori_rounds_U896 ( .B1(Midori_rounds_n1748), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1747), .ZN(Midori_rounds_n895)
         );
  AOI22_X1 Midori_rounds_U895 ( .A1(reset), .A2(Midori_add_Result_Start2[42]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[42]), .ZN(
        Midori_rounds_n1747) );
  XOR2_X1 Midori_rounds_U894 ( .A(Midori_rounds_SR_Inv_Result2[46]), .B(
        Midori_rounds_n1746), .Z(Midori_rounds_n1748) );
  OAI21_X1 Midori_rounds_U893 ( .B1(Midori_rounds_n1745), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1744), .ZN(
        Midori_rounds_sub_Sub_10_F_in2[2]) );
  AOI22_X1 Midori_rounds_U892 ( .A1(reset), .A2(Midori_add_Result_Start2[43]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[43]), .ZN(
        Midori_rounds_n1744) );
  XOR2_X1 Midori_rounds_U891 ( .A(Midori_rounds_SR_Inv_Result2[47]), .B(
        Midori_rounds_n1743), .Z(Midori_rounds_n1745) );
  OAI21_X1 Midori_rounds_U890 ( .B1(Midori_rounds_n1742), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1741), .ZN(Midori_rounds_n897)
         );
  AOI22_X1 Midori_rounds_U889 ( .A1(reset), .A2(Midori_add_Result_Start2[44]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[44]), .ZN(
        Midori_rounds_n1741) );
  XOR2_X1 Midori_rounds_U888 ( .A(Midori_rounds_SR_Inv_Result2[4]), .B(
        Midori_rounds_n1740), .Z(Midori_rounds_n1742) );
  OAI21_X1 Midori_rounds_U887 ( .B1(Midori_rounds_n1739), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1738), .ZN(
        Midori_rounds_sub_Sub_11_F_in2[0]) );
  AOI22_X1 Midori_rounds_U886 ( .A1(reset), .A2(Midori_add_Result_Start2[45]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[45]), .ZN(
        Midori_rounds_n1738) );
  XOR2_X1 Midori_rounds_U885 ( .A(Midori_rounds_SR_Inv_Result2[5]), .B(
        Midori_rounds_n1737), .Z(Midori_rounds_n1739) );
  OAI21_X1 Midori_rounds_U884 ( .B1(Midori_rounds_n1736), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1735), .ZN(Midori_rounds_n899)
         );
  AOI22_X1 Midori_rounds_U883 ( .A1(reset), .A2(Midori_add_Result_Start2[46]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[46]), .ZN(
        Midori_rounds_n1735) );
  XOR2_X1 Midori_rounds_U882 ( .A(Midori_rounds_SR_Inv_Result2[6]), .B(
        Midori_rounds_n1734), .Z(Midori_rounds_n1736) );
  OAI21_X1 Midori_rounds_U881 ( .B1(Midori_rounds_n1733), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1732), .ZN(
        Midori_rounds_sub_Sub_11_F_in2[2]) );
  AOI22_X1 Midori_rounds_U880 ( .A1(reset), .A2(Midori_add_Result_Start2[47]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[47]), .ZN(
        Midori_rounds_n1732) );
  XOR2_X1 Midori_rounds_U879 ( .A(Midori_rounds_SR_Inv_Result2[7]), .B(
        Midori_rounds_n1731), .Z(Midori_rounds_n1733) );
  OAI21_X1 Midori_rounds_U878 ( .B1(Midori_rounds_n1730), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1729), .ZN(Midori_rounds_n901)
         );
  AOI22_X1 Midori_rounds_U877 ( .A1(reset), .A2(Midori_add_Result_Start2[48]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[48]), .ZN(
        Midori_rounds_n1729) );
  XOR2_X1 Midori_rounds_U876 ( .A(Midori_rounds_SR_Inv_Result2[0]), .B(
        Midori_rounds_n1728), .Z(Midori_rounds_n1730) );
  OAI21_X1 Midori_rounds_U875 ( .B1(Midori_rounds_n1727), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1726), .ZN(
        Midori_rounds_sub_Sub_12_F_in2[0]) );
  AOI22_X1 Midori_rounds_U874 ( .A1(reset), .A2(Midori_add_Result_Start2[49]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[49]), .ZN(
        Midori_rounds_n1726) );
  XOR2_X1 Midori_rounds_U873 ( .A(Midori_rounds_SR_Inv_Result2[1]), .B(
        Midori_rounds_n1725), .Z(Midori_rounds_n1727) );
  OAI21_X1 Midori_rounds_U872 ( .B1(Midori_rounds_n1724), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1723), .ZN(Midori_rounds_n903)
         );
  AOI22_X1 Midori_rounds_U871 ( .A1(reset), .A2(Midori_add_Result_Start2[50]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[50]), .ZN(
        Midori_rounds_n1723) );
  XOR2_X1 Midori_rounds_U870 ( .A(Midori_rounds_SR_Inv_Result2[2]), .B(
        Midori_rounds_n1722), .Z(Midori_rounds_n1724) );
  OAI21_X1 Midori_rounds_U869 ( .B1(Midori_rounds_n1721), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1720), .ZN(
        Midori_rounds_sub_Sub_12_F_in2[2]) );
  AOI22_X1 Midori_rounds_U868 ( .A1(reset), .A2(Midori_add_Result_Start2[51]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[51]), .ZN(
        Midori_rounds_n1720) );
  XOR2_X1 Midori_rounds_U867 ( .A(Midori_rounds_SR_Inv_Result2[3]), .B(
        Midori_rounds_n1719), .Z(Midori_rounds_n1721) );
  OAI21_X1 Midori_rounds_U866 ( .B1(Midori_rounds_n1718), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1717), .ZN(Midori_rounds_n905)
         );
  AOI22_X1 Midori_rounds_U865 ( .A1(reset), .A2(Midori_add_Result_Start2[52]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[52]), .ZN(
        Midori_rounds_n1717) );
  XOR2_X1 Midori_rounds_U864 ( .A(Midori_rounds_SR_Inv_Result2[40]), .B(
        Midori_rounds_n1716), .Z(Midori_rounds_n1718) );
  OAI21_X1 Midori_rounds_U863 ( .B1(Midori_rounds_n1715), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1714), .ZN(
        Midori_rounds_sub_Sub_13_F_in2[0]) );
  AOI22_X1 Midori_rounds_U862 ( .A1(reset), .A2(Midori_add_Result_Start2[53]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[53]), .ZN(
        Midori_rounds_n1714) );
  XOR2_X1 Midori_rounds_U861 ( .A(Midori_rounds_SR_Inv_Result2[41]), .B(
        Midori_rounds_n1713), .Z(Midori_rounds_n1715) );
  OAI21_X1 Midori_rounds_U860 ( .B1(Midori_rounds_n1712), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1711), .ZN(Midori_rounds_n907)
         );
  AOI22_X1 Midori_rounds_U859 ( .A1(reset), .A2(Midori_add_Result_Start2[54]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[54]), .ZN(
        Midori_rounds_n1711) );
  XOR2_X1 Midori_rounds_U858 ( .A(Midori_rounds_SR_Inv_Result2[42]), .B(
        Midori_rounds_n1710), .Z(Midori_rounds_n1712) );
  OAI21_X1 Midori_rounds_U857 ( .B1(Midori_rounds_n1709), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1708), .ZN(
        Midori_rounds_sub_Sub_13_F_in2[2]) );
  AOI22_X1 Midori_rounds_U856 ( .A1(reset), .A2(Midori_add_Result_Start2[55]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[55]), .ZN(
        Midori_rounds_n1708) );
  XOR2_X1 Midori_rounds_U855 ( .A(Midori_rounds_SR_Inv_Result2[43]), .B(
        Midori_rounds_n1707), .Z(Midori_rounds_n1709) );
  OAI21_X1 Midori_rounds_U854 ( .B1(Midori_rounds_n1706), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1705), .ZN(Midori_rounds_n909)
         );
  AOI22_X1 Midori_rounds_U853 ( .A1(reset), .A2(Midori_add_Result_Start2[56]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[56]), .ZN(
        Midori_rounds_n1705) );
  XOR2_X1 Midori_rounds_U852 ( .A(Midori_rounds_SR_Inv_Result2[20]), .B(
        Midori_rounds_n1704), .Z(Midori_rounds_n1706) );
  OAI21_X1 Midori_rounds_U851 ( .B1(Midori_rounds_n1703), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1702), .ZN(
        Midori_rounds_sub_Sub_14_F_in2[0]) );
  AOI22_X1 Midori_rounds_U850 ( .A1(reset), .A2(Midori_add_Result_Start2[57]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[57]), .ZN(
        Midori_rounds_n1702) );
  XOR2_X1 Midori_rounds_U849 ( .A(Midori_rounds_SR_Inv_Result2[21]), .B(
        Midori_rounds_n1701), .Z(Midori_rounds_n1703) );
  OAI21_X1 Midori_rounds_U848 ( .B1(Midori_rounds_n1700), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1699), .ZN(Midori_rounds_n911)
         );
  AOI22_X1 Midori_rounds_U847 ( .A1(reset), .A2(Midori_add_Result_Start2[58]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[58]), .ZN(
        Midori_rounds_n1699) );
  XOR2_X1 Midori_rounds_U846 ( .A(Midori_rounds_SR_Inv_Result2[22]), .B(
        Midori_rounds_n1698), .Z(Midori_rounds_n1700) );
  OAI21_X1 Midori_rounds_U845 ( .B1(Midori_rounds_n1697), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1696), .ZN(
        Midori_rounds_sub_Sub_14_F_in2[2]) );
  AOI22_X1 Midori_rounds_U844 ( .A1(reset), .A2(Midori_add_Result_Start2[59]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[59]), .ZN(
        Midori_rounds_n1696) );
  XOR2_X1 Midori_rounds_U843 ( .A(Midori_rounds_SR_Inv_Result2[23]), .B(
        Midori_rounds_n1695), .Z(Midori_rounds_n1697) );
  OAI21_X1 Midori_rounds_U842 ( .B1(Midori_rounds_n1694), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1693), .ZN(Midori_rounds_n913)
         );
  AOI22_X1 Midori_rounds_U841 ( .A1(reset), .A2(Midori_add_Result_Start2[60]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[60]), .ZN(
        Midori_rounds_n1693) );
  XOR2_X1 Midori_rounds_U840 ( .A(Midori_rounds_SR_Inv_Result2[60]), .B(
        Midori_rounds_n1692), .Z(Midori_rounds_n1694) );
  OAI21_X1 Midori_rounds_U839 ( .B1(Midori_rounds_n1691), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1690), .ZN(
        Midori_rounds_sub_Sub_15_F_in2[0]) );
  AOI22_X1 Midori_rounds_U838 ( .A1(reset), .A2(Midori_add_Result_Start2[61]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[61]), .ZN(
        Midori_rounds_n1690) );
  XOR2_X1 Midori_rounds_U837 ( .A(Midori_rounds_SR_Inv_Result2[61]), .B(
        Midori_rounds_n1689), .Z(Midori_rounds_n1691) );
  OAI21_X1 Midori_rounds_U836 ( .B1(Midori_rounds_n1688), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1687), .ZN(Midori_rounds_n915)
         );
  AOI22_X1 Midori_rounds_U835 ( .A1(reset), .A2(Midori_add_Result_Start2[62]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[62]), .ZN(
        Midori_rounds_n1687) );
  XOR2_X1 Midori_rounds_U834 ( .A(Midori_rounds_SR_Inv_Result2[62]), .B(
        Midori_rounds_n1686), .Z(Midori_rounds_n1688) );
  OAI21_X1 Midori_rounds_U833 ( .B1(Midori_rounds_n1685), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1684), .ZN(
        Midori_rounds_sub_Sub_15_F_in2[2]) );
  AOI22_X1 Midori_rounds_U832 ( .A1(reset), .A2(Midori_add_Result_Start2[63]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[63]), .ZN(
        Midori_rounds_n1684) );
  XOR2_X1 Midori_rounds_U831 ( .A(Midori_rounds_SR_Inv_Result2[63]), .B(
        Midori_rounds_n1683), .Z(Midori_rounds_n1685) );
  OAI21_X1 Midori_rounds_U830 ( .B1(Midori_rounds_n1682), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1681), .ZN(Midori_rounds_n917)
         );
  AOI22_X1 Midori_rounds_U829 ( .A1(reset), .A2(Midori_add_Result_Start3[0]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[0]), .ZN(
        Midori_rounds_n1681) );
  XOR2_X1 Midori_rounds_U828 ( .A(Midori_rounds_SR_Inv_Result3[28]), .B(
        Midori_rounds_n1680), .Z(Midori_rounds_n1682) );
  OAI21_X1 Midori_rounds_U827 ( .B1(Midori_rounds_n1679), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1678), .ZN(
        Midori_rounds_sub_Sub_0_F_in3[0]) );
  AOI22_X1 Midori_rounds_U826 ( .A1(reset), .A2(Midori_add_Result_Start3[1]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[1]), .ZN(
        Midori_rounds_n1678) );
  XOR2_X1 Midori_rounds_U825 ( .A(Midori_rounds_SR_Inv_Result3[29]), .B(
        Midori_rounds_n1677), .Z(Midori_rounds_n1679) );
  OAI21_X1 Midori_rounds_U824 ( .B1(Midori_rounds_n1676), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1675), .ZN(Midori_rounds_n919)
         );
  AOI22_X1 Midori_rounds_U823 ( .A1(reset), .A2(Midori_add_Result_Start3[2]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[2]), .ZN(
        Midori_rounds_n1675) );
  XOR2_X1 Midori_rounds_U822 ( .A(Midori_rounds_SR_Inv_Result3[30]), .B(
        Midori_rounds_n1674), .Z(Midori_rounds_n1676) );
  OAI21_X1 Midori_rounds_U821 ( .B1(Midori_rounds_n1673), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1672), .ZN(
        Midori_rounds_sub_Sub_0_F_in3[2]) );
  AOI22_X1 Midori_rounds_U820 ( .A1(reset), .A2(Midori_add_Result_Start3[3]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[3]), .ZN(
        Midori_rounds_n1672) );
  XOR2_X1 Midori_rounds_U819 ( .A(Midori_rounds_SR_Inv_Result3[31]), .B(
        Midori_rounds_n1671), .Z(Midori_rounds_n1673) );
  OAI21_X1 Midori_rounds_U818 ( .B1(Midori_rounds_n1670), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1669), .ZN(Midori_rounds_n921)
         );
  AOI22_X1 Midori_rounds_U817 ( .A1(reset), .A2(Midori_add_Result_Start3[4]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[4]), .ZN(
        Midori_rounds_n1669) );
  XOR2_X1 Midori_rounds_U816 ( .A(Midori_rounds_SR_Inv_Result3[52]), .B(
        Midori_rounds_n1668), .Z(Midori_rounds_n1670) );
  OAI21_X1 Midori_rounds_U815 ( .B1(Midori_rounds_n1667), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1666), .ZN(
        Midori_rounds_sub_Sub_1_F_in3[0]) );
  AOI22_X1 Midori_rounds_U814 ( .A1(reset), .A2(Midori_add_Result_Start3[5]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[5]), .ZN(
        Midori_rounds_n1666) );
  XOR2_X1 Midori_rounds_U813 ( .A(Midori_rounds_SR_Inv_Result3[53]), .B(
        Midori_rounds_n1665), .Z(Midori_rounds_n1667) );
  OAI21_X1 Midori_rounds_U812 ( .B1(Midori_rounds_n1664), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1663), .ZN(Midori_rounds_n923)
         );
  AOI22_X1 Midori_rounds_U811 ( .A1(reset), .A2(Midori_add_Result_Start3[6]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[6]), .ZN(
        Midori_rounds_n1663) );
  XOR2_X1 Midori_rounds_U810 ( .A(Midori_rounds_SR_Inv_Result3[54]), .B(
        Midori_rounds_n1662), .Z(Midori_rounds_n1664) );
  OAI21_X1 Midori_rounds_U809 ( .B1(Midori_rounds_n1661), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1660), .ZN(
        Midori_rounds_sub_Sub_1_F_in3[2]) );
  AOI22_X1 Midori_rounds_U808 ( .A1(reset), .A2(Midori_add_Result_Start3[7]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[7]), .ZN(
        Midori_rounds_n1660) );
  XOR2_X1 Midori_rounds_U807 ( .A(Midori_rounds_SR_Inv_Result3[55]), .B(
        Midori_rounds_n1659), .Z(Midori_rounds_n1661) );
  OAI21_X1 Midori_rounds_U806 ( .B1(Midori_rounds_n1658), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1657), .ZN(Midori_rounds_n925)
         );
  AOI22_X1 Midori_rounds_U805 ( .A1(reset), .A2(Midori_add_Result_Start3[8]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[8]), .ZN(
        Midori_rounds_n1657) );
  XOR2_X1 Midori_rounds_U804 ( .A(Midori_rounds_SR_Inv_Result3[8]), .B(
        Midori_rounds_n1656), .Z(Midori_rounds_n1658) );
  OAI21_X1 Midori_rounds_U803 ( .B1(Midori_rounds_n1655), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1654), .ZN(
        Midori_rounds_sub_Sub_2_F_in3[0]) );
  AOI22_X1 Midori_rounds_U802 ( .A1(reset), .A2(Midori_add_Result_Start3[9]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[9]), .ZN(
        Midori_rounds_n1654) );
  XOR2_X1 Midori_rounds_U801 ( .A(Midori_rounds_SR_Inv_Result3[9]), .B(
        Midori_rounds_n1653), .Z(Midori_rounds_n1655) );
  OAI21_X1 Midori_rounds_U800 ( .B1(Midori_rounds_n1652), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1651), .ZN(Midori_rounds_n927)
         );
  AOI22_X1 Midori_rounds_U799 ( .A1(reset), .A2(Midori_add_Result_Start3[10]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[10]), .ZN(
        Midori_rounds_n1651) );
  XOR2_X1 Midori_rounds_U798 ( .A(Midori_rounds_SR_Inv_Result3[10]), .B(
        Midori_rounds_n1650), .Z(Midori_rounds_n1652) );
  OAI21_X1 Midori_rounds_U797 ( .B1(Midori_rounds_n1649), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1648), .ZN(
        Midori_rounds_sub_Sub_2_F_in3[2]) );
  AOI22_X1 Midori_rounds_U796 ( .A1(reset), .A2(Midori_add_Result_Start3[11]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[11]), .ZN(
        Midori_rounds_n1648) );
  XOR2_X1 Midori_rounds_U795 ( .A(Midori_rounds_SR_Inv_Result3[11]), .B(
        Midori_rounds_n1647), .Z(Midori_rounds_n1649) );
  OAI21_X1 Midori_rounds_U794 ( .B1(Midori_rounds_n1646), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1645), .ZN(Midori_rounds_n929)
         );
  AOI22_X1 Midori_rounds_U793 ( .A1(reset), .A2(Midori_add_Result_Start3[12]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[12]), .ZN(
        Midori_rounds_n1645) );
  XOR2_X1 Midori_rounds_U792 ( .A(Midori_rounds_SR_Inv_Result3[32]), .B(
        Midori_rounds_n1644), .Z(Midori_rounds_n1646) );
  OAI21_X1 Midori_rounds_U791 ( .B1(Midori_rounds_n1643), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1642), .ZN(
        Midori_rounds_sub_Sub_3_F_in3[0]) );
  AOI22_X1 Midori_rounds_U790 ( .A1(reset), .A2(Midori_add_Result_Start3[13]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[13]), .ZN(
        Midori_rounds_n1642) );
  XOR2_X1 Midori_rounds_U789 ( .A(Midori_rounds_SR_Inv_Result3[33]), .B(
        Midori_rounds_n1641), .Z(Midori_rounds_n1643) );
  OAI21_X1 Midori_rounds_U788 ( .B1(Midori_rounds_n1640), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1639), .ZN(Midori_rounds_n931)
         );
  AOI22_X1 Midori_rounds_U787 ( .A1(reset), .A2(Midori_add_Result_Start3[14]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[14]), .ZN(
        Midori_rounds_n1639) );
  XOR2_X1 Midori_rounds_U786 ( .A(Midori_rounds_SR_Inv_Result3[34]), .B(
        Midori_rounds_n1638), .Z(Midori_rounds_n1640) );
  OAI21_X1 Midori_rounds_U785 ( .B1(Midori_rounds_n1637), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1636), .ZN(
        Midori_rounds_sub_Sub_3_F_in3[2]) );
  AOI22_X1 Midori_rounds_U784 ( .A1(reset), .A2(Midori_add_Result_Start3[15]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[15]), .ZN(
        Midori_rounds_n1636) );
  XOR2_X1 Midori_rounds_U783 ( .A(Midori_rounds_SR_Inv_Result3[35]), .B(
        Midori_rounds_n1635), .Z(Midori_rounds_n1637) );
  OAI21_X1 Midori_rounds_U782 ( .B1(Midori_rounds_n1634), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1633), .ZN(Midori_rounds_n933)
         );
  AOI22_X1 Midori_rounds_U781 ( .A1(reset), .A2(Midori_add_Result_Start3[16]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[16]), .ZN(
        Midori_rounds_n1633) );
  XOR2_X1 Midori_rounds_U780 ( .A(Midori_rounds_SR_Inv_Result3[36]), .B(
        Midori_rounds_n1632), .Z(Midori_rounds_n1634) );
  OAI21_X1 Midori_rounds_U779 ( .B1(Midori_rounds_n1631), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1630), .ZN(
        Midori_rounds_sub_Sub_4_F_in3[0]) );
  AOI22_X1 Midori_rounds_U778 ( .A1(reset), .A2(Midori_add_Result_Start3[17]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[17]), .ZN(
        Midori_rounds_n1630) );
  XOR2_X1 Midori_rounds_U777 ( .A(Midori_rounds_SR_Inv_Result3[37]), .B(
        Midori_rounds_n1629), .Z(Midori_rounds_n1631) );
  OAI21_X1 Midori_rounds_U776 ( .B1(Midori_rounds_n1628), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1627), .ZN(Midori_rounds_n935)
         );
  AOI22_X1 Midori_rounds_U775 ( .A1(reset), .A2(Midori_add_Result_Start3[18]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[18]), .ZN(
        Midori_rounds_n1627) );
  XOR2_X1 Midori_rounds_U774 ( .A(Midori_rounds_SR_Inv_Result3[38]), .B(
        Midori_rounds_n1626), .Z(Midori_rounds_n1628) );
  OAI21_X1 Midori_rounds_U773 ( .B1(Midori_rounds_n1625), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1624), .ZN(
        Midori_rounds_sub_Sub_4_F_in3[2]) );
  AOI22_X1 Midori_rounds_U772 ( .A1(reset), .A2(Midori_add_Result_Start3[19]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[19]), .ZN(
        Midori_rounds_n1624) );
  XOR2_X1 Midori_rounds_U771 ( .A(Midori_rounds_SR_Inv_Result3[39]), .B(
        Midori_rounds_n1623), .Z(Midori_rounds_n1625) );
  OAI21_X1 Midori_rounds_U770 ( .B1(Midori_rounds_n1622), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1621), .ZN(Midori_rounds_n937)
         );
  AOI22_X1 Midori_rounds_U769 ( .A1(reset), .A2(Midori_add_Result_Start3[20]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[20]), .ZN(
        Midori_rounds_n1621) );
  XOR2_X1 Midori_rounds_U768 ( .A(Midori_rounds_SR_Inv_Result3[12]), .B(
        Midori_rounds_n1620), .Z(Midori_rounds_n1622) );
  OAI21_X1 Midori_rounds_U767 ( .B1(Midori_rounds_n1619), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1618), .ZN(
        Midori_rounds_sub_Sub_5_F_in3[0]) );
  AOI22_X1 Midori_rounds_U766 ( .A1(reset), .A2(Midori_add_Result_Start3[21]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[21]), .ZN(
        Midori_rounds_n1618) );
  XOR2_X1 Midori_rounds_U765 ( .A(Midori_rounds_SR_Inv_Result3[13]), .B(
        Midori_rounds_n1617), .Z(Midori_rounds_n1619) );
  OAI21_X1 Midori_rounds_U764 ( .B1(Midori_rounds_n1616), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1615), .ZN(Midori_rounds_n939)
         );
  AOI22_X1 Midori_rounds_U763 ( .A1(reset), .A2(Midori_add_Result_Start3[22]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[22]), .ZN(
        Midori_rounds_n1615) );
  XOR2_X1 Midori_rounds_U762 ( .A(Midori_rounds_SR_Inv_Result3[14]), .B(
        Midori_rounds_n1614), .Z(Midori_rounds_n1616) );
  OAI21_X1 Midori_rounds_U761 ( .B1(Midori_rounds_n1613), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1612), .ZN(
        Midori_rounds_sub_Sub_5_F_in3[2]) );
  AOI22_X1 Midori_rounds_U760 ( .A1(reset), .A2(Midori_add_Result_Start3[23]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[23]), .ZN(
        Midori_rounds_n1612) );
  XOR2_X1 Midori_rounds_U759 ( .A(Midori_rounds_SR_Inv_Result3[15]), .B(
        Midori_rounds_n1611), .Z(Midori_rounds_n1613) );
  OAI21_X1 Midori_rounds_U758 ( .B1(Midori_rounds_n1610), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1609), .ZN(Midori_rounds_n941)
         );
  AOI22_X1 Midori_rounds_U757 ( .A1(reset), .A2(Midori_add_Result_Start3[24]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[24]), .ZN(
        Midori_rounds_n1609) );
  XOR2_X1 Midori_rounds_U756 ( .A(Midori_rounds_SR_Inv_Result3[48]), .B(
        Midori_rounds_n1608), .Z(Midori_rounds_n1610) );
  OAI21_X1 Midori_rounds_U755 ( .B1(Midori_rounds_n1607), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1606), .ZN(
        Midori_rounds_sub_Sub_6_F_in3[0]) );
  AOI22_X1 Midori_rounds_U754 ( .A1(reset), .A2(Midori_add_Result_Start3[25]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[25]), .ZN(
        Midori_rounds_n1606) );
  XOR2_X1 Midori_rounds_U753 ( .A(Midori_rounds_SR_Inv_Result3[49]), .B(
        Midori_rounds_n1605), .Z(Midori_rounds_n1607) );
  OAI21_X1 Midori_rounds_U752 ( .B1(Midori_rounds_n1604), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1603), .ZN(Midori_rounds_n943)
         );
  AOI22_X1 Midori_rounds_U751 ( .A1(reset), .A2(Midori_add_Result_Start3[26]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[26]), .ZN(
        Midori_rounds_n1603) );
  XOR2_X1 Midori_rounds_U750 ( .A(Midori_rounds_SR_Inv_Result3[50]), .B(
        Midori_rounds_n1602), .Z(Midori_rounds_n1604) );
  OAI21_X1 Midori_rounds_U749 ( .B1(Midori_rounds_n1601), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1600), .ZN(
        Midori_rounds_sub_Sub_6_F_in3[2]) );
  AOI22_X1 Midori_rounds_U748 ( .A1(reset), .A2(Midori_add_Result_Start3[27]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[27]), .ZN(
        Midori_rounds_n1600) );
  XOR2_X1 Midori_rounds_U747 ( .A(Midori_rounds_SR_Inv_Result3[51]), .B(
        Midori_rounds_n1599), .Z(Midori_rounds_n1601) );
  OAI21_X1 Midori_rounds_U746 ( .B1(Midori_rounds_n1598), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1597), .ZN(Midori_rounds_n945)
         );
  AOI22_X1 Midori_rounds_U745 ( .A1(reset), .A2(Midori_add_Result_Start3[28]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[28]), .ZN(
        Midori_rounds_n1597) );
  XOR2_X1 Midori_rounds_U744 ( .A(Midori_rounds_SR_Inv_Result3[24]), .B(
        Midori_rounds_n1596), .Z(Midori_rounds_n1598) );
  OAI21_X1 Midori_rounds_U743 ( .B1(Midori_rounds_n1595), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1594), .ZN(
        Midori_rounds_sub_Sub_7_F_in3[0]) );
  AOI22_X1 Midori_rounds_U742 ( .A1(reset), .A2(Midori_add_Result_Start3[29]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[29]), .ZN(
        Midori_rounds_n1594) );
  XOR2_X1 Midori_rounds_U741 ( .A(Midori_rounds_SR_Inv_Result3[25]), .B(
        Midori_rounds_n1593), .Z(Midori_rounds_n1595) );
  OAI21_X1 Midori_rounds_U740 ( .B1(Midori_rounds_n1592), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1591), .ZN(Midori_rounds_n947)
         );
  AOI22_X1 Midori_rounds_U739 ( .A1(reset), .A2(Midori_add_Result_Start3[30]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[30]), .ZN(
        Midori_rounds_n1591) );
  XOR2_X1 Midori_rounds_U738 ( .A(Midori_rounds_SR_Inv_Result3[26]), .B(
        Midori_rounds_n1590), .Z(Midori_rounds_n1592) );
  OAI21_X1 Midori_rounds_U737 ( .B1(Midori_rounds_n1589), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1588), .ZN(
        Midori_rounds_sub_Sub_7_F_in3[2]) );
  AOI22_X1 Midori_rounds_U736 ( .A1(reset), .A2(Midori_add_Result_Start3[31]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[31]), .ZN(
        Midori_rounds_n1588) );
  XOR2_X1 Midori_rounds_U735 ( .A(Midori_rounds_SR_Inv_Result3[27]), .B(
        Midori_rounds_n1587), .Z(Midori_rounds_n1589) );
  OAI21_X1 Midori_rounds_U734 ( .B1(Midori_rounds_n1586), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1585), .ZN(Midori_rounds_n949)
         );
  AOI22_X1 Midori_rounds_U733 ( .A1(reset), .A2(Midori_add_Result_Start3[32]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[32]), .ZN(
        Midori_rounds_n1585) );
  XOR2_X1 Midori_rounds_U732 ( .A(Midori_rounds_SR_Inv_Result3[56]), .B(
        Midori_rounds_n1584), .Z(Midori_rounds_n1586) );
  OAI21_X1 Midori_rounds_U731 ( .B1(Midori_rounds_n1583), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1582), .ZN(
        Midori_rounds_sub_Sub_8_F_in3[0]) );
  AOI22_X1 Midori_rounds_U730 ( .A1(reset), .A2(Midori_add_Result_Start3[33]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[33]), .ZN(
        Midori_rounds_n1582) );
  XOR2_X1 Midori_rounds_U729 ( .A(Midori_rounds_SR_Inv_Result3[57]), .B(
        Midori_rounds_n1581), .Z(Midori_rounds_n1583) );
  OAI21_X1 Midori_rounds_U728 ( .B1(Midori_rounds_n1580), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1579), .ZN(Midori_rounds_n951)
         );
  AOI22_X1 Midori_rounds_U727 ( .A1(reset), .A2(Midori_add_Result_Start3[34]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[34]), .ZN(
        Midori_rounds_n1579) );
  XOR2_X1 Midori_rounds_U726 ( .A(Midori_rounds_SR_Inv_Result3[58]), .B(
        Midori_rounds_n1578), .Z(Midori_rounds_n1580) );
  OAI21_X1 Midori_rounds_U725 ( .B1(Midori_rounds_n1577), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1576), .ZN(
        Midori_rounds_sub_Sub_8_F_in3[2]) );
  AOI22_X1 Midori_rounds_U724 ( .A1(reset), .A2(Midori_add_Result_Start3[35]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[35]), .ZN(
        Midori_rounds_n1576) );
  XOR2_X1 Midori_rounds_U723 ( .A(Midori_rounds_SR_Inv_Result3[59]), .B(
        Midori_rounds_n1575), .Z(Midori_rounds_n1577) );
  OAI21_X1 Midori_rounds_U722 ( .B1(Midori_rounds_n1574), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1573), .ZN(Midori_rounds_n953)
         );
  AOI22_X1 Midori_rounds_U721 ( .A1(reset), .A2(Midori_add_Result_Start3[36]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[36]), .ZN(
        Midori_rounds_n1573) );
  XOR2_X1 Midori_rounds_U720 ( .A(Midori_rounds_SR_Inv_Result3[16]), .B(
        Midori_rounds_n1572), .Z(Midori_rounds_n1574) );
  OAI21_X1 Midori_rounds_U719 ( .B1(Midori_rounds_n1571), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1570), .ZN(
        Midori_rounds_sub_Sub_9_F_in3[0]) );
  AOI22_X1 Midori_rounds_U718 ( .A1(reset), .A2(Midori_add_Result_Start3[37]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[37]), .ZN(
        Midori_rounds_n1570) );
  XOR2_X1 Midori_rounds_U717 ( .A(Midori_rounds_SR_Inv_Result3[17]), .B(
        Midori_rounds_n1569), .Z(Midori_rounds_n1571) );
  OAI21_X1 Midori_rounds_U716 ( .B1(Midori_rounds_n1568), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1567), .ZN(Midori_rounds_n955)
         );
  AOI22_X1 Midori_rounds_U715 ( .A1(reset), .A2(Midori_add_Result_Start3[38]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[38]), .ZN(
        Midori_rounds_n1567) );
  XOR2_X1 Midori_rounds_U714 ( .A(Midori_rounds_SR_Inv_Result3[18]), .B(
        Midori_rounds_n1566), .Z(Midori_rounds_n1568) );
  OAI21_X1 Midori_rounds_U713 ( .B1(Midori_rounds_n1565), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1564), .ZN(
        Midori_rounds_sub_Sub_9_F_in3[2]) );
  AOI22_X1 Midori_rounds_U712 ( .A1(reset), .A2(Midori_add_Result_Start3[39]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[39]), .ZN(
        Midori_rounds_n1564) );
  XOR2_X1 Midori_rounds_U711 ( .A(Midori_rounds_SR_Inv_Result3[19]), .B(
        Midori_rounds_n1563), .Z(Midori_rounds_n1565) );
  OAI21_X1 Midori_rounds_U710 ( .B1(Midori_rounds_n1562), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1561), .ZN(Midori_rounds_n957)
         );
  AOI22_X1 Midori_rounds_U709 ( .A1(reset), .A2(Midori_add_Result_Start3[40]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[40]), .ZN(
        Midori_rounds_n1561) );
  XOR2_X1 Midori_rounds_U708 ( .A(Midori_rounds_SR_Inv_Result3[44]), .B(
        Midori_rounds_n1560), .Z(Midori_rounds_n1562) );
  OAI21_X1 Midori_rounds_U707 ( .B1(Midori_rounds_n1559), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1558), .ZN(
        Midori_rounds_sub_Sub_10_F_in3[0]) );
  AOI22_X1 Midori_rounds_U706 ( .A1(reset), .A2(Midori_add_Result_Start3[41]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[41]), .ZN(
        Midori_rounds_n1558) );
  XOR2_X1 Midori_rounds_U705 ( .A(Midori_rounds_SR_Inv_Result3[45]), .B(
        Midori_rounds_n1557), .Z(Midori_rounds_n1559) );
  OAI21_X1 Midori_rounds_U704 ( .B1(Midori_rounds_n1556), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1555), .ZN(Midori_rounds_n959)
         );
  AOI22_X1 Midori_rounds_U703 ( .A1(reset), .A2(Midori_add_Result_Start3[42]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[42]), .ZN(
        Midori_rounds_n1555) );
  XOR2_X1 Midori_rounds_U702 ( .A(Midori_rounds_SR_Inv_Result3[46]), .B(
        Midori_rounds_n1554), .Z(Midori_rounds_n1556) );
  OAI21_X1 Midori_rounds_U701 ( .B1(Midori_rounds_n1553), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1552), .ZN(
        Midori_rounds_sub_Sub_10_F_in3[2]) );
  AOI22_X1 Midori_rounds_U700 ( .A1(reset), .A2(Midori_add_Result_Start3[43]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[43]), .ZN(
        Midori_rounds_n1552) );
  XOR2_X1 Midori_rounds_U699 ( .A(Midori_rounds_SR_Inv_Result3[47]), .B(
        Midori_rounds_n1551), .Z(Midori_rounds_n1553) );
  OAI21_X1 Midori_rounds_U698 ( .B1(Midori_rounds_n1550), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1549), .ZN(Midori_rounds_n961)
         );
  AOI22_X1 Midori_rounds_U697 ( .A1(reset), .A2(Midori_add_Result_Start3[44]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[44]), .ZN(
        Midori_rounds_n1549) );
  XOR2_X1 Midori_rounds_U696 ( .A(Midori_rounds_SR_Inv_Result3[4]), .B(
        Midori_rounds_n1548), .Z(Midori_rounds_n1550) );
  OAI21_X1 Midori_rounds_U695 ( .B1(Midori_rounds_n1547), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1546), .ZN(
        Midori_rounds_sub_Sub_11_F_in3[0]) );
  AOI22_X1 Midori_rounds_U694 ( .A1(reset), .A2(Midori_add_Result_Start3[45]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[45]), .ZN(
        Midori_rounds_n1546) );
  XOR2_X1 Midori_rounds_U693 ( .A(Midori_rounds_SR_Inv_Result3[5]), .B(
        Midori_rounds_n1545), .Z(Midori_rounds_n1547) );
  OAI21_X1 Midori_rounds_U692 ( .B1(Midori_rounds_n1544), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1543), .ZN(Midori_rounds_n963)
         );
  AOI22_X1 Midori_rounds_U691 ( .A1(reset), .A2(Midori_add_Result_Start3[46]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[46]), .ZN(
        Midori_rounds_n1543) );
  XOR2_X1 Midori_rounds_U690 ( .A(Midori_rounds_SR_Inv_Result3[6]), .B(
        Midori_rounds_n1542), .Z(Midori_rounds_n1544) );
  OAI21_X1 Midori_rounds_U689 ( .B1(Midori_rounds_n1541), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1540), .ZN(
        Midori_rounds_sub_Sub_11_F_in3[2]) );
  AOI22_X1 Midori_rounds_U688 ( .A1(reset), .A2(Midori_add_Result_Start3[47]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[47]), .ZN(
        Midori_rounds_n1540) );
  XOR2_X1 Midori_rounds_U687 ( .A(Midori_rounds_SR_Inv_Result3[7]), .B(
        Midori_rounds_n1539), .Z(Midori_rounds_n1541) );
  OAI21_X1 Midori_rounds_U686 ( .B1(Midori_rounds_n1538), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1537), .ZN(Midori_rounds_n965)
         );
  AOI22_X1 Midori_rounds_U685 ( .A1(reset), .A2(Midori_add_Result_Start3[48]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[48]), .ZN(
        Midori_rounds_n1537) );
  XOR2_X1 Midori_rounds_U684 ( .A(Midori_rounds_SR_Inv_Result3[0]), .B(
        Midori_rounds_n1536), .Z(Midori_rounds_n1538) );
  OAI21_X1 Midori_rounds_U683 ( .B1(Midori_rounds_n1535), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1534), .ZN(
        Midori_rounds_sub_Sub_12_F_in3[0]) );
  AOI22_X1 Midori_rounds_U682 ( .A1(reset), .A2(Midori_add_Result_Start3[49]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[49]), .ZN(
        Midori_rounds_n1534) );
  XOR2_X1 Midori_rounds_U681 ( .A(Midori_rounds_SR_Inv_Result3[1]), .B(
        Midori_rounds_n1533), .Z(Midori_rounds_n1535) );
  OAI21_X1 Midori_rounds_U680 ( .B1(Midori_rounds_n1532), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1531), .ZN(Midori_rounds_n967)
         );
  AOI22_X1 Midori_rounds_U679 ( .A1(reset), .A2(Midori_add_Result_Start3[50]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[50]), .ZN(
        Midori_rounds_n1531) );
  XOR2_X1 Midori_rounds_U678 ( .A(Midori_rounds_SR_Inv_Result3[2]), .B(
        Midori_rounds_n1530), .Z(Midori_rounds_n1532) );
  OAI21_X1 Midori_rounds_U677 ( .B1(Midori_rounds_n1529), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1528), .ZN(
        Midori_rounds_sub_Sub_12_F_in3[2]) );
  AOI22_X1 Midori_rounds_U676 ( .A1(reset), .A2(Midori_add_Result_Start3[51]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[51]), .ZN(
        Midori_rounds_n1528) );
  XOR2_X1 Midori_rounds_U675 ( .A(Midori_rounds_SR_Inv_Result3[3]), .B(
        Midori_rounds_n1527), .Z(Midori_rounds_n1529) );
  OAI21_X1 Midori_rounds_U674 ( .B1(Midori_rounds_n1526), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1525), .ZN(Midori_rounds_n969)
         );
  AOI22_X1 Midori_rounds_U673 ( .A1(reset), .A2(Midori_add_Result_Start3[52]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[52]), .ZN(
        Midori_rounds_n1525) );
  XOR2_X1 Midori_rounds_U672 ( .A(Midori_rounds_SR_Inv_Result3[40]), .B(
        Midori_rounds_n1524), .Z(Midori_rounds_n1526) );
  OAI21_X1 Midori_rounds_U671 ( .B1(Midori_rounds_n1523), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1522), .ZN(
        Midori_rounds_sub_Sub_13_F_in3[0]) );
  AOI22_X1 Midori_rounds_U670 ( .A1(reset), .A2(Midori_add_Result_Start3[53]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[53]), .ZN(
        Midori_rounds_n1522) );
  XOR2_X1 Midori_rounds_U669 ( .A(Midori_rounds_SR_Inv_Result3[41]), .B(
        Midori_rounds_n1521), .Z(Midori_rounds_n1523) );
  OAI21_X1 Midori_rounds_U668 ( .B1(Midori_rounds_n1520), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1519), .ZN(Midori_rounds_n971)
         );
  AOI22_X1 Midori_rounds_U667 ( .A1(reset), .A2(Midori_add_Result_Start3[54]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[54]), .ZN(
        Midori_rounds_n1519) );
  XOR2_X1 Midori_rounds_U666 ( .A(Midori_rounds_SR_Inv_Result3[42]), .B(
        Midori_rounds_n1518), .Z(Midori_rounds_n1520) );
  OAI21_X1 Midori_rounds_U665 ( .B1(Midori_rounds_n1517), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1516), .ZN(
        Midori_rounds_sub_Sub_13_F_in3[2]) );
  AOI22_X1 Midori_rounds_U664 ( .A1(reset), .A2(Midori_add_Result_Start3[55]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[55]), .ZN(
        Midori_rounds_n1516) );
  XOR2_X1 Midori_rounds_U663 ( .A(Midori_rounds_SR_Inv_Result3[43]), .B(
        Midori_rounds_n1515), .Z(Midori_rounds_n1517) );
  OAI21_X1 Midori_rounds_U662 ( .B1(Midori_rounds_n1514), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1513), .ZN(Midori_rounds_n973)
         );
  AOI22_X1 Midori_rounds_U661 ( .A1(reset), .A2(Midori_add_Result_Start3[56]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[56]), .ZN(
        Midori_rounds_n1513) );
  XOR2_X1 Midori_rounds_U660 ( .A(Midori_rounds_SR_Inv_Result3[20]), .B(
        Midori_rounds_n1512), .Z(Midori_rounds_n1514) );
  OAI21_X1 Midori_rounds_U659 ( .B1(Midori_rounds_n1511), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1510), .ZN(
        Midori_rounds_sub_Sub_14_F_in3[0]) );
  AOI22_X1 Midori_rounds_U658 ( .A1(reset), .A2(Midori_add_Result_Start3[57]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[57]), .ZN(
        Midori_rounds_n1510) );
  XOR2_X1 Midori_rounds_U657 ( .A(Midori_rounds_SR_Inv_Result3[21]), .B(
        Midori_rounds_n1509), .Z(Midori_rounds_n1511) );
  OAI21_X1 Midori_rounds_U656 ( .B1(Midori_rounds_n1508), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1507), .ZN(Midori_rounds_n975)
         );
  AOI22_X1 Midori_rounds_U655 ( .A1(reset), .A2(Midori_add_Result_Start3[58]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[58]), .ZN(
        Midori_rounds_n1507) );
  XOR2_X1 Midori_rounds_U654 ( .A(Midori_rounds_SR_Inv_Result3[22]), .B(
        Midori_rounds_n1506), .Z(Midori_rounds_n1508) );
  OAI21_X1 Midori_rounds_U653 ( .B1(Midori_rounds_n1505), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1504), .ZN(
        Midori_rounds_sub_Sub_14_F_in3[2]) );
  AOI22_X1 Midori_rounds_U652 ( .A1(reset), .A2(Midori_add_Result_Start3[59]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[59]), .ZN(
        Midori_rounds_n1504) );
  XOR2_X1 Midori_rounds_U651 ( .A(Midori_rounds_SR_Inv_Result3[23]), .B(
        Midori_rounds_n1503), .Z(Midori_rounds_n1505) );
  OAI21_X1 Midori_rounds_U650 ( .B1(Midori_rounds_n1502), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1501), .ZN(Midori_rounds_n977)
         );
  AOI22_X1 Midori_rounds_U649 ( .A1(reset), .A2(Midori_add_Result_Start3[60]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[60]), .ZN(
        Midori_rounds_n1501) );
  XOR2_X1 Midori_rounds_U648 ( .A(Midori_rounds_SR_Inv_Result3[60]), .B(
        Midori_rounds_n1500), .Z(Midori_rounds_n1502) );
  OAI21_X1 Midori_rounds_U647 ( .B1(Midori_rounds_n1499), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1498), .ZN(
        Midori_rounds_sub_Sub_15_F_in3[0]) );
  AOI22_X1 Midori_rounds_U646 ( .A1(reset), .A2(Midori_add_Result_Start3[61]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[61]), .ZN(
        Midori_rounds_n1498) );
  XOR2_X1 Midori_rounds_U645 ( .A(Midori_rounds_SR_Inv_Result3[61]), .B(
        Midori_rounds_n1497), .Z(Midori_rounds_n1499) );
  OAI21_X1 Midori_rounds_U644 ( .B1(Midori_rounds_n1496), .B2(
        Midori_rounds_n2067), .A(Midori_rounds_n1495), .ZN(Midori_rounds_n979)
         );
  AOI22_X1 Midori_rounds_U643 ( .A1(reset), .A2(Midori_add_Result_Start3[62]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[62]), .ZN(
        Midori_rounds_n1495) );
  XOR2_X1 Midori_rounds_U642 ( .A(Midori_rounds_SR_Inv_Result3[62]), .B(
        Midori_rounds_n1494), .Z(Midori_rounds_n1496) );
  OAI21_X1 Midori_rounds_U641 ( .B1(Midori_rounds_n1493), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1492), .ZN(
        Midori_rounds_sub_Sub_15_F_in3[2]) );
  AOI22_X1 Midori_rounds_U640 ( .A1(reset), .A2(Midori_add_Result_Start3[63]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[63]), .ZN(
        Midori_rounds_n1492) );
  XOR2_X1 Midori_rounds_U639 ( .A(Midori_rounds_SR_Inv_Result3[63]), .B(
        Midori_rounds_n1490), .Z(Midori_rounds_n1493) );
  MUX2_X1 Midori_rounds_U638 ( .A(Midori_rounds_n1489), .B(
        Midori_rounds_SR_Result3[9]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[9]) );
  XNOR2_X1 Midori_rounds_U637 ( .A(Midori_rounds_SR_Result3[9]), .B(
        Midori_rounds_n1653), .ZN(Midori_rounds_n1489) );
  AOI22_X1 Midori_rounds_U636 ( .A1(Midori_rounds_n1272), .A2(Key3[9]), .B1(
        Key3[73]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1653) );
  MUX2_X1 Midori_rounds_U635 ( .A(Midori_rounds_n1488), .B(
        Midori_rounds_SR_Result3[8]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[8]) );
  XNOR2_X1 Midori_rounds_U634 ( .A(Midori_rounds_SR_Result3[8]), .B(
        Midori_rounds_n1656), .ZN(Midori_rounds_n1488) );
  AOI22_X1 Midori_rounds_U633 ( .A1(Midori_rounds_n1271), .A2(Key3[8]), .B1(
        Key3[72]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1656) );
  MUX2_X1 Midori_rounds_U632 ( .A(Midori_rounds_n1487), .B(
        Midori_rounds_SR_Result3[7]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[7]) );
  XNOR2_X1 Midori_rounds_U631 ( .A(Midori_rounds_SR_Result3[47]), .B(
        Midori_rounds_n1659), .ZN(Midori_rounds_n1487) );
  AOI22_X1 Midori_rounds_U630 ( .A1(Midori_rounds_n1272), .A2(Key3[7]), .B1(
        Key3[71]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1659) );
  MUX2_X1 Midori_rounds_U629 ( .A(Midori_rounds_n1486), .B(
        Midori_rounds_SR_Result3[6]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[6]) );
  XNOR2_X1 Midori_rounds_U628 ( .A(Midori_rounds_SR_Result3[46]), .B(
        Midori_rounds_n1662), .ZN(Midori_rounds_n1486) );
  AOI22_X1 Midori_rounds_U627 ( .A1(Midori_rounds_n1269), .A2(Key3[6]), .B1(
        Key3[70]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1662) );
  MUX2_X1 Midori_rounds_U626 ( .A(Midori_rounds_n1485), .B(
        Midori_rounds_SR_Result3[63]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[63]) );
  XNOR2_X1 Midori_rounds_U625 ( .A(Midori_rounds_SR_Result3[63]), .B(
        Midori_rounds_n1490), .ZN(Midori_rounds_n1485) );
  AOI22_X1 Midori_rounds_U624 ( .A1(Midori_rounds_n1275), .A2(Key3[63]), .B1(
        Key3[127]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1490) );
  MUX2_X1 Midori_rounds_U623 ( .A(Midori_rounds_n1484), .B(
        Midori_rounds_SR_Result3[62]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[62]) );
  XNOR2_X1 Midori_rounds_U622 ( .A(Midori_rounds_SR_Result3[62]), .B(
        Midori_rounds_n1494), .ZN(Midori_rounds_n1484) );
  AOI22_X1 Midori_rounds_U621 ( .A1(Midori_rounds_n1275), .A2(Key3[62]), .B1(
        Key3[126]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1494) );
  MUX2_X1 Midori_rounds_U620 ( .A(Midori_rounds_n1483), .B(
        Midori_rounds_SR_Result3[61]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[61]) );
  XNOR2_X1 Midori_rounds_U619 ( .A(Midori_rounds_SR_Result3[61]), .B(
        Midori_rounds_n1497), .ZN(Midori_rounds_n1483) );
  AOI22_X1 Midori_rounds_U618 ( .A1(Midori_rounds_n1274), .A2(Key3[61]), .B1(
        Key3[125]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1497) );
  MUX2_X1 Midori_rounds_U617 ( .A(Midori_rounds_n1482), .B(
        Midori_rounds_SR_Result3[60]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[60]) );
  XNOR2_X1 Midori_rounds_U616 ( .A(Midori_rounds_SR_Result3[60]), .B(
        Midori_rounds_n1500), .ZN(Midori_rounds_n1482) );
  AOI22_X1 Midori_rounds_U615 ( .A1(Midori_rounds_n1274), .A2(Key3[60]), .B1(
        Key3[124]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1500) );
  MUX2_X1 Midori_rounds_U614 ( .A(Midori_rounds_n1481), .B(
        Midori_rounds_SR_Result3[5]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[5]) );
  XNOR2_X1 Midori_rounds_U613 ( .A(Midori_rounds_SR_Result3[45]), .B(
        Midori_rounds_n1665), .ZN(Midori_rounds_n1481) );
  AOI22_X1 Midori_rounds_U612 ( .A1(Midori_rounds_n1271), .A2(Key3[5]), .B1(
        Key3[69]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1665) );
  MUX2_X1 Midori_rounds_U611 ( .A(Midori_rounds_n1480), .B(
        Midori_rounds_SR_Result3[59]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[59]) );
  XNOR2_X1 Midori_rounds_U610 ( .A(Midori_rounds_SR_Result3[35]), .B(
        Midori_rounds_n1503), .ZN(Midori_rounds_n1480) );
  AOI22_X1 Midori_rounds_U609 ( .A1(Midori_rounds_n1273), .A2(Key3[59]), .B1(
        Key3[123]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1503) );
  MUX2_X1 Midori_rounds_U608 ( .A(Midori_rounds_n1479), .B(
        Midori_rounds_SR_Result3[58]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[58]) );
  XNOR2_X1 Midori_rounds_U607 ( .A(Midori_rounds_SR_Result3[34]), .B(
        Midori_rounds_n1506), .ZN(Midori_rounds_n1479) );
  AOI22_X1 Midori_rounds_U606 ( .A1(Midori_rounds_n1272), .A2(Key3[58]), .B1(
        Key3[122]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1506) );
  MUX2_X1 Midori_rounds_U605 ( .A(Midori_rounds_n1478), .B(
        Midori_rounds_SR_Result3[57]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[57]) );
  XNOR2_X1 Midori_rounds_U604 ( .A(Midori_rounds_SR_Result3[33]), .B(
        Midori_rounds_n1509), .ZN(Midori_rounds_n1478) );
  AOI22_X1 Midori_rounds_U603 ( .A1(Midori_rounds_n1275), .A2(Key3[57]), .B1(
        Key3[121]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1509) );
  MUX2_X1 Midori_rounds_U602 ( .A(Midori_rounds_n1477), .B(
        Midori_rounds_SR_Result3[56]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input3[56]) );
  XNOR2_X1 Midori_rounds_U601 ( .A(Midori_rounds_SR_Result3[32]), .B(
        Midori_rounds_n1512), .ZN(Midori_rounds_n1477) );
  AOI22_X1 Midori_rounds_U600 ( .A1(Midori_rounds_n1272), .A2(Key3[56]), .B1(
        Key3[120]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1512) );
  MUX2_X1 Midori_rounds_U599 ( .A(Midori_rounds_n1476), .B(
        Midori_rounds_SR_Result3[55]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input3[55]) );
  XNOR2_X1 Midori_rounds_U598 ( .A(Midori_rounds_SR_Result3[7]), .B(
        Midori_rounds_n1515), .ZN(Midori_rounds_n1476) );
  AOI22_X1 Midori_rounds_U597 ( .A1(Midori_rounds_n1273), .A2(Key3[55]), .B1(
        Key3[119]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1515) );
  MUX2_X1 Midori_rounds_U596 ( .A(Midori_rounds_n1475), .B(
        Midori_rounds_SR_Result3[54]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[54]) );
  XNOR2_X1 Midori_rounds_U595 ( .A(Midori_rounds_SR_Result3[6]), .B(
        Midori_rounds_n1518), .ZN(Midori_rounds_n1475) );
  AOI22_X1 Midori_rounds_U594 ( .A1(Midori_rounds_n1272), .A2(Key3[54]), .B1(
        Key3[118]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1518) );
  MUX2_X1 Midori_rounds_U593 ( .A(Midori_rounds_n1474), .B(
        Midori_rounds_SR_Result3[53]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input3[53]) );
  XNOR2_X1 Midori_rounds_U592 ( .A(Midori_rounds_SR_Result3[5]), .B(
        Midori_rounds_n1521), .ZN(Midori_rounds_n1474) );
  AOI22_X1 Midori_rounds_U591 ( .A1(Midori_rounds_n1273), .A2(Key3[53]), .B1(
        Key3[117]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1521) );
  MUX2_X1 Midori_rounds_U590 ( .A(Midori_rounds_n1473), .B(
        Midori_rounds_SR_Result3[52]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input3[52]) );
  XNOR2_X1 Midori_rounds_U589 ( .A(Midori_rounds_SR_Result3[4]), .B(
        Midori_rounds_n1524), .ZN(Midori_rounds_n1473) );
  AOI22_X1 Midori_rounds_U588 ( .A1(Midori_rounds_n1274), .A2(Key3[52]), .B1(
        Key3[116]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1524) );
  MUX2_X1 Midori_rounds_U587 ( .A(Midori_rounds_n1472), .B(
        Midori_rounds_SR_Result3[51]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[51]) );
  XNOR2_X1 Midori_rounds_U586 ( .A(Midori_rounds_SR_Result3[27]), .B(
        Midori_rounds_n1527), .ZN(Midori_rounds_n1472) );
  AOI22_X1 Midori_rounds_U585 ( .A1(Midori_rounds_n1270), .A2(Key3[51]), .B1(
        Key3[115]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1527) );
  MUX2_X1 Midori_rounds_U584 ( .A(Midori_rounds_n1471), .B(
        Midori_rounds_SR_Result3[50]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input3[50]) );
  XNOR2_X1 Midori_rounds_U583 ( .A(Midori_rounds_SR_Result3[26]), .B(
        Midori_rounds_n1530), .ZN(Midori_rounds_n1471) );
  AOI22_X1 Midori_rounds_U582 ( .A1(Midori_rounds_n1272), .A2(Key3[50]), .B1(
        Key3[114]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1530) );
  MUX2_X1 Midori_rounds_U581 ( .A(Midori_rounds_n1470), .B(
        Midori_rounds_SR_Result3[4]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[4]) );
  XNOR2_X1 Midori_rounds_U580 ( .A(Midori_rounds_SR_Result3[44]), .B(
        Midori_rounds_n1668), .ZN(Midori_rounds_n1470) );
  AOI22_X1 Midori_rounds_U579 ( .A1(Midori_rounds_n1275), .A2(Key3[4]), .B1(
        Key3[68]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1668) );
  MUX2_X1 Midori_rounds_U578 ( .A(Midori_rounds_n1469), .B(
        Midori_rounds_SR_Result3[49]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[49]) );
  XNOR2_X1 Midori_rounds_U577 ( .A(Midori_rounds_SR_Result3[25]), .B(
        Midori_rounds_n1533), .ZN(Midori_rounds_n1469) );
  AOI22_X1 Midori_rounds_U576 ( .A1(Midori_rounds_n1269), .A2(Key3[49]), .B1(
        Key3[113]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1533) );
  MUX2_X1 Midori_rounds_U575 ( .A(Midori_rounds_n1468), .B(
        Midori_rounds_SR_Result3[48]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input3[48]) );
  XNOR2_X1 Midori_rounds_U574 ( .A(Midori_rounds_SR_Result3[24]), .B(
        Midori_rounds_n1536), .ZN(Midori_rounds_n1468) );
  AOI22_X1 Midori_rounds_U573 ( .A1(Midori_rounds_n1273), .A2(Key3[48]), .B1(
        Key3[112]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1536) );
  MUX2_X1 Midori_rounds_U572 ( .A(Midori_rounds_n1467), .B(
        Midori_rounds_SR_Result3[47]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input3[47]) );
  XNOR2_X1 Midori_rounds_U571 ( .A(Midori_rounds_SR_Result3[43]), .B(
        Midori_rounds_n1539), .ZN(Midori_rounds_n1467) );
  AOI22_X1 Midori_rounds_U570 ( .A1(Midori_rounds_n1273), .A2(Key3[47]), .B1(
        Key3[111]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1539) );
  MUX2_X1 Midori_rounds_U569 ( .A(Midori_rounds_n1466), .B(
        Midori_rounds_SR_Result3[46]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input3[46]) );
  XNOR2_X1 Midori_rounds_U568 ( .A(Midori_rounds_SR_Result3[42]), .B(
        Midori_rounds_n1542), .ZN(Midori_rounds_n1466) );
  AOI22_X1 Midori_rounds_U567 ( .A1(Midori_rounds_n1271), .A2(Key3[46]), .B1(
        Key3[110]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1542) );
  MUX2_X1 Midori_rounds_U566 ( .A(Midori_rounds_n1465), .B(
        Midori_rounds_SR_Result3[45]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[45]) );
  XNOR2_X1 Midori_rounds_U565 ( .A(Midori_rounds_SR_Result3[41]), .B(
        Midori_rounds_n1545), .ZN(Midori_rounds_n1465) );
  AOI22_X1 Midori_rounds_U564 ( .A1(Midori_rounds_n1269), .A2(Key3[45]), .B1(
        Key3[109]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1545) );
  MUX2_X1 Midori_rounds_U563 ( .A(Midori_rounds_n1464), .B(
        Midori_rounds_SR_Result3[44]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[44]) );
  XNOR2_X1 Midori_rounds_U562 ( .A(Midori_rounds_SR_Result3[40]), .B(
        Midori_rounds_n1548), .ZN(Midori_rounds_n1464) );
  AOI22_X1 Midori_rounds_U561 ( .A1(Midori_rounds_n1269), .A2(Key3[44]), .B1(
        Key3[108]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1548) );
  MUX2_X1 Midori_rounds_U560 ( .A(Midori_rounds_n1463), .B(
        Midori_rounds_SR_Result3[43]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[43]) );
  XNOR2_X1 Midori_rounds_U559 ( .A(Midori_rounds_SR_Result3[55]), .B(
        Midori_rounds_n1551), .ZN(Midori_rounds_n1463) );
  AOI22_X1 Midori_rounds_U558 ( .A1(Midori_rounds_n1275), .A2(Key3[43]), .B1(
        Key3[107]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1551) );
  MUX2_X1 Midori_rounds_U557 ( .A(Midori_rounds_n1462), .B(
        Midori_rounds_SR_Result3[42]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[42]) );
  XNOR2_X1 Midori_rounds_U556 ( .A(Midori_rounds_SR_Result3[54]), .B(
        Midori_rounds_n1554), .ZN(Midori_rounds_n1462) );
  AOI22_X1 Midori_rounds_U555 ( .A1(Midori_rounds_n1270), .A2(Key3[42]), .B1(
        Key3[106]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1554) );
  MUX2_X1 Midori_rounds_U554 ( .A(Midori_rounds_n1461), .B(
        Midori_rounds_SR_Result3[41]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[41]) );
  XNOR2_X1 Midori_rounds_U553 ( .A(Midori_rounds_SR_Result3[53]), .B(
        Midori_rounds_n1557), .ZN(Midori_rounds_n1461) );
  AOI22_X1 Midori_rounds_U552 ( .A1(Midori_rounds_n1270), .A2(Key3[41]), .B1(
        Key3[105]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1557) );
  MUX2_X1 Midori_rounds_U551 ( .A(Midori_rounds_n1460), .B(
        Midori_rounds_SR_Result3[40]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[40]) );
  XNOR2_X1 Midori_rounds_U550 ( .A(Midori_rounds_SR_Result3[52]), .B(
        Midori_rounds_n1560), .ZN(Midori_rounds_n1460) );
  AOI22_X1 Midori_rounds_U549 ( .A1(Midori_rounds_n1273), .A2(Key3[40]), .B1(
        Key3[104]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1560) );
  MUX2_X1 Midori_rounds_U548 ( .A(Midori_rounds_n1459), .B(
        Midori_rounds_SR_Result3[3]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[3]) );
  XNOR2_X1 Midori_rounds_U547 ( .A(Midori_rounds_SR_Result3[51]), .B(
        Midori_rounds_n1671), .ZN(Midori_rounds_n1459) );
  AOI22_X1 Midori_rounds_U546 ( .A1(Midori_rounds_n1270), .A2(Key3[3]), .B1(
        Key3[67]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1671) );
  MUX2_X1 Midori_rounds_U545 ( .A(Midori_rounds_n1458), .B(
        Midori_rounds_SR_Result3[39]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[39]) );
  XNOR2_X1 Midori_rounds_U544 ( .A(Midori_rounds_SR_Result3[19]), .B(
        Midori_rounds_n1563), .ZN(Midori_rounds_n1458) );
  AOI22_X1 Midori_rounds_U543 ( .A1(Midori_rounds_n1274), .A2(Key3[39]), .B1(
        Key3[103]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1563) );
  MUX2_X1 Midori_rounds_U542 ( .A(Midori_rounds_n1457), .B(
        Midori_rounds_SR_Result3[38]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[38]) );
  XNOR2_X1 Midori_rounds_U541 ( .A(Midori_rounds_SR_Result3[18]), .B(
        Midori_rounds_n1566), .ZN(Midori_rounds_n1457) );
  AOI22_X1 Midori_rounds_U540 ( .A1(Midori_rounds_n1269), .A2(Key3[38]), .B1(
        Key3[102]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1566) );
  MUX2_X1 Midori_rounds_U539 ( .A(Midori_rounds_n1456), .B(
        Midori_rounds_SR_Result3[37]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[37]) );
  XNOR2_X1 Midori_rounds_U538 ( .A(Midori_rounds_SR_Result3[17]), .B(
        Midori_rounds_n1569), .ZN(Midori_rounds_n1456) );
  AOI22_X1 Midori_rounds_U537 ( .A1(Midori_rounds_n1270), .A2(Key3[37]), .B1(
        Key3[101]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1569) );
  MUX2_X1 Midori_rounds_U536 ( .A(Midori_rounds_n1455), .B(
        Midori_rounds_SR_Result3[36]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[36]) );
  XNOR2_X1 Midori_rounds_U535 ( .A(Midori_rounds_SR_Result3[16]), .B(
        Midori_rounds_n1572), .ZN(Midori_rounds_n1455) );
  AOI22_X1 Midori_rounds_U534 ( .A1(Midori_rounds_n1270), .A2(Key3[36]), .B1(
        Key3[100]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1572) );
  MUX2_X1 Midori_rounds_U533 ( .A(Midori_rounds_n1454), .B(
        Midori_rounds_SR_Result3[35]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[35]) );
  XNOR2_X1 Midori_rounds_U532 ( .A(Midori_rounds_SR_Result3[15]), .B(
        Midori_rounds_n1575), .ZN(Midori_rounds_n1454) );
  AOI22_X1 Midori_rounds_U531 ( .A1(Midori_rounds_n1269), .A2(Key3[35]), .B1(
        Key3[99]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1575) );
  MUX2_X1 Midori_rounds_U530 ( .A(Midori_rounds_n1453), .B(
        Midori_rounds_SR_Result3[34]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[34]) );
  XNOR2_X1 Midori_rounds_U529 ( .A(Midori_rounds_SR_Result3[14]), .B(
        Midori_rounds_n1578), .ZN(Midori_rounds_n1453) );
  AOI22_X1 Midori_rounds_U528 ( .A1(Midori_rounds_n1270), .A2(Key3[34]), .B1(
        Key3[98]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1578) );
  MUX2_X1 Midori_rounds_U527 ( .A(Midori_rounds_n1452), .B(
        Midori_rounds_SR_Result3[33]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[33]) );
  XNOR2_X1 Midori_rounds_U526 ( .A(Midori_rounds_SR_Result3[13]), .B(
        Midori_rounds_n1581), .ZN(Midori_rounds_n1452) );
  AOI22_X1 Midori_rounds_U525 ( .A1(Midori_rounds_n1275), .A2(Key3[33]), .B1(
        Key3[97]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1581) );
  MUX2_X1 Midori_rounds_U524 ( .A(Midori_rounds_n1451), .B(
        Midori_rounds_SR_Result3[32]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[32]) );
  XNOR2_X1 Midori_rounds_U523 ( .A(Midori_rounds_SR_Result3[12]), .B(
        Midori_rounds_n1584), .ZN(Midori_rounds_n1451) );
  AOI22_X1 Midori_rounds_U522 ( .A1(Midori_rounds_n1275), .A2(Key3[32]), .B1(
        Key3[96]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1584) );
  MUX2_X1 Midori_rounds_U521 ( .A(Midori_rounds_n1450), .B(
        Midori_rounds_SR_Result3[31]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[31]) );
  XNOR2_X1 Midori_rounds_U520 ( .A(Midori_rounds_SR_Result3[3]), .B(
        Midori_rounds_n1587), .ZN(Midori_rounds_n1450) );
  AOI22_X1 Midori_rounds_U519 ( .A1(Midori_rounds_n1275), .A2(Key3[31]), .B1(
        Key3[95]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1587) );
  MUX2_X1 Midori_rounds_U518 ( .A(Midori_rounds_n1449), .B(
        Midori_rounds_SR_Result3[30]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[30]) );
  XNOR2_X1 Midori_rounds_U517 ( .A(Midori_rounds_SR_Result3[2]), .B(
        Midori_rounds_n1590), .ZN(Midori_rounds_n1449) );
  AOI22_X1 Midori_rounds_U516 ( .A1(Midori_rounds_n1275), .A2(Key3[30]), .B1(
        Key3[94]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1590) );
  MUX2_X1 Midori_rounds_U515 ( .A(Midori_rounds_n1448), .B(
        Midori_rounds_SR_Result3[2]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[2]) );
  XNOR2_X1 Midori_rounds_U514 ( .A(Midori_rounds_SR_Result3[50]), .B(
        Midori_rounds_n1674), .ZN(Midori_rounds_n1448) );
  AOI22_X1 Midori_rounds_U513 ( .A1(Midori_rounds_n1275), .A2(Key3[2]), .B1(
        Key3[66]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1674) );
  MUX2_X1 Midori_rounds_U512 ( .A(Midori_rounds_n1447), .B(
        Midori_rounds_SR_Result3[29]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[29]) );
  XNOR2_X1 Midori_rounds_U511 ( .A(Midori_rounds_SR_Result3[1]), .B(
        Midori_rounds_n1593), .ZN(Midori_rounds_n1447) );
  AOI22_X1 Midori_rounds_U510 ( .A1(Midori_rounds_n1275), .A2(Key3[29]), .B1(
        Key3[93]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1593) );
  MUX2_X1 Midori_rounds_U509 ( .A(Midori_rounds_n1446), .B(
        Midori_rounds_SR_Result3[28]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[28]) );
  XNOR2_X1 Midori_rounds_U508 ( .A(Midori_rounds_SR_Result3[0]), .B(
        Midori_rounds_n1596), .ZN(Midori_rounds_n1446) );
  AOI22_X1 Midori_rounds_U507 ( .A1(Midori_rounds_n1275), .A2(Key3[28]), .B1(
        Key3[92]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1596) );
  MUX2_X1 Midori_rounds_U506 ( .A(Midori_rounds_n1445), .B(
        Midori_rounds_SR_Result3[27]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[27]) );
  XNOR2_X1 Midori_rounds_U505 ( .A(Midori_rounds_SR_Result3[31]), .B(
        Midori_rounds_n1599), .ZN(Midori_rounds_n1445) );
  AOI22_X1 Midori_rounds_U504 ( .A1(Midori_rounds_n1275), .A2(Key3[27]), .B1(
        Key3[91]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1599) );
  MUX2_X1 Midori_rounds_U503 ( .A(Midori_rounds_n1444), .B(
        Midori_rounds_SR_Result3[26]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[26]) );
  XNOR2_X1 Midori_rounds_U502 ( .A(Midori_rounds_SR_Result3[30]), .B(
        Midori_rounds_n1602), .ZN(Midori_rounds_n1444) );
  AOI22_X1 Midori_rounds_U501 ( .A1(Midori_rounds_n1275), .A2(Key3[26]), .B1(
        Key3[90]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1602) );
  MUX2_X1 Midori_rounds_U500 ( .A(Midori_rounds_n1443), .B(
        Midori_rounds_SR_Result3[25]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[25]) );
  XNOR2_X1 Midori_rounds_U499 ( .A(Midori_rounds_SR_Result3[29]), .B(
        Midori_rounds_n1605), .ZN(Midori_rounds_n1443) );
  AOI22_X1 Midori_rounds_U498 ( .A1(Midori_rounds_n1275), .A2(Key3[25]), .B1(
        Key3[89]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1605) );
  MUX2_X1 Midori_rounds_U497 ( .A(Midori_rounds_n1442), .B(
        Midori_rounds_SR_Result3[24]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[24]) );
  XNOR2_X1 Midori_rounds_U496 ( .A(Midori_rounds_SR_Result3[28]), .B(
        Midori_rounds_n1608), .ZN(Midori_rounds_n1442) );
  AOI22_X1 Midori_rounds_U495 ( .A1(Midori_rounds_n1275), .A2(Key3[24]), .B1(
        Key3[88]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1608) );
  MUX2_X1 Midori_rounds_U494 ( .A(Midori_rounds_n1441), .B(
        Midori_rounds_SR_Result3[23]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[23]) );
  XNOR2_X1 Midori_rounds_U493 ( .A(Midori_rounds_SR_Result3[59]), .B(
        Midori_rounds_n1611), .ZN(Midori_rounds_n1441) );
  AOI22_X1 Midori_rounds_U492 ( .A1(Midori_rounds_n1275), .A2(Key3[23]), .B1(
        Key3[87]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1611) );
  MUX2_X1 Midori_rounds_U491 ( .A(Midori_rounds_n1440), .B(
        Midori_rounds_SR_Result3[22]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[22]) );
  XNOR2_X1 Midori_rounds_U490 ( .A(Midori_rounds_SR_Result3[58]), .B(
        Midori_rounds_n1614), .ZN(Midori_rounds_n1440) );
  AOI22_X1 Midori_rounds_U489 ( .A1(Midori_rounds_n1275), .A2(Key3[22]), .B1(
        Key3[86]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1614) );
  MUX2_X1 Midori_rounds_U488 ( .A(Midori_rounds_n1439), .B(
        Midori_rounds_SR_Result3[21]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[21]) );
  XNOR2_X1 Midori_rounds_U487 ( .A(Midori_rounds_SR_Result3[57]), .B(
        Midori_rounds_n1617), .ZN(Midori_rounds_n1439) );
  AOI22_X1 Midori_rounds_U486 ( .A1(Midori_rounds_n1274), .A2(Key3[21]), .B1(
        Key3[85]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1617) );
  MUX2_X1 Midori_rounds_U485 ( .A(Midori_rounds_n1438), .B(
        Midori_rounds_SR_Result3[20]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[20]) );
  XNOR2_X1 Midori_rounds_U484 ( .A(Midori_rounds_SR_Result3[56]), .B(
        Midori_rounds_n1620), .ZN(Midori_rounds_n1438) );
  AOI22_X1 Midori_rounds_U483 ( .A1(Midori_rounds_n1274), .A2(Key3[20]), .B1(
        Key3[84]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1620) );
  MUX2_X1 Midori_rounds_U482 ( .A(Midori_rounds_n1437), .B(
        Midori_rounds_SR_Result3[1]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[1]) );
  XNOR2_X1 Midori_rounds_U481 ( .A(Midori_rounds_SR_Result3[49]), .B(
        Midori_rounds_n1677), .ZN(Midori_rounds_n1437) );
  AOI22_X1 Midori_rounds_U480 ( .A1(Midori_rounds_n1274), .A2(Key3[1]), .B1(
        Key3[65]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1677) );
  MUX2_X1 Midori_rounds_U479 ( .A(Midori_rounds_n1436), .B(
        Midori_rounds_SR_Result3[19]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[19]) );
  XNOR2_X1 Midori_rounds_U478 ( .A(Midori_rounds_SR_Result3[39]), .B(
        Midori_rounds_n1623), .ZN(Midori_rounds_n1436) );
  AOI22_X1 Midori_rounds_U477 ( .A1(Midori_rounds_n1274), .A2(Key3[19]), .B1(
        Key3[83]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1623) );
  MUX2_X1 Midori_rounds_U476 ( .A(Midori_rounds_n1435), .B(
        Midori_rounds_SR_Result3[18]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[18]) );
  XNOR2_X1 Midori_rounds_U475 ( .A(Midori_rounds_SR_Result3[38]), .B(
        Midori_rounds_n1626), .ZN(Midori_rounds_n1435) );
  AOI22_X1 Midori_rounds_U474 ( .A1(Midori_rounds_n1274), .A2(Key3[18]), .B1(
        Key3[82]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1626) );
  MUX2_X1 Midori_rounds_U473 ( .A(Midori_rounds_n1434), .B(
        Midori_rounds_SR_Result3[17]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[17]) );
  XNOR2_X1 Midori_rounds_U472 ( .A(Midori_rounds_SR_Result3[37]), .B(
        Midori_rounds_n1629), .ZN(Midori_rounds_n1434) );
  AOI22_X1 Midori_rounds_U471 ( .A1(Midori_rounds_n1274), .A2(Key3[17]), .B1(
        Key3[81]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1629) );
  MUX2_X1 Midori_rounds_U470 ( .A(Midori_rounds_n1433), .B(
        Midori_rounds_SR_Result3[16]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[16]) );
  XNOR2_X1 Midori_rounds_U469 ( .A(Midori_rounds_SR_Result3[36]), .B(
        Midori_rounds_n1632), .ZN(Midori_rounds_n1433) );
  AOI22_X1 Midori_rounds_U468 ( .A1(Midori_rounds_n1274), .A2(Key3[16]), .B1(
        Key3[80]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1632) );
  MUX2_X1 Midori_rounds_U467 ( .A(Midori_rounds_n1432), .B(
        Midori_rounds_SR_Result3[15]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[15]) );
  XNOR2_X1 Midori_rounds_U466 ( .A(Midori_rounds_SR_Result3[23]), .B(
        Midori_rounds_n1635), .ZN(Midori_rounds_n1432) );
  AOI22_X1 Midori_rounds_U465 ( .A1(Midori_rounds_n1274), .A2(Key3[15]), .B1(
        Key3[79]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1635) );
  MUX2_X1 Midori_rounds_U464 ( .A(Midori_rounds_n1431), .B(
        Midori_rounds_SR_Result3[14]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[14]) );
  XNOR2_X1 Midori_rounds_U463 ( .A(Midori_rounds_SR_Result3[22]), .B(
        Midori_rounds_n1638), .ZN(Midori_rounds_n1431) );
  AOI22_X1 Midori_rounds_U462 ( .A1(Midori_rounds_n1274), .A2(Key3[14]), .B1(
        Key3[78]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1638) );
  MUX2_X1 Midori_rounds_U461 ( .A(Midori_rounds_n1430), .B(
        Midori_rounds_SR_Result3[13]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[13]) );
  XNOR2_X1 Midori_rounds_U460 ( .A(Midori_rounds_SR_Result3[21]), .B(
        Midori_rounds_n1641), .ZN(Midori_rounds_n1430) );
  AOI22_X1 Midori_rounds_U459 ( .A1(Midori_rounds_n1274), .A2(Key3[13]), .B1(
        Key3[77]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1641) );
  MUX2_X1 Midori_rounds_U458 ( .A(Midori_rounds_n1429), .B(
        Midori_rounds_SR_Result3[12]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[12]) );
  XNOR2_X1 Midori_rounds_U457 ( .A(Midori_rounds_SR_Result3[20]), .B(
        Midori_rounds_n1644), .ZN(Midori_rounds_n1429) );
  AOI22_X1 Midori_rounds_U456 ( .A1(Midori_rounds_n1274), .A2(Key3[12]), .B1(
        Key3[76]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1644) );
  MUX2_X1 Midori_rounds_U455 ( .A(Midori_rounds_n1428), .B(
        Midori_rounds_SR_Result3[11]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[11]) );
  XNOR2_X1 Midori_rounds_U454 ( .A(Midori_rounds_SR_Result3[11]), .B(
        Midori_rounds_n1647), .ZN(Midori_rounds_n1428) );
  AOI22_X1 Midori_rounds_U453 ( .A1(Midori_rounds_n1274), .A2(Key3[11]), .B1(
        Key3[75]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1647) );
  MUX2_X1 Midori_rounds_U452 ( .A(Midori_rounds_n1427), .B(
        Midori_rounds_SR_Result3[10]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[10]) );
  XNOR2_X1 Midori_rounds_U451 ( .A(Midori_rounds_SR_Result3[10]), .B(
        Midori_rounds_n1650), .ZN(Midori_rounds_n1427) );
  AOI22_X1 Midori_rounds_U450 ( .A1(Midori_rounds_n1274), .A2(Key3[10]), .B1(
        Key3[74]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1650) );
  MUX2_X1 Midori_rounds_U449 ( .A(Midori_rounds_n1426), .B(
        Midori_rounds_SR_Result3[0]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input3[0]) );
  XNOR2_X1 Midori_rounds_U448 ( .A(Midori_rounds_SR_Result3[48]), .B(
        Midori_rounds_n1680), .ZN(Midori_rounds_n1426) );
  AOI22_X1 Midori_rounds_U447 ( .A1(Midori_rounds_n1273), .A2(Key3[0]), .B1(
        Key3[64]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1680) );
  MUX2_X1 Midori_rounds_U446 ( .A(Midori_rounds_n1425), .B(
        Midori_rounds_SR_Result2[9]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[9]) );
  XNOR2_X1 Midori_rounds_U445 ( .A(Midori_rounds_SR_Result2[9]), .B(
        Midori_rounds_n1845), .ZN(Midori_rounds_n1425) );
  AOI22_X1 Midori_rounds_U444 ( .A1(Midori_rounds_n1273), .A2(Key2[9]), .B1(
        Key2[73]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1845) );
  MUX2_X1 Midori_rounds_U443 ( .A(Midori_rounds_n1424), .B(
        Midori_rounds_SR_Result2[8]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[8]) );
  XNOR2_X1 Midori_rounds_U442 ( .A(Midori_rounds_SR_Result2[8]), .B(
        Midori_rounds_n1848), .ZN(Midori_rounds_n1424) );
  AOI22_X1 Midori_rounds_U441 ( .A1(Midori_rounds_n1273), .A2(Key2[8]), .B1(
        Key2[72]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1848) );
  MUX2_X1 Midori_rounds_U440 ( .A(Midori_rounds_n1423), .B(
        Midori_rounds_SR_Result2[7]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[7]) );
  XNOR2_X1 Midori_rounds_U439 ( .A(Midori_rounds_SR_Result2[47]), .B(
        Midori_rounds_n1851), .ZN(Midori_rounds_n1423) );
  AOI22_X1 Midori_rounds_U438 ( .A1(Midori_rounds_n1273), .A2(Key2[7]), .B1(
        Key2[71]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1851) );
  MUX2_X1 Midori_rounds_U437 ( .A(Midori_rounds_n1422), .B(
        Midori_rounds_SR_Result2[6]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input2[6]) );
  XNOR2_X1 Midori_rounds_U436 ( .A(Midori_rounds_SR_Result2[46]), .B(
        Midori_rounds_n1854), .ZN(Midori_rounds_n1422) );
  AOI22_X1 Midori_rounds_U435 ( .A1(Midori_rounds_n1273), .A2(Key2[6]), .B1(
        Key2[70]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1854) );
  MUX2_X1 Midori_rounds_U434 ( .A(Midori_rounds_n1421), .B(
        Midori_rounds_SR_Result2[63]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[63]) );
  XNOR2_X1 Midori_rounds_U433 ( .A(Midori_rounds_SR_Result2[63]), .B(
        Midori_rounds_n1683), .ZN(Midori_rounds_n1421) );
  AOI22_X1 Midori_rounds_U432 ( .A1(Midori_rounds_n1273), .A2(Key2[63]), .B1(
        Key2[127]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1683) );
  MUX2_X1 Midori_rounds_U431 ( .A(Midori_rounds_n1420), .B(
        Midori_rounds_SR_Result2[62]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[62]) );
  XNOR2_X1 Midori_rounds_U430 ( .A(Midori_rounds_SR_Result2[62]), .B(
        Midori_rounds_n1686), .ZN(Midori_rounds_n1420) );
  AOI22_X1 Midori_rounds_U429 ( .A1(Midori_rounds_n1273), .A2(Key2[62]), .B1(
        Key2[126]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1686) );
  MUX2_X1 Midori_rounds_U428 ( .A(Midori_rounds_n1419), .B(
        Midori_rounds_SR_Result2[61]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[61]) );
  XNOR2_X1 Midori_rounds_U427 ( .A(Midori_rounds_SR_Result2[61]), .B(
        Midori_rounds_n1689), .ZN(Midori_rounds_n1419) );
  AOI22_X1 Midori_rounds_U426 ( .A1(Midori_rounds_n1273), .A2(Key2[61]), .B1(
        Key2[125]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1689) );
  MUX2_X1 Midori_rounds_U425 ( .A(Midori_rounds_n1418), .B(
        Midori_rounds_SR_Result2[60]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[60]) );
  XNOR2_X1 Midori_rounds_U424 ( .A(Midori_rounds_SR_Result2[60]), .B(
        Midori_rounds_n1692), .ZN(Midori_rounds_n1418) );
  AOI22_X1 Midori_rounds_U423 ( .A1(Midori_rounds_n1273), .A2(Key2[60]), .B1(
        Key2[124]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1692) );
  MUX2_X1 Midori_rounds_U422 ( .A(Midori_rounds_n1417), .B(
        Midori_rounds_SR_Result2[5]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[5]) );
  XNOR2_X1 Midori_rounds_U421 ( .A(Midori_rounds_SR_Result2[45]), .B(
        Midori_rounds_n1857), .ZN(Midori_rounds_n1417) );
  AOI22_X1 Midori_rounds_U420 ( .A1(Midori_rounds_n1273), .A2(Key2[5]), .B1(
        Key2[69]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1857) );
  MUX2_X1 Midori_rounds_U419 ( .A(Midori_rounds_n1416), .B(
        Midori_rounds_SR_Result2[59]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input2[59]) );
  XNOR2_X1 Midori_rounds_U418 ( .A(Midori_rounds_SR_Result2[35]), .B(
        Midori_rounds_n1695), .ZN(Midori_rounds_n1416) );
  AOI22_X1 Midori_rounds_U417 ( .A1(Midori_rounds_n1273), .A2(Key2[59]), .B1(
        Key2[123]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1695) );
  MUX2_X1 Midori_rounds_U416 ( .A(Midori_rounds_n1415), .B(
        Midori_rounds_SR_Result2[58]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[58]) );
  XNOR2_X1 Midori_rounds_U415 ( .A(Midori_rounds_SR_Result2[34]), .B(
        Midori_rounds_n1698), .ZN(Midori_rounds_n1415) );
  AOI22_X1 Midori_rounds_U414 ( .A1(Midori_rounds_n1273), .A2(Key2[58]), .B1(
        Key2[122]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1698) );
  MUX2_X1 Midori_rounds_U413 ( .A(Midori_rounds_n1414), .B(
        Midori_rounds_SR_Result2[57]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[57]) );
  XNOR2_X1 Midori_rounds_U412 ( .A(Midori_rounds_SR_Result2[33]), .B(
        Midori_rounds_n1701), .ZN(Midori_rounds_n1414) );
  AOI22_X1 Midori_rounds_U411 ( .A1(Midori_rounds_n1273), .A2(Key2[57]), .B1(
        Key2[121]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1701) );
  MUX2_X1 Midori_rounds_U410 ( .A(Midori_rounds_n1413), .B(
        Midori_rounds_SR_Result2[56]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input2[56]) );
  XNOR2_X1 Midori_rounds_U409 ( .A(Midori_rounds_SR_Result2[32]), .B(
        Midori_rounds_n1704), .ZN(Midori_rounds_n1413) );
  AOI22_X1 Midori_rounds_U408 ( .A1(Midori_rounds_n1272), .A2(Key2[56]), .B1(
        Key2[120]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1704) );
  MUX2_X1 Midori_rounds_U407 ( .A(Midori_rounds_n1412), .B(
        Midori_rounds_SR_Result2[55]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[55]) );
  XNOR2_X1 Midori_rounds_U406 ( .A(Midori_rounds_SR_Result2[7]), .B(
        Midori_rounds_n1707), .ZN(Midori_rounds_n1412) );
  AOI22_X1 Midori_rounds_U405 ( .A1(Midori_rounds_n1272), .A2(Key2[55]), .B1(
        Key2[119]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1707) );
  MUX2_X1 Midori_rounds_U404 ( .A(Midori_rounds_n1411), .B(
        Midori_rounds_SR_Result2[54]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[54]) );
  XNOR2_X1 Midori_rounds_U403 ( .A(Midori_rounds_SR_Result2[6]), .B(
        Midori_rounds_n1710), .ZN(Midori_rounds_n1411) );
  AOI22_X1 Midori_rounds_U402 ( .A1(Midori_rounds_n1272), .A2(Key2[54]), .B1(
        Key2[118]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1710) );
  MUX2_X1 Midori_rounds_U401 ( .A(Midori_rounds_n1410), .B(
        Midori_rounds_SR_Result2[53]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[53]) );
  XNOR2_X1 Midori_rounds_U400 ( .A(Midori_rounds_SR_Result2[5]), .B(
        Midori_rounds_n1713), .ZN(Midori_rounds_n1410) );
  AOI22_X1 Midori_rounds_U399 ( .A1(Midori_rounds_n1272), .A2(Key2[53]), .B1(
        Key2[117]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1713) );
  MUX2_X1 Midori_rounds_U398 ( .A(Midori_rounds_n1409), .B(
        Midori_rounds_SR_Result2[52]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[52]) );
  XNOR2_X1 Midori_rounds_U397 ( .A(Midori_rounds_SR_Result2[4]), .B(
        Midori_rounds_n1716), .ZN(Midori_rounds_n1409) );
  AOI22_X1 Midori_rounds_U396 ( .A1(Midori_rounds_n1272), .A2(Key2[52]), .B1(
        Key2[116]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1716) );
  MUX2_X1 Midori_rounds_U395 ( .A(Midori_rounds_n1408), .B(
        Midori_rounds_SR_Result2[51]), .S(Midori_rounds_n1491), .Z(
        Midori_rounds_mul_input2[51]) );
  XNOR2_X1 Midori_rounds_U394 ( .A(Midori_rounds_SR_Result2[27]), .B(
        Midori_rounds_n1719), .ZN(Midori_rounds_n1408) );
  AOI22_X1 Midori_rounds_U393 ( .A1(Midori_rounds_n1272), .A2(Key2[51]), .B1(
        Key2[115]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1719) );
  MUX2_X1 Midori_rounds_U392 ( .A(Midori_rounds_n1407), .B(
        Midori_rounds_SR_Result2[50]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[50]) );
  XNOR2_X1 Midori_rounds_U391 ( .A(Midori_rounds_SR_Result2[26]), .B(
        Midori_rounds_n1722), .ZN(Midori_rounds_n1407) );
  AOI22_X1 Midori_rounds_U390 ( .A1(Midori_rounds_n1272), .A2(Key2[50]), .B1(
        Key2[114]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1722) );
  MUX2_X1 Midori_rounds_U389 ( .A(Midori_rounds_n1406), .B(
        Midori_rounds_SR_Result2[4]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[4]) );
  XNOR2_X1 Midori_rounds_U388 ( .A(Midori_rounds_SR_Result2[44]), .B(
        Midori_rounds_n1860), .ZN(Midori_rounds_n1406) );
  AOI22_X1 Midori_rounds_U387 ( .A1(Midori_rounds_n1272), .A2(Key2[4]), .B1(
        Key2[68]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1860) );
  MUX2_X1 Midori_rounds_U386 ( .A(Midori_rounds_n1405), .B(
        Midori_rounds_SR_Result2[49]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[49]) );
  XNOR2_X1 Midori_rounds_U385 ( .A(Midori_rounds_SR_Result2[25]), .B(
        Midori_rounds_n1725), .ZN(Midori_rounds_n1405) );
  AOI22_X1 Midori_rounds_U384 ( .A1(Midori_rounds_n1272), .A2(Key2[49]), .B1(
        Key2[113]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1725) );
  MUX2_X1 Midori_rounds_U383 ( .A(Midori_rounds_n1404), .B(
        Midori_rounds_SR_Result2[48]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[48]) );
  XNOR2_X1 Midori_rounds_U382 ( .A(Midori_rounds_SR_Result2[24]), .B(
        Midori_rounds_n1728), .ZN(Midori_rounds_n1404) );
  AOI22_X1 Midori_rounds_U381 ( .A1(Midori_rounds_n1272), .A2(Key2[48]), .B1(
        Key2[112]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1728) );
  MUX2_X1 Midori_rounds_U380 ( .A(Midori_rounds_n1403), .B(
        Midori_rounds_SR_Result2[47]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[47]) );
  XNOR2_X1 Midori_rounds_U379 ( .A(Midori_rounds_SR_Result2[43]), .B(
        Midori_rounds_n1731), .ZN(Midori_rounds_n1403) );
  AOI22_X1 Midori_rounds_U378 ( .A1(Midori_rounds_n1272), .A2(Key2[47]), .B1(
        Key2[111]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1731) );
  MUX2_X1 Midori_rounds_U377 ( .A(Midori_rounds_n1402), .B(
        Midori_rounds_SR_Result2[46]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[46]) );
  XNOR2_X1 Midori_rounds_U376 ( .A(Midori_rounds_SR_Result2[42]), .B(
        Midori_rounds_n1734), .ZN(Midori_rounds_n1402) );
  AOI22_X1 Midori_rounds_U375 ( .A1(Midori_rounds_n1272), .A2(Key2[46]), .B1(
        Key2[110]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1734) );
  MUX2_X1 Midori_rounds_U374 ( .A(Midori_rounds_n1401), .B(
        Midori_rounds_SR_Result2[45]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[45]) );
  XNOR2_X1 Midori_rounds_U373 ( .A(Midori_rounds_SR_Result2[41]), .B(
        Midori_rounds_n1737), .ZN(Midori_rounds_n1401) );
  AOI22_X1 Midori_rounds_U372 ( .A1(Midori_rounds_n1272), .A2(Key2[45]), .B1(
        Key2[109]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1737) );
  MUX2_X1 Midori_rounds_U371 ( .A(Midori_rounds_n1400), .B(
        Midori_rounds_SR_Result2[44]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[44]) );
  XNOR2_X1 Midori_rounds_U370 ( .A(Midori_rounds_SR_Result2[40]), .B(
        Midori_rounds_n1740), .ZN(Midori_rounds_n1400) );
  AOI22_X1 Midori_rounds_U369 ( .A1(Midori_rounds_n1271), .A2(Key2[44]), .B1(
        Key2[108]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1740) );
  MUX2_X1 Midori_rounds_U368 ( .A(Midori_rounds_n1399), .B(
        Midori_rounds_SR_Result2[43]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[43]) );
  XNOR2_X1 Midori_rounds_U367 ( .A(Midori_rounds_SR_Result2[55]), .B(
        Midori_rounds_n1743), .ZN(Midori_rounds_n1399) );
  AOI22_X1 Midori_rounds_U366 ( .A1(Midori_rounds_n1271), .A2(Key2[43]), .B1(
        Key2[107]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1743) );
  MUX2_X1 Midori_rounds_U365 ( .A(Midori_rounds_n1398), .B(
        Midori_rounds_SR_Result2[42]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[42]) );
  XNOR2_X1 Midori_rounds_U364 ( .A(Midori_rounds_SR_Result2[54]), .B(
        Midori_rounds_n1746), .ZN(Midori_rounds_n1398) );
  AOI22_X1 Midori_rounds_U363 ( .A1(Midori_rounds_n1271), .A2(Key2[42]), .B1(
        Key2[106]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1746) );
  MUX2_X1 Midori_rounds_U362 ( .A(Midori_rounds_n1397), .B(
        Midori_rounds_SR_Result2[41]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[41]) );
  XNOR2_X1 Midori_rounds_U361 ( .A(Midori_rounds_SR_Result2[53]), .B(
        Midori_rounds_n1749), .ZN(Midori_rounds_n1397) );
  AOI22_X1 Midori_rounds_U360 ( .A1(Midori_rounds_n1271), .A2(Key2[41]), .B1(
        Key2[105]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1749) );
  MUX2_X1 Midori_rounds_U359 ( .A(Midori_rounds_n1396), .B(
        Midori_rounds_SR_Result2[40]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[40]) );
  XNOR2_X1 Midori_rounds_U358 ( .A(Midori_rounds_SR_Result2[52]), .B(
        Midori_rounds_n1752), .ZN(Midori_rounds_n1396) );
  AOI22_X1 Midori_rounds_U357 ( .A1(Midori_rounds_n1271), .A2(Key2[40]), .B1(
        Key2[104]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1752) );
  MUX2_X1 Midori_rounds_U356 ( .A(Midori_rounds_n1395), .B(
        Midori_rounds_SR_Result2[3]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[3]) );
  XNOR2_X1 Midori_rounds_U355 ( .A(Midori_rounds_SR_Result2[51]), .B(
        Midori_rounds_n1863), .ZN(Midori_rounds_n1395) );
  AOI22_X1 Midori_rounds_U354 ( .A1(Midori_rounds_n1271), .A2(Key2[3]), .B1(
        Key2[67]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1863) );
  MUX2_X1 Midori_rounds_U353 ( .A(Midori_rounds_n1394), .B(
        Midori_rounds_SR_Result2[39]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[39]) );
  XNOR2_X1 Midori_rounds_U352 ( .A(Midori_rounds_SR_Result2[19]), .B(
        Midori_rounds_n1755), .ZN(Midori_rounds_n1394) );
  AOI22_X1 Midori_rounds_U351 ( .A1(Midori_rounds_n1271), .A2(Key2[39]), .B1(
        Key2[103]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1755) );
  MUX2_X1 Midori_rounds_U350 ( .A(Midori_rounds_n1393), .B(
        Midori_rounds_SR_Result2[38]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[38]) );
  XNOR2_X1 Midori_rounds_U349 ( .A(Midori_rounds_SR_Result2[18]), .B(
        Midori_rounds_n1758), .ZN(Midori_rounds_n1393) );
  AOI22_X1 Midori_rounds_U348 ( .A1(Midori_rounds_n1271), .A2(Key2[38]), .B1(
        Key2[102]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1758) );
  MUX2_X1 Midori_rounds_U347 ( .A(Midori_rounds_n1392), .B(
        Midori_rounds_SR_Result2[37]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[37]) );
  XNOR2_X1 Midori_rounds_U346 ( .A(Midori_rounds_SR_Result2[17]), .B(
        Midori_rounds_n1761), .ZN(Midori_rounds_n1392) );
  AOI22_X1 Midori_rounds_U345 ( .A1(Midori_rounds_n1271), .A2(Key2[37]), .B1(
        Key2[101]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1761) );
  MUX2_X1 Midori_rounds_U344 ( .A(Midori_rounds_n1391), .B(
        Midori_rounds_SR_Result2[36]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[36]) );
  XNOR2_X1 Midori_rounds_U343 ( .A(Midori_rounds_SR_Result2[16]), .B(
        Midori_rounds_n1764), .ZN(Midori_rounds_n1391) );
  AOI22_X1 Midori_rounds_U342 ( .A1(Midori_rounds_n1271), .A2(Key2[36]), .B1(
        Key2[100]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1764) );
  MUX2_X1 Midori_rounds_U341 ( .A(Midori_rounds_n1390), .B(
        Midori_rounds_SR_Result2[35]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[35]) );
  XNOR2_X1 Midori_rounds_U340 ( .A(Midori_rounds_SR_Result2[15]), .B(
        Midori_rounds_n1767), .ZN(Midori_rounds_n1390) );
  AOI22_X1 Midori_rounds_U339 ( .A1(Midori_rounds_n1271), .A2(Key2[35]), .B1(
        Key2[99]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1767) );
  MUX2_X1 Midori_rounds_U338 ( .A(Midori_rounds_n1389), .B(
        Midori_rounds_SR_Result2[34]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[34]) );
  XNOR2_X1 Midori_rounds_U337 ( .A(Midori_rounds_SR_Result2[14]), .B(
        Midori_rounds_n1770), .ZN(Midori_rounds_n1389) );
  AOI22_X1 Midori_rounds_U336 ( .A1(Midori_rounds_n1271), .A2(Key2[34]), .B1(
        Key2[98]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1770) );
  MUX2_X1 Midori_rounds_U335 ( .A(Midori_rounds_n1388), .B(
        Midori_rounds_SR_Result2[33]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[33]) );
  XNOR2_X1 Midori_rounds_U334 ( .A(Midori_rounds_SR_Result2[13]), .B(
        Midori_rounds_n1773), .ZN(Midori_rounds_n1388) );
  AOI22_X1 Midori_rounds_U333 ( .A1(Midori_rounds_n1271), .A2(Key2[33]), .B1(
        Key2[97]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1773) );
  MUX2_X1 Midori_rounds_U332 ( .A(Midori_rounds_n1387), .B(
        Midori_rounds_SR_Result2[32]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[32]) );
  XNOR2_X1 Midori_rounds_U331 ( .A(Midori_rounds_SR_Result2[12]), .B(
        Midori_rounds_n1776), .ZN(Midori_rounds_n1387) );
  AOI22_X1 Midori_rounds_U330 ( .A1(Midori_rounds_n1271), .A2(Key2[32]), .B1(
        Key2[96]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1776) );
  MUX2_X1 Midori_rounds_U329 ( .A(Midori_rounds_n1386), .B(
        Midori_rounds_SR_Result2[31]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[31]) );
  XNOR2_X1 Midori_rounds_U328 ( .A(Midori_rounds_SR_Result2[3]), .B(
        Midori_rounds_n1779), .ZN(Midori_rounds_n1386) );
  AOI22_X1 Midori_rounds_U327 ( .A1(Midori_rounds_n1269), .A2(Key2[31]), .B1(
        Key2[95]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1779) );
  MUX2_X1 Midori_rounds_U326 ( .A(Midori_rounds_n1385), .B(
        Midori_rounds_SR_Result2[30]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[30]) );
  XNOR2_X1 Midori_rounds_U325 ( .A(Midori_rounds_SR_Result2[2]), .B(
        Midori_rounds_n1782), .ZN(Midori_rounds_n1385) );
  AOI22_X1 Midori_rounds_U324 ( .A1(Midori_rounds_n1273), .A2(Key2[30]), .B1(
        Key2[94]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1782) );
  MUX2_X1 Midori_rounds_U323 ( .A(Midori_rounds_n1384), .B(
        Midori_rounds_SR_Result2[2]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[2]) );
  XNOR2_X1 Midori_rounds_U322 ( .A(Midori_rounds_SR_Result2[50]), .B(
        Midori_rounds_n1866), .ZN(Midori_rounds_n1384) );
  AOI22_X1 Midori_rounds_U321 ( .A1(Midori_rounds_n1274), .A2(Key2[2]), .B1(
        Key2[66]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1866) );
  MUX2_X1 Midori_rounds_U320 ( .A(Midori_rounds_n1383), .B(
        Midori_rounds_SR_Result2[29]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[29]) );
  XNOR2_X1 Midori_rounds_U319 ( .A(Midori_rounds_SR_Result2[1]), .B(
        Midori_rounds_n1785), .ZN(Midori_rounds_n1383) );
  AOI22_X1 Midori_rounds_U318 ( .A1(Midori_rounds_n1269), .A2(Key2[29]), .B1(
        Key2[93]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1785) );
  MUX2_X1 Midori_rounds_U317 ( .A(Midori_rounds_n1382), .B(
        Midori_rounds_SR_Result2[28]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[28]) );
  XNOR2_X1 Midori_rounds_U316 ( .A(Midori_rounds_SR_Result2[0]), .B(
        Midori_rounds_n1788), .ZN(Midori_rounds_n1382) );
  AOI22_X1 Midori_rounds_U315 ( .A1(Midori_rounds_n1275), .A2(Key2[28]), .B1(
        Key2[92]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1788) );
  MUX2_X1 Midori_rounds_U314 ( .A(Midori_rounds_n1381), .B(
        Midori_rounds_SR_Result2[27]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[27]) );
  XNOR2_X1 Midori_rounds_U313 ( .A(Midori_rounds_SR_Result2[31]), .B(
        Midori_rounds_n1791), .ZN(Midori_rounds_n1381) );
  AOI22_X1 Midori_rounds_U312 ( .A1(Midori_rounds_n1273), .A2(Key2[27]), .B1(
        Key2[91]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1791) );
  MUX2_X1 Midori_rounds_U311 ( .A(Midori_rounds_n1380), .B(
        Midori_rounds_SR_Result2[26]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[26]) );
  XNOR2_X1 Midori_rounds_U310 ( .A(Midori_rounds_SR_Result2[30]), .B(
        Midori_rounds_n1794), .ZN(Midori_rounds_n1380) );
  AOI22_X1 Midori_rounds_U309 ( .A1(Midori_rounds_n1270), .A2(Key2[26]), .B1(
        Key2[90]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1794) );
  MUX2_X1 Midori_rounds_U308 ( .A(Midori_rounds_n1379), .B(
        Midori_rounds_SR_Result2[25]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[25]) );
  XNOR2_X1 Midori_rounds_U307 ( .A(Midori_rounds_SR_Result2[29]), .B(
        Midori_rounds_n1797), .ZN(Midori_rounds_n1379) );
  AOI22_X1 Midori_rounds_U306 ( .A1(Midori_rounds_n1271), .A2(Key2[25]), .B1(
        Key2[89]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1797) );
  MUX2_X1 Midori_rounds_U305 ( .A(Midori_rounds_n1378), .B(
        Midori_rounds_SR_Result2[24]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[24]) );
  XNOR2_X1 Midori_rounds_U304 ( .A(Midori_rounds_SR_Result2[28]), .B(
        Midori_rounds_n1800), .ZN(Midori_rounds_n1378) );
  AOI22_X1 Midori_rounds_U303 ( .A1(Midori_rounds_n1272), .A2(Key2[24]), .B1(
        Key2[88]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1800) );
  MUX2_X1 Midori_rounds_U302 ( .A(Midori_rounds_n1377), .B(
        Midori_rounds_SR_Result2[23]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[23]) );
  XNOR2_X1 Midori_rounds_U301 ( .A(Midori_rounds_SR_Result2[59]), .B(
        Midori_rounds_n1803), .ZN(Midori_rounds_n1377) );
  AOI22_X1 Midori_rounds_U300 ( .A1(Midori_rounds_n1274), .A2(Key2[23]), .B1(
        Key2[87]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1803) );
  MUX2_X1 Midori_rounds_U299 ( .A(Midori_rounds_n1376), .B(
        Midori_rounds_SR_Result2[22]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[22]) );
  XNOR2_X1 Midori_rounds_U298 ( .A(Midori_rounds_SR_Result2[58]), .B(
        Midori_rounds_n1806), .ZN(Midori_rounds_n1376) );
  AOI22_X1 Midori_rounds_U297 ( .A1(Midori_rounds_n1271), .A2(Key2[22]), .B1(
        Key2[86]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1806) );
  MUX2_X1 Midori_rounds_U296 ( .A(Midori_rounds_n1375), .B(
        Midori_rounds_SR_Result2[21]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[21]) );
  XNOR2_X1 Midori_rounds_U295 ( .A(Midori_rounds_SR_Result2[57]), .B(
        Midori_rounds_n1809), .ZN(Midori_rounds_n1375) );
  AOI22_X1 Midori_rounds_U294 ( .A1(Midori_rounds_n1275), .A2(Key2[21]), .B1(
        Key2[85]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1809) );
  MUX2_X1 Midori_rounds_U293 ( .A(Midori_rounds_n1374), .B(
        Midori_rounds_SR_Result2[20]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[20]) );
  XNOR2_X1 Midori_rounds_U292 ( .A(Midori_rounds_SR_Result2[56]), .B(
        Midori_rounds_n1812), .ZN(Midori_rounds_n1374) );
  AOI22_X1 Midori_rounds_U291 ( .A1(Midori_rounds_n1271), .A2(Key2[20]), .B1(
        Key2[84]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1812) );
  MUX2_X1 Midori_rounds_U290 ( .A(Midori_rounds_n1373), .B(
        Midori_rounds_SR_Result2[1]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[1]) );
  XNOR2_X1 Midori_rounds_U289 ( .A(Midori_rounds_SR_Result2[49]), .B(
        Midori_rounds_n1869), .ZN(Midori_rounds_n1373) );
  AOI22_X1 Midori_rounds_U288 ( .A1(Midori_rounds_n1271), .A2(Key2[1]), .B1(
        Key2[65]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1869) );
  MUX2_X1 Midori_rounds_U287 ( .A(Midori_rounds_n1372), .B(
        Midori_rounds_SR_Result2[19]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[19]) );
  XNOR2_X1 Midori_rounds_U286 ( .A(Midori_rounds_SR_Result2[39]), .B(
        Midori_rounds_n1815), .ZN(Midori_rounds_n1372) );
  AOI22_X1 Midori_rounds_U285 ( .A1(Midori_rounds_n1274), .A2(Key2[19]), .B1(
        Key2[83]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1815) );
  MUX2_X1 Midori_rounds_U284 ( .A(Midori_rounds_n1371), .B(
        Midori_rounds_SR_Result2[18]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[18]) );
  XNOR2_X1 Midori_rounds_U283 ( .A(Midori_rounds_SR_Result2[38]), .B(
        Midori_rounds_n1818), .ZN(Midori_rounds_n1371) );
  AOI22_X1 Midori_rounds_U282 ( .A1(Midori_rounds_n1273), .A2(Key2[18]), .B1(
        Key2[82]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1818) );
  MUX2_X1 Midori_rounds_U281 ( .A(Midori_rounds_n1370), .B(
        Midori_rounds_SR_Result2[17]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[17]) );
  XNOR2_X1 Midori_rounds_U280 ( .A(Midori_rounds_SR_Result2[37]), .B(
        Midori_rounds_n1821), .ZN(Midori_rounds_n1370) );
  AOI22_X1 Midori_rounds_U279 ( .A1(Midori_rounds_n1272), .A2(Key2[17]), .B1(
        Key2[81]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1821) );
  MUX2_X1 Midori_rounds_U278 ( .A(Midori_rounds_n1369), .B(
        Midori_rounds_SR_Result2[16]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[16]) );
  XNOR2_X1 Midori_rounds_U277 ( .A(Midori_rounds_SR_Result2[36]), .B(
        Midori_rounds_n1824), .ZN(Midori_rounds_n1369) );
  AOI22_X1 Midori_rounds_U276 ( .A1(Midori_rounds_n1274), .A2(Key2[16]), .B1(
        Key2[80]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1824) );
  MUX2_X1 Midori_rounds_U275 ( .A(Midori_rounds_n1368), .B(
        Midori_rounds_SR_Result2[15]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[15]) );
  XNOR2_X1 Midori_rounds_U274 ( .A(Midori_rounds_SR_Result2[23]), .B(
        Midori_rounds_n1827), .ZN(Midori_rounds_n1368) );
  AOI22_X1 Midori_rounds_U273 ( .A1(Midori_rounds_n1275), .A2(Key2[15]), .B1(
        Key2[79]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1827) );
  MUX2_X1 Midori_rounds_U272 ( .A(Midori_rounds_n1367), .B(
        Midori_rounds_SR_Result2[14]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[14]) );
  XNOR2_X1 Midori_rounds_U271 ( .A(Midori_rounds_SR_Result2[22]), .B(
        Midori_rounds_n1830), .ZN(Midori_rounds_n1367) );
  AOI22_X1 Midori_rounds_U270 ( .A1(Midori_rounds_n1274), .A2(Key2[14]), .B1(
        Key2[78]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1830) );
  MUX2_X1 Midori_rounds_U269 ( .A(Midori_rounds_n1366), .B(
        Midori_rounds_SR_Result2[13]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[13]) );
  XNOR2_X1 Midori_rounds_U268 ( .A(Midori_rounds_SR_Result2[21]), .B(
        Midori_rounds_n1833), .ZN(Midori_rounds_n1366) );
  AOI22_X1 Midori_rounds_U267 ( .A1(Midori_rounds_n1270), .A2(Key2[13]), .B1(
        Key2[77]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1833) );
  MUX2_X1 Midori_rounds_U266 ( .A(Midori_rounds_n1365), .B(
        Midori_rounds_SR_Result2[12]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[12]) );
  XNOR2_X1 Midori_rounds_U265 ( .A(Midori_rounds_SR_Result2[20]), .B(
        Midori_rounds_n1836), .ZN(Midori_rounds_n1365) );
  AOI22_X1 Midori_rounds_U264 ( .A1(Midori_rounds_n1272), .A2(Key2[12]), .B1(
        Key2[76]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1836) );
  MUX2_X1 Midori_rounds_U263 ( .A(Midori_rounds_n1364), .B(
        Midori_rounds_SR_Result2[11]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[11]) );
  XNOR2_X1 Midori_rounds_U262 ( .A(Midori_rounds_SR_Result2[11]), .B(
        Midori_rounds_n1839), .ZN(Midori_rounds_n1364) );
  AOI22_X1 Midori_rounds_U261 ( .A1(Midori_rounds_n1269), .A2(Key2[11]), .B1(
        Key2[75]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1839) );
  MUX2_X1 Midori_rounds_U260 ( .A(Midori_rounds_n1363), .B(
        Midori_rounds_SR_Result2[10]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[10]) );
  XNOR2_X1 Midori_rounds_U259 ( .A(Midori_rounds_SR_Result2[10]), .B(
        Midori_rounds_n1842), .ZN(Midori_rounds_n1363) );
  AOI22_X1 Midori_rounds_U258 ( .A1(Midori_rounds_n1271), .A2(Key2[10]), .B1(
        Key2[74]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1842) );
  MUX2_X1 Midori_rounds_U257 ( .A(Midori_rounds_n1362), .B(
        Midori_rounds_SR_Result2[0]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[0]) );
  XNOR2_X1 Midori_rounds_U256 ( .A(Midori_rounds_SR_Result2[48]), .B(
        Midori_rounds_n1872), .ZN(Midori_rounds_n1362) );
  AOI22_X1 Midori_rounds_U255 ( .A1(Midori_rounds_n1275), .A2(Key2[0]), .B1(
        Key2[64]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1872) );
  MUX2_X1 Midori_rounds_U254 ( .A(Midori_rounds_n1361), .B(
        Midori_rounds_SR_Result1[9]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[9]) );
  XNOR2_X1 Midori_rounds_U253 ( .A(Midori_rounds_SR_Result1[9]), .B(
        Midori_rounds_n1998), .ZN(Midori_rounds_n1361) );
  AOI22_X1 Midori_rounds_U252 ( .A1(Midori_rounds_n1270), .A2(Key1[9]), .B1(
        Key1[73]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1998) );
  MUX2_X1 Midori_rounds_U251 ( .A(Midori_rounds_n1360), .B(
        Midori_rounds_SR_Result1[8]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[8]) );
  XNOR2_X1 Midori_rounds_U250 ( .A(Midori_rounds_SR_Result1[8]), .B(
        Midori_rounds_n2058), .ZN(Midori_rounds_n1360) );
  XOR2_X1 Midori_rounds_U249 ( .A(Midori_rounds_round_Constant[2]), .B(
        Midori_rounds_n1359), .Z(Midori_rounds_n2058) );
  AOI22_X1 Midori_rounds_U248 ( .A1(Midori_rounds_n1270), .A2(Key1[8]), .B1(
        Key1[72]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1359) );
  MUX2_X1 Midori_rounds_U247 ( .A(Midori_rounds_n1358), .B(
        Midori_rounds_SR_Result1[7]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[7]) );
  XNOR2_X1 Midori_rounds_U246 ( .A(Midori_rounds_SR_Result1[47]), .B(
        Midori_rounds_n2001), .ZN(Midori_rounds_n1358) );
  AOI22_X1 Midori_rounds_U245 ( .A1(Midori_rounds_n1270), .A2(Key1[7]), .B1(
        Key1[71]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n2001) );
  MUX2_X1 Midori_rounds_U244 ( .A(Midori_rounds_n1357), .B(
        Midori_rounds_SR_Result1[6]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[6]) );
  XNOR2_X1 Midori_rounds_U243 ( .A(Midori_rounds_SR_Result1[46]), .B(
        Midori_rounds_n2004), .ZN(Midori_rounds_n1357) );
  AOI22_X1 Midori_rounds_U242 ( .A1(Midori_rounds_n1270), .A2(Key1[6]), .B1(
        Key1[70]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n2004) );
  MUX2_X1 Midori_rounds_U241 ( .A(Midori_rounds_n1356), .B(
        Midori_rounds_SR_Result1[63]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[63]) );
  XNOR2_X1 Midori_rounds_U240 ( .A(Midori_rounds_SR_Result1[63]), .B(
        Midori_rounds_n1875), .ZN(Midori_rounds_n1356) );
  AOI22_X1 Midori_rounds_U239 ( .A1(Midori_rounds_n1270), .A2(Key1[63]), .B1(
        Key1[127]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1875) );
  MUX2_X1 Midori_rounds_U238 ( .A(Midori_rounds_n1355), .B(
        Midori_rounds_SR_Result1[62]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[62]) );
  XNOR2_X1 Midori_rounds_U237 ( .A(Midori_rounds_SR_Result1[62]), .B(
        Midori_rounds_n1878), .ZN(Midori_rounds_n1355) );
  AOI22_X1 Midori_rounds_U236 ( .A1(Midori_rounds_n1270), .A2(Key1[62]), .B1(
        Key1[126]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1878) );
  MUX2_X1 Midori_rounds_U235 ( .A(Midori_rounds_n1354), .B(
        Midori_rounds_SR_Result1[61]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[61]) );
  XNOR2_X1 Midori_rounds_U234 ( .A(Midori_rounds_SR_Result1[61]), .B(
        Midori_rounds_n1881), .ZN(Midori_rounds_n1354) );
  AOI22_X1 Midori_rounds_U233 ( .A1(Midori_rounds_n1270), .A2(Key1[61]), .B1(
        Key1[125]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1881) );
  MUX2_X1 Midori_rounds_U232 ( .A(Midori_rounds_n1353), .B(
        Midori_rounds_SR_Result1[60]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[60]) );
  XNOR2_X1 Midori_rounds_U231 ( .A(Midori_rounds_SR_Result1[60]), .B(
        Midori_rounds_n2019), .ZN(Midori_rounds_n1353) );
  XOR2_X1 Midori_rounds_U230 ( .A(Midori_rounds_round_Constant[15]), .B(
        Midori_rounds_n1352), .Z(Midori_rounds_n2019) );
  AOI22_X1 Midori_rounds_U229 ( .A1(Midori_rounds_n1270), .A2(Key1[60]), .B1(
        Key1[124]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1352) );
  MUX2_X1 Midori_rounds_U228 ( .A(Midori_rounds_n1351), .B(
        Midori_rounds_SR_Result1[5]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[5]) );
  XNOR2_X1 Midori_rounds_U227 ( .A(Midori_rounds_SR_Result1[45]), .B(
        Midori_rounds_n2007), .ZN(Midori_rounds_n1351) );
  AOI22_X1 Midori_rounds_U226 ( .A1(Midori_rounds_n1270), .A2(Key1[5]), .B1(
        Key1[69]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n2007) );
  MUX2_X1 Midori_rounds_U225 ( .A(Midori_rounds_n1350), .B(
        Midori_rounds_SR_Result1[59]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[59]) );
  XNOR2_X1 Midori_rounds_U224 ( .A(Midori_rounds_SR_Result1[35]), .B(
        Midori_rounds_n1884), .ZN(Midori_rounds_n1350) );
  AOI22_X1 Midori_rounds_U223 ( .A1(Midori_rounds_n1270), .A2(Key1[59]), .B1(
        Key1[123]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1884) );
  MUX2_X1 Midori_rounds_U222 ( .A(Midori_rounds_n1349), .B(
        Midori_rounds_SR_Result1[58]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[58]) );
  XNOR2_X1 Midori_rounds_U221 ( .A(Midori_rounds_SR_Result1[34]), .B(
        Midori_rounds_n1887), .ZN(Midori_rounds_n1349) );
  AOI22_X1 Midori_rounds_U220 ( .A1(Midori_rounds_n1270), .A2(Key1[58]), .B1(
        Key1[122]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1887) );
  MUX2_X1 Midori_rounds_U219 ( .A(Midori_rounds_n1348), .B(
        Midori_rounds_SR_Result1[57]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[57]) );
  XNOR2_X1 Midori_rounds_U218 ( .A(Midori_rounds_SR_Result1[33]), .B(
        Midori_rounds_n1890), .ZN(Midori_rounds_n1348) );
  AOI22_X1 Midori_rounds_U217 ( .A1(Midori_rounds_n1270), .A2(Key1[57]), .B1(
        Key1[121]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1890) );
  MUX2_X1 Midori_rounds_U216 ( .A(Midori_rounds_n1347), .B(
        Midori_rounds_SR_Result1[56]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[56]) );
  XNOR2_X1 Midori_rounds_U215 ( .A(Midori_rounds_SR_Result1[32]), .B(
        Midori_rounds_n2022), .ZN(Midori_rounds_n1347) );
  XOR2_X1 Midori_rounds_U214 ( .A(Midori_rounds_round_Constant[14]), .B(
        Midori_rounds_n1346), .Z(Midori_rounds_n2022) );
  AOI22_X1 Midori_rounds_U213 ( .A1(Midori_rounds_n1270), .A2(Key1[56]), .B1(
        Key1[120]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1346) );
  MUX2_X1 Midori_rounds_U212 ( .A(Midori_rounds_n1345), .B(
        Midori_rounds_SR_Result1[55]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[55]) );
  XNOR2_X1 Midori_rounds_U211 ( .A(Midori_rounds_SR_Result1[7]), .B(
        Midori_rounds_n1893), .ZN(Midori_rounds_n1345) );
  AOI22_X1 Midori_rounds_U210 ( .A1(Midori_rounds_n1269), .A2(Key1[55]), .B1(
        Key1[119]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1893) );
  MUX2_X1 Midori_rounds_U209 ( .A(Midori_rounds_n1344), .B(
        Midori_rounds_SR_Result1[54]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[54]) );
  XNOR2_X1 Midori_rounds_U208 ( .A(Midori_rounds_SR_Result1[6]), .B(
        Midori_rounds_n1896), .ZN(Midori_rounds_n1344) );
  AOI22_X1 Midori_rounds_U207 ( .A1(Midori_rounds_n1269), .A2(Key1[54]), .B1(
        Key1[118]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1896) );
  MUX2_X1 Midori_rounds_U206 ( .A(Midori_rounds_n1343), .B(
        Midori_rounds_SR_Result1[53]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[53]) );
  XNOR2_X1 Midori_rounds_U205 ( .A(Midori_rounds_SR_Result1[5]), .B(
        Midori_rounds_n1899), .ZN(Midori_rounds_n1343) );
  AOI22_X1 Midori_rounds_U204 ( .A1(Midori_rounds_n1269), .A2(Key1[53]), .B1(
        Key1[117]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1899) );
  MUX2_X1 Midori_rounds_U203 ( .A(Midori_rounds_n1342), .B(
        Midori_rounds_SR_Result1[52]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[52]) );
  XNOR2_X1 Midori_rounds_U202 ( .A(Midori_rounds_SR_Result1[4]), .B(
        Midori_rounds_n2025), .ZN(Midori_rounds_n1342) );
  XOR2_X1 Midori_rounds_U201 ( .A(Midori_rounds_round_Constant[13]), .B(
        Midori_rounds_n1341), .Z(Midori_rounds_n2025) );
  AOI22_X1 Midori_rounds_U200 ( .A1(Midori_rounds_n1269), .A2(Key1[52]), .B1(
        Key1[116]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1341) );
  MUX2_X1 Midori_rounds_U199 ( .A(Midori_rounds_n1340), .B(
        Midori_rounds_SR_Result1[51]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[51]) );
  XNOR2_X1 Midori_rounds_U198 ( .A(Midori_rounds_SR_Result1[27]), .B(
        Midori_rounds_n1902), .ZN(Midori_rounds_n1340) );
  AOI22_X1 Midori_rounds_U197 ( .A1(Midori_rounds_n1269), .A2(Key1[51]), .B1(
        Key1[115]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1902) );
  MUX2_X1 Midori_rounds_U196 ( .A(Midori_rounds_n1339), .B(
        Midori_rounds_SR_Result1[50]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[50]) );
  XNOR2_X1 Midori_rounds_U195 ( .A(Midori_rounds_SR_Result1[26]), .B(
        Midori_rounds_n1905), .ZN(Midori_rounds_n1339) );
  AOI22_X1 Midori_rounds_U194 ( .A1(Midori_rounds_n1269), .A2(Key1[50]), .B1(
        Key1[114]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1905) );
  MUX2_X1 Midori_rounds_U193 ( .A(Midori_rounds_n1338), .B(
        Midori_rounds_SR_Result1[4]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[4]) );
  XNOR2_X1 Midori_rounds_U192 ( .A(Midori_rounds_SR_Result1[44]), .B(
        Midori_rounds_n2061), .ZN(Midori_rounds_n1338) );
  XOR2_X1 Midori_rounds_U191 ( .A(Midori_rounds_round_Constant[1]), .B(
        Midori_rounds_n1337), .Z(Midori_rounds_n2061) );
  AOI22_X1 Midori_rounds_U190 ( .A1(Midori_rounds_n1269), .A2(Key1[4]), .B1(
        Key1[68]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1337) );
  MUX2_X1 Midori_rounds_U189 ( .A(Midori_rounds_n1336), .B(
        Midori_rounds_SR_Result1[49]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[49]) );
  XNOR2_X1 Midori_rounds_U188 ( .A(Midori_rounds_SR_Result1[25]), .B(
        Midori_rounds_n1908), .ZN(Midori_rounds_n1336) );
  AOI22_X1 Midori_rounds_U187 ( .A1(Midori_rounds_n1269), .A2(Key1[49]), .B1(
        Key1[113]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1908) );
  MUX2_X1 Midori_rounds_U186 ( .A(Midori_rounds_n1335), .B(
        Midori_rounds_SR_Result1[48]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[48]) );
  XNOR2_X1 Midori_rounds_U185 ( .A(Midori_rounds_SR_Result1[24]), .B(
        Midori_rounds_n2028), .ZN(Midori_rounds_n1335) );
  XOR2_X1 Midori_rounds_U184 ( .A(Midori_rounds_round_Constant[12]), .B(
        Midori_rounds_n1334), .Z(Midori_rounds_n2028) );
  AOI22_X1 Midori_rounds_U183 ( .A1(Midori_rounds_n1269), .A2(Key1[48]), .B1(
        Key1[112]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1334) );
  MUX2_X1 Midori_rounds_U182 ( .A(Midori_rounds_n1333), .B(
        Midori_rounds_SR_Result1[47]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[47]) );
  XNOR2_X1 Midori_rounds_U181 ( .A(Midori_rounds_SR_Result1[43]), .B(
        Midori_rounds_n1911), .ZN(Midori_rounds_n1333) );
  AOI22_X1 Midori_rounds_U180 ( .A1(Midori_rounds_n1269), .A2(Key1[47]), .B1(
        Key1[111]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1911) );
  MUX2_X1 Midori_rounds_U179 ( .A(Midori_rounds_n1332), .B(
        Midori_rounds_SR_Result1[46]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[46]) );
  XNOR2_X1 Midori_rounds_U178 ( .A(Midori_rounds_SR_Result1[42]), .B(
        Midori_rounds_n1914), .ZN(Midori_rounds_n1332) );
  AOI22_X1 Midori_rounds_U177 ( .A1(Midori_rounds_n1269), .A2(Key1[46]), .B1(
        Key1[110]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1914) );
  MUX2_X1 Midori_rounds_U176 ( .A(Midori_rounds_n1331), .B(
        Midori_rounds_SR_Result1[45]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[45]) );
  XNOR2_X1 Midori_rounds_U175 ( .A(Midori_rounds_SR_Result1[41]), .B(
        Midori_rounds_n1917), .ZN(Midori_rounds_n1331) );
  AOI22_X1 Midori_rounds_U174 ( .A1(Midori_rounds_n1269), .A2(Key1[45]), .B1(
        Key1[109]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1917) );
  MUX2_X1 Midori_rounds_U173 ( .A(Midori_rounds_n1330), .B(
        Midori_rounds_SR_Result1[44]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[44]) );
  XNOR2_X1 Midori_rounds_U172 ( .A(Midori_rounds_SR_Result1[40]), .B(
        Midori_rounds_n2031), .ZN(Midori_rounds_n1330) );
  XOR2_X1 Midori_rounds_U171 ( .A(Midori_rounds_round_Constant[11]), .B(
        Midori_rounds_n1329), .Z(Midori_rounds_n2031) );
  AOI22_X1 Midori_rounds_U170 ( .A1(Midori_rounds_n1269), .A2(Key1[44]), .B1(
        Key1[108]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1329) );
  MUX2_X1 Midori_rounds_U169 ( .A(Midori_rounds_n1328), .B(
        Midori_rounds_SR_Result1[43]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[43]) );
  XNOR2_X1 Midori_rounds_U168 ( .A(Midori_rounds_SR_Result1[55]), .B(
        Midori_rounds_n1920), .ZN(Midori_rounds_n1328) );
  AOI22_X1 Midori_rounds_U167 ( .A1(Midori_rounds_n1268), .A2(Key1[43]), .B1(
        Key1[107]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1920) );
  MUX2_X1 Midori_rounds_U166 ( .A(Midori_rounds_n1327), .B(
        Midori_rounds_SR_Result1[42]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[42]) );
  XNOR2_X1 Midori_rounds_U165 ( .A(Midori_rounds_SR_Result1[54]), .B(
        Midori_rounds_n1923), .ZN(Midori_rounds_n1327) );
  AOI22_X1 Midori_rounds_U164 ( .A1(Midori_rounds_n1268), .A2(Key1[42]), .B1(
        Key1[106]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1923) );
  MUX2_X1 Midori_rounds_U163 ( .A(Midori_rounds_n1326), .B(
        Midori_rounds_SR_Result1[41]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[41]) );
  XNOR2_X1 Midori_rounds_U162 ( .A(Midori_rounds_SR_Result1[53]), .B(
        Midori_rounds_n1926), .ZN(Midori_rounds_n1326) );
  AOI22_X1 Midori_rounds_U161 ( .A1(Midori_rounds_n1268), .A2(Key1[41]), .B1(
        Key1[105]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1926) );
  MUX2_X1 Midori_rounds_U160 ( .A(Midori_rounds_n1325), .B(
        Midori_rounds_SR_Result1[40]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[40]) );
  XNOR2_X1 Midori_rounds_U159 ( .A(Midori_rounds_SR_Result1[52]), .B(
        Midori_rounds_n2034), .ZN(Midori_rounds_n1325) );
  XOR2_X1 Midori_rounds_U158 ( .A(Midori_rounds_round_Constant[10]), .B(
        Midori_rounds_n1324), .Z(Midori_rounds_n2034) );
  AOI22_X1 Midori_rounds_U157 ( .A1(Midori_rounds_n1268), .A2(Key1[40]), .B1(
        Key1[104]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1324) );
  MUX2_X1 Midori_rounds_U156 ( .A(Midori_rounds_n1323), .B(
        Midori_rounds_SR_Result1[3]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[3]) );
  XNOR2_X1 Midori_rounds_U155 ( .A(Midori_rounds_SR_Result1[51]), .B(
        Midori_rounds_n2010), .ZN(Midori_rounds_n1323) );
  AOI22_X1 Midori_rounds_U154 ( .A1(Midori_rounds_n1268), .A2(Key1[3]), .B1(
        Key1[67]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n2010) );
  MUX2_X1 Midori_rounds_U153 ( .A(Midori_rounds_n1322), .B(
        Midori_rounds_SR_Result1[39]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[39]) );
  XNOR2_X1 Midori_rounds_U152 ( .A(Midori_rounds_SR_Result1[19]), .B(
        Midori_rounds_n1929), .ZN(Midori_rounds_n1322) );
  AOI22_X1 Midori_rounds_U151 ( .A1(Midori_rounds_n1268), .A2(Key1[39]), .B1(
        Key1[103]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1929) );
  MUX2_X1 Midori_rounds_U150 ( .A(Midori_rounds_n1321), .B(
        Midori_rounds_SR_Result1[38]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[38]) );
  XNOR2_X1 Midori_rounds_U149 ( .A(Midori_rounds_SR_Result1[18]), .B(
        Midori_rounds_n1932), .ZN(Midori_rounds_n1321) );
  AOI22_X1 Midori_rounds_U148 ( .A1(Midori_rounds_n1268), .A2(Key1[38]), .B1(
        Key1[102]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1932) );
  MUX2_X1 Midori_rounds_U147 ( .A(Midori_rounds_n1320), .B(
        Midori_rounds_SR_Result1[37]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[37]) );
  XNOR2_X1 Midori_rounds_U146 ( .A(Midori_rounds_SR_Result1[17]), .B(
        Midori_rounds_n1935), .ZN(Midori_rounds_n1320) );
  AOI22_X1 Midori_rounds_U145 ( .A1(Midori_rounds_n1268), .A2(Key1[37]), .B1(
        Key1[101]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1935) );
  MUX2_X1 Midori_rounds_U144 ( .A(Midori_rounds_n1319), .B(
        Midori_rounds_SR_Result1[36]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[36]) );
  XNOR2_X1 Midori_rounds_U143 ( .A(Midori_rounds_SR_Result1[16]), .B(
        Midori_rounds_n2037), .ZN(Midori_rounds_n1319) );
  XOR2_X1 Midori_rounds_U142 ( .A(Midori_rounds_round_Constant[9]), .B(
        Midori_rounds_n1318), .Z(Midori_rounds_n2037) );
  AOI22_X1 Midori_rounds_U141 ( .A1(Midori_rounds_n1268), .A2(Key1[36]), .B1(
        Key1[100]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1318) );
  MUX2_X1 Midori_rounds_U140 ( .A(Midori_rounds_n1317), .B(
        Midori_rounds_SR_Result1[35]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[35]) );
  XNOR2_X1 Midori_rounds_U139 ( .A(Midori_rounds_SR_Result1[15]), .B(
        Midori_rounds_n1938), .ZN(Midori_rounds_n1317) );
  AOI22_X1 Midori_rounds_U138 ( .A1(Midori_rounds_n1268), .A2(Key1[35]), .B1(
        Key1[99]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1938) );
  MUX2_X1 Midori_rounds_U137 ( .A(Midori_rounds_n1316), .B(
        Midori_rounds_SR_Result1[34]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[34]) );
  XNOR2_X1 Midori_rounds_U136 ( .A(Midori_rounds_SR_Result1[14]), .B(
        Midori_rounds_n1941), .ZN(Midori_rounds_n1316) );
  AOI22_X1 Midori_rounds_U135 ( .A1(Midori_rounds_n1268), .A2(Key1[34]), .B1(
        Key1[98]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1941) );
  MUX2_X1 Midori_rounds_U134 ( .A(Midori_rounds_n1315), .B(
        Midori_rounds_SR_Result1[33]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[33]) );
  XNOR2_X1 Midori_rounds_U133 ( .A(Midori_rounds_SR_Result1[13]), .B(
        Midori_rounds_n1944), .ZN(Midori_rounds_n1315) );
  AOI22_X1 Midori_rounds_U132 ( .A1(Midori_rounds_n1268), .A2(Key1[33]), .B1(
        Key1[97]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1944) );
  MUX2_X1 Midori_rounds_U131 ( .A(Midori_rounds_n1314), .B(
        Midori_rounds_SR_Result1[32]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[32]) );
  XNOR2_X1 Midori_rounds_U130 ( .A(Midori_rounds_SR_Result1[12]), .B(
        Midori_rounds_n2040), .ZN(Midori_rounds_n1314) );
  XOR2_X1 Midori_rounds_U129 ( .A(Midori_rounds_round_Constant[8]), .B(
        Midori_rounds_n1313), .Z(Midori_rounds_n2040) );
  AOI22_X1 Midori_rounds_U128 ( .A1(Midori_rounds_n1268), .A2(Key1[32]), .B1(
        Key1[96]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1313) );
  MUX2_X1 Midori_rounds_U127 ( .A(Midori_rounds_n1312), .B(
        Midori_rounds_SR_Result1[31]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[31]) );
  XNOR2_X1 Midori_rounds_U126 ( .A(Midori_rounds_SR_Result1[3]), .B(
        Midori_rounds_n1947), .ZN(Midori_rounds_n1312) );
  AOI22_X1 Midori_rounds_U125 ( .A1(Midori_rounds_n1268), .A2(Key1[31]), .B1(
        Key1[95]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1947) );
  MUX2_X1 Midori_rounds_U124 ( .A(Midori_rounds_n1311), .B(
        Midori_rounds_SR_Result1[30]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[30]) );
  XNOR2_X1 Midori_rounds_U123 ( .A(Midori_rounds_SR_Result1[2]), .B(
        Midori_rounds_n1950), .ZN(Midori_rounds_n1311) );
  AOI22_X1 Midori_rounds_U122 ( .A1(Midori_rounds_n1268), .A2(Key1[30]), .B1(
        Key1[94]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1950) );
  MUX2_X1 Midori_rounds_U121 ( .A(Midori_rounds_n1310), .B(
        Midori_rounds_SR_Result1[2]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[2]) );
  XNOR2_X1 Midori_rounds_U120 ( .A(Midori_rounds_SR_Result1[50]), .B(
        Midori_rounds_n2013), .ZN(Midori_rounds_n1310) );
  AOI22_X1 Midori_rounds_U119 ( .A1(Midori_rounds_n1267), .A2(Key1[2]), .B1(
        Key1[66]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n2013) );
  MUX2_X1 Midori_rounds_U118 ( .A(Midori_rounds_n1309), .B(
        Midori_rounds_SR_Result1[29]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[29]) );
  XNOR2_X1 Midori_rounds_U117 ( .A(Midori_rounds_SR_Result1[1]), .B(
        Midori_rounds_n1953), .ZN(Midori_rounds_n1309) );
  AOI22_X1 Midori_rounds_U116 ( .A1(Midori_rounds_n1267), .A2(Key1[29]), .B1(
        Key1[93]), .B2(Midori_rounds_n1282), .ZN(Midori_rounds_n1953) );
  MUX2_X1 Midori_rounds_U115 ( .A(Midori_rounds_n1308), .B(
        Midori_rounds_SR_Result1[28]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[28]) );
  XNOR2_X1 Midori_rounds_U114 ( .A(Midori_rounds_SR_Result1[0]), .B(
        Midori_rounds_n2043), .ZN(Midori_rounds_n1308) );
  XOR2_X1 Midori_rounds_U113 ( .A(Midori_rounds_round_Constant[7]), .B(
        Midori_rounds_n1307), .Z(Midori_rounds_n2043) );
  AOI22_X1 Midori_rounds_U112 ( .A1(Midori_rounds_n1268), .A2(Key1[28]), .B1(
        Key1[92]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1307) );
  MUX2_X1 Midori_rounds_U111 ( .A(Midori_rounds_n1306), .B(
        Midori_rounds_SR_Result1[27]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[27]) );
  XNOR2_X1 Midori_rounds_U110 ( .A(Midori_rounds_SR_Result1[31]), .B(
        Midori_rounds_n1956), .ZN(Midori_rounds_n1306) );
  AOI22_X1 Midori_rounds_U109 ( .A1(Midori_rounds_n1268), .A2(Key1[27]), .B1(
        Key1[91]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1956) );
  MUX2_X1 Midori_rounds_U108 ( .A(Midori_rounds_n1305), .B(
        Midori_rounds_SR_Result1[26]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[26]) );
  XNOR2_X1 Midori_rounds_U107 ( .A(Midori_rounds_SR_Result1[30]), .B(
        Midori_rounds_n1959), .ZN(Midori_rounds_n1305) );
  AOI22_X1 Midori_rounds_U106 ( .A1(Midori_rounds_n1268), .A2(Key1[26]), .B1(
        Key1[90]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1959) );
  MUX2_X1 Midori_rounds_U105 ( .A(Midori_rounds_n1304), .B(
        Midori_rounds_SR_Result1[25]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[25]) );
  XNOR2_X1 Midori_rounds_U104 ( .A(Midori_rounds_SR_Result1[29]), .B(
        Midori_rounds_n1962), .ZN(Midori_rounds_n1304) );
  AOI22_X1 Midori_rounds_U103 ( .A1(Midori_rounds_n1267), .A2(Key1[25]), .B1(
        Key1[89]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1962) );
  MUX2_X1 Midori_rounds_U102 ( .A(Midori_rounds_n1303), .B(
        Midori_rounds_SR_Result1[24]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[24]) );
  XNOR2_X1 Midori_rounds_U101 ( .A(Midori_rounds_SR_Result1[28]), .B(
        Midori_rounds_n2046), .ZN(Midori_rounds_n1303) );
  XOR2_X1 Midori_rounds_U100 ( .A(Midori_rounds_round_Constant[6]), .B(
        Midori_rounds_n1302), .Z(Midori_rounds_n2046) );
  AOI22_X1 Midori_rounds_U99 ( .A1(Midori_rounds_n1268), .A2(Key1[24]), .B1(
        Key1[88]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1302) );
  MUX2_X1 Midori_rounds_U98 ( .A(Midori_rounds_n1301), .B(
        Midori_rounds_SR_Result1[23]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[23]) );
  XNOR2_X1 Midori_rounds_U97 ( .A(Midori_rounds_SR_Result1[59]), .B(
        Midori_rounds_n1965), .ZN(Midori_rounds_n1301) );
  AOI22_X1 Midori_rounds_U96 ( .A1(Midori_rounds_n1268), .A2(Key1[23]), .B1(
        Key1[87]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1965) );
  MUX2_X1 Midori_rounds_U95 ( .A(Midori_rounds_n1300), .B(
        Midori_rounds_SR_Result1[22]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[22]) );
  XNOR2_X1 Midori_rounds_U94 ( .A(Midori_rounds_SR_Result1[58]), .B(
        Midori_rounds_n1968), .ZN(Midori_rounds_n1300) );
  AOI22_X1 Midori_rounds_U93 ( .A1(Midori_rounds_n1268), .A2(Key1[22]), .B1(
        Key1[86]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1968) );
  MUX2_X1 Midori_rounds_U92 ( .A(Midori_rounds_n1299), .B(
        Midori_rounds_SR_Result1[21]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[21]) );
  XNOR2_X1 Midori_rounds_U91 ( .A(Midori_rounds_SR_Result1[57]), .B(
        Midori_rounds_n1971), .ZN(Midori_rounds_n1299) );
  AOI22_X1 Midori_rounds_U90 ( .A1(Midori_rounds_n1267), .A2(Key1[21]), .B1(
        Key1[85]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1971) );
  MUX2_X1 Midori_rounds_U89 ( .A(Midori_rounds_n1298), .B(
        Midori_rounds_SR_Result1[20]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[20]) );
  XNOR2_X1 Midori_rounds_U88 ( .A(Midori_rounds_SR_Result1[56]), .B(
        Midori_rounds_n2049), .ZN(Midori_rounds_n1298) );
  MUX2_X1 Midori_rounds_U87 ( .A(Midori_rounds_n1297), .B(
        Midori_rounds_SR_Result1[1]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[1]) );
  XNOR2_X1 Midori_rounds_U86 ( .A(Midori_rounds_SR_Result1[49]), .B(
        Midori_rounds_n2016), .ZN(Midori_rounds_n1297) );
  AOI22_X1 Midori_rounds_U85 ( .A1(Midori_rounds_n1267), .A2(Key1[1]), .B1(
        Key1[65]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n2016) );
  MUX2_X1 Midori_rounds_U84 ( .A(Midori_rounds_n1296), .B(
        Midori_rounds_SR_Result1[19]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[19]) );
  XNOR2_X1 Midori_rounds_U83 ( .A(Midori_rounds_SR_Result1[39]), .B(
        Midori_rounds_n1974), .ZN(Midori_rounds_n1296) );
  AOI22_X1 Midori_rounds_U82 ( .A1(Midori_rounds_n1267), .A2(Key1[19]), .B1(
        Key1[83]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1974) );
  MUX2_X1 Midori_rounds_U81 ( .A(Midori_rounds_n1295), .B(
        Midori_rounds_SR_Result1[18]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[18]) );
  XNOR2_X1 Midori_rounds_U80 ( .A(Midori_rounds_SR_Result1[38]), .B(
        Midori_rounds_n1977), .ZN(Midori_rounds_n1295) );
  AOI22_X1 Midori_rounds_U79 ( .A1(Midori_rounds_n1267), .A2(Key1[18]), .B1(
        Key1[82]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1977) );
  MUX2_X1 Midori_rounds_U78 ( .A(Midori_rounds_n1294), .B(
        Midori_rounds_SR_Result1[17]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[17]) );
  XNOR2_X1 Midori_rounds_U77 ( .A(Midori_rounds_SR_Result1[37]), .B(
        Midori_rounds_n1980), .ZN(Midori_rounds_n1294) );
  AOI22_X1 Midori_rounds_U76 ( .A1(Midori_rounds_n1267), .A2(Key1[17]), .B1(
        Key1[81]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1980) );
  MUX2_X1 Midori_rounds_U75 ( .A(Midori_rounds_n1293), .B(
        Midori_rounds_SR_Result1[16]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[16]) );
  XNOR2_X1 Midori_rounds_U74 ( .A(Midori_rounds_SR_Result1[36]), .B(
        Midori_rounds_n2052), .ZN(Midori_rounds_n1293) );
  XOR2_X1 Midori_rounds_U73 ( .A(Midori_rounds_round_Constant[4]), .B(
        Midori_rounds_n1292), .Z(Midori_rounds_n2052) );
  AOI22_X1 Midori_rounds_U72 ( .A1(Midori_rounds_n1267), .A2(Key1[16]), .B1(
        Key1[80]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1292) );
  MUX2_X1 Midori_rounds_U71 ( .A(Midori_rounds_n1291), .B(
        Midori_rounds_SR_Result1[15]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[15]) );
  XNOR2_X1 Midori_rounds_U70 ( .A(Midori_rounds_SR_Result1[23]), .B(
        Midori_rounds_n1983), .ZN(Midori_rounds_n1291) );
  AOI22_X1 Midori_rounds_U69 ( .A1(Midori_rounds_n1267), .A2(Key1[15]), .B1(
        Key1[79]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1983) );
  MUX2_X1 Midori_rounds_U68 ( .A(Midori_rounds_n1290), .B(
        Midori_rounds_SR_Result1[14]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[14]) );
  XNOR2_X1 Midori_rounds_U67 ( .A(Midori_rounds_SR_Result1[22]), .B(
        Midori_rounds_n1986), .ZN(Midori_rounds_n1290) );
  AOI22_X1 Midori_rounds_U66 ( .A1(Midori_rounds_n1267), .A2(Key1[14]), .B1(
        Key1[78]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1986) );
  MUX2_X1 Midori_rounds_U65 ( .A(Midori_rounds_n1289), .B(
        Midori_rounds_SR_Result1[13]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[13]) );
  XNOR2_X1 Midori_rounds_U64 ( .A(Midori_rounds_SR_Result1[21]), .B(
        Midori_rounds_n1989), .ZN(Midori_rounds_n1289) );
  AOI22_X1 Midori_rounds_U63 ( .A1(Midori_rounds_n1267), .A2(Key1[13]), .B1(
        Key1[77]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1989) );
  MUX2_X1 Midori_rounds_U62 ( .A(Midori_rounds_n1288), .B(
        Midori_rounds_SR_Result1[12]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[12]) );
  XNOR2_X1 Midori_rounds_U61 ( .A(Midori_rounds_SR_Result1[20]), .B(
        Midori_rounds_n2055), .ZN(Midori_rounds_n1288) );
  XOR2_X1 Midori_rounds_U60 ( .A(Midori_rounds_round_Constant[3]), .B(
        Midori_rounds_n1287), .Z(Midori_rounds_n2055) );
  AOI22_X1 Midori_rounds_U59 ( .A1(Midori_rounds_n1267), .A2(Key1[12]), .B1(
        Key1[76]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1287) );
  MUX2_X1 Midori_rounds_U58 ( .A(Midori_rounds_n1286), .B(
        Midori_rounds_SR_Result1[11]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[11]) );
  XNOR2_X1 Midori_rounds_U57 ( .A(Midori_rounds_SR_Result1[11]), .B(
        Midori_rounds_n1992), .ZN(Midori_rounds_n1286) );
  AOI22_X1 Midori_rounds_U56 ( .A1(Midori_rounds_n1267), .A2(Key1[11]), .B1(
        Key1[75]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1992) );
  MUX2_X1 Midori_rounds_U55 ( .A(Midori_rounds_n1285), .B(
        Midori_rounds_SR_Result1[10]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[10]) );
  XNOR2_X1 Midori_rounds_U54 ( .A(Midori_rounds_SR_Result1[10]), .B(
        Midori_rounds_n1995), .ZN(Midori_rounds_n1285) );
  AOI22_X1 Midori_rounds_U53 ( .A1(Midori_rounds_n1267), .A2(Key1[10]), .B1(
        Key1[74]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1995) );
  MUX2_X1 Midori_rounds_U52 ( .A(Midori_rounds_n1284), .B(
        Midori_rounds_SR_Result1[0]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[0]) );
  XNOR2_X1 Midori_rounds_U51 ( .A(Midori_rounds_SR_Result1[48]), .B(
        Midori_rounds_n2064), .ZN(Midori_rounds_n1284) );
  XOR2_X1 Midori_rounds_U50 ( .A(Midori_rounds_round_Constant[0]), .B(
        Midori_rounds_n1283), .Z(Midori_rounds_n2064) );
  AOI22_X1 Midori_rounds_U49 ( .A1(Midori_rounds_n1267), .A2(Key1[0]), .B1(
        Key1[64]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1283) );
  INV_X1 Midori_rounds_U48 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1269)
         );
  INV_X1 Midori_rounds_U47 ( .A(enc_dec), .ZN(Midori_rounds_n1491) );
  BUF_X1 Midori_rounds_U46 ( .A(Midori_rounds_n1491), .Z(Midori_rounds_n1247)
         );
  BUF_X1 Midori_rounds_U45 ( .A(Midori_rounds_n1247), .Z(Midori_rounds_n1243)
         );
  BUF_X1 Midori_rounds_U44 ( .A(Midori_rounds_n1243), .Z(Midori_rounds_n1249)
         );
  INV_X1 Midori_rounds_U43 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1270)
         );
  BUF_X1 Midori_rounds_U42 ( .A(Midori_rounds_n1276), .Z(Midori_rounds_n1280)
         );
  BUF_X2 Midori_rounds_U41 ( .A(Midori_rounds_n2067), .Z(Midori_rounds_n1265)
         );
  BUF_X1 Midori_rounds_U40 ( .A(Midori_rounds_n1491), .Z(Midori_rounds_n1246)
         );
  NOR2_X1 Midori_rounds_U39 ( .A1(reset), .A2(Midori_rounds_n1246), .ZN(
        Midori_rounds_n2065) );
  BUF_X1 Midori_rounds_U38 ( .A(Midori_rounds_n1247), .Z(Midori_rounds_n1242)
         );
  BUF_X1 Midori_rounds_U37 ( .A(Midori_rounds_n1242), .Z(Midori_rounds_n1248)
         );
  BUF_X1 Midori_rounds_U36 ( .A(Midori_rounds_n2067), .Z(Midori_rounds_n1262)
         );
  BUF_X1 Midori_rounds_U35 ( .A(Midori_rounds_n2065), .Z(Midori_rounds_n1258)
         );
  BUF_X1 Midori_rounds_U34 ( .A(Midori_rounds_n1258), .Z(Midori_rounds_n1252)
         );
  INV_X1 Midori_rounds_U33 ( .A(Midori_rounds_n1277), .ZN(Midori_rounds_n1268)
         );
  BUF_X1 Midori_rounds_U32 ( .A(Midori_rounds_n2065), .Z(Midori_rounds_n1257)
         );
  BUF_X1 Midori_rounds_U31 ( .A(Midori_rounds_n1257), .Z(Midori_rounds_n1251)
         );
  BUF_X1 Midori_rounds_U30 ( .A(Midori_rounds_n2065), .Z(Midori_rounds_n1255)
         );
  BUF_X1 Midori_rounds_U29 ( .A(Midori_rounds_n2065), .Z(Midori_rounds_n1254)
         );
  BUF_X1 Midori_rounds_U28 ( .A(Midori_rounds_n2067), .Z(Midori_rounds_n1266)
         );
  BUF_X1 Midori_rounds_U27 ( .A(Midori_rounds_n1257), .Z(Midori_rounds_n1253)
         );
  BUF_X1 Midori_rounds_U26 ( .A(Midori_rounds_n2067), .Z(Midori_rounds_n1264)
         );
  BUF_X1 Midori_rounds_U25 ( .A(Midori_rounds_n2065), .Z(Midori_rounds_n1256)
         );
  BUF_X1 Midori_rounds_U24 ( .A(Midori_rounds_n1256), .Z(Midori_rounds_n1259)
         );
  BUF_X1 Midori_rounds_U23 ( .A(Midori_rounds_n2067), .Z(Midori_rounds_n1263)
         );
  INV_X1 Midori_rounds_U22 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1271)
         );
  INV_X1 Midori_rounds_U21 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1272)
         );
  BUF_X1 Midori_rounds_U20 ( .A(Midori_rounds_n1247), .Z(Midori_rounds_n1244)
         );
  INV_X1 Midori_rounds_U19 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1273)
         );
  BUF_X1 Midori_rounds_U18 ( .A(Midori_rounds_n1282), .Z(Midori_rounds_n1281)
         );
  BUF_X1 Midori_rounds_U17 ( .A(Midori_rounds_n1246), .Z(Midori_rounds_n1245)
         );
  BUF_X1 Midori_rounds_U16 ( .A(Midori_rounds_n1491), .Z(Midori_rounds_n1250)
         );
  BUF_X1 Midori_rounds_U15 ( .A(Midori_rounds_n1262), .Z(Midori_rounds_n1260)
         );
  BUF_X1 Midori_rounds_U14 ( .A(Midori_rounds_n1265), .Z(Midori_rounds_n1261)
         );
  BUF_X1 Midori_rounds_U13 ( .A(Midori_rounds_n1282), .Z(Midori_rounds_n1277)
         );
  INV_X1 Midori_rounds_U12 ( .A(Midori_rounds_n1277), .ZN(Midori_rounds_n1267)
         );
  BUF_X1 Midori_rounds_U11 ( .A(Midori_rounds_n1282), .Z(Midori_rounds_n1278)
         );
  BUF_X1 Midori_rounds_U10 ( .A(Midori_rounds_n1278), .Z(Midori_rounds_n1279)
         );
  OR2_X1 Midori_rounds_U9 ( .A1(enc_dec), .A2(reset), .ZN(Midori_rounds_n2067)
         );
  INV_X1 Midori_rounds_U8 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1275)
         );
  INV_X1 Midori_rounds_U7 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1274)
         );
  BUF_X1 Midori_rounds_U6 ( .A(Midori_rounds_n1282), .Z(Midori_rounds_n1276)
         );
  INV_X4 Midori_rounds_U5 ( .A(round_Signal[0]), .ZN(Midori_rounds_n1282) );
  XOR2_X1 Midori_rounds_U4 ( .A(Midori_rounds_n1241), .B(
        Midori_rounds_round_Constant[5]), .Z(Midori_rounds_n2049) );
  AOI22_X1 Midori_rounds_U3 ( .A1(Midori_rounds_n1278), .A2(Key1[84]), .B1(
        Key1[20]), .B2(Midori_rounds_n1268), .ZN(Midori_rounds_n1241) );
  NAND3_X1 Midori_rounds_constant_MUX_U77 ( .A1(Midori_rounds_constant_MUX_n70), .A2(Midori_rounds_constant_MUX_n69), .A3(Midori_rounds_constant_MUX_n68), 
        .ZN(Midori_rounds_round_Constant[9]) );
  INV_X1 Midori_rounds_constant_MUX_U76 ( .A(Midori_rounds_constant_MUX_n67), 
        .ZN(Midori_rounds_constant_MUX_n70) );
  OR3_X1 Midori_rounds_constant_MUX_U75 ( .A1(Midori_rounds_constant_MUX_n66), 
        .A2(Midori_rounds_constant_MUX_n65), .A3(
        Midori_rounds_constant_MUX_n64), .ZN(Midori_rounds_round_Constant[8])
         );
  NAND4_X1 Midori_rounds_constant_MUX_U74 ( .A1(Midori_rounds_constant_MUX_n63), .A2(Midori_rounds_constant_MUX_n62), .A3(Midori_rounds_constant_MUX_n61), 
        .A4(Midori_rounds_constant_MUX_n60), .ZN(
        Midori_rounds_round_Constant[7]) );
  NAND3_X1 Midori_rounds_constant_MUX_U73 ( .A1(Midori_rounds_constant_MUX_n59), .A2(Midori_rounds_constant_MUX_n58), .A3(Midori_rounds_constant_MUX_n69), 
        .ZN(Midori_rounds_round_Constant[6]) );
  NAND2_X1 Midori_rounds_constant_MUX_U72 ( .A1(Midori_rounds_constant_MUX_n54), .A2(Midori_rounds_constant_MUX_n55), .ZN(Midori_rounds_round_Constant[4]) );
  NOR3_X1 Midori_rounds_constant_MUX_U71 ( .A1(Midori_rounds_constant_MUX_n53), 
        .A2(Midori_rounds_constant_MUX_n66), .A3(
        Midori_rounds_constant_MUX_n52), .ZN(Midori_rounds_constant_MUX_n55)
         );
  NAND2_X1 Midori_rounds_constant_MUX_U70 ( .A1(Midori_rounds_constant_MUX_n51), .A2(Midori_rounds_constant_MUX_n50), .ZN(Midori_rounds_round_Constant[3]) );
  NOR4_X1 Midori_rounds_constant_MUX_U69 ( .A1(Midori_rounds_constant_MUX_n49), 
        .A2(Midori_rounds_constant_MUX_n64), .A3(
        Midori_rounds_constant_MUX_n48), .A4(Midori_rounds_constant_MUX_n53), 
        .ZN(Midori_rounds_constant_MUX_n50) );
  NAND3_X1 Midori_rounds_constant_MUX_U68 ( .A1(Midori_rounds_constant_MUX_n61), .A2(Midori_rounds_constant_MUX_n47), .A3(Midori_rounds_constant_MUX_n69), 
        .ZN(Midori_rounds_round_Constant[2]) );
  NOR2_X1 Midori_rounds_constant_MUX_U67 ( .A1(Midori_rounds_constant_MUX_n64), 
        .A2(Midori_rounds_constant_MUX_n56), .ZN(
        Midori_rounds_constant_MUX_n69) );
  NAND4_X1 Midori_rounds_constant_MUX_U66 ( .A1(Midori_rounds_constant_MUX_n51), .A2(Midori_rounds_constant_MUX_n46), .A3(Midori_rounds_constant_MUX_n61), 
        .A4(Midori_rounds_constant_MUX_n45), .ZN(
        Midori_rounds_round_Constant[1]) );
  NOR3_X1 Midori_rounds_constant_MUX_U65 ( .A1(Midori_rounds_constant_MUX_n44), 
        .A2(Midori_rounds_constant_MUX_n48), .A3(
        Midori_rounds_constant_MUX_n56), .ZN(Midori_rounds_constant_MUX_n45)
         );
  OAI22_X1 Midori_rounds_constant_MUX_U64 ( .A1(Midori_rounds_constant_MUX_n43), .A2(Midori_rounds_constant_MUX_n42), .B1(Midori_rounds_constant_MUX_n41), 
        .B2(Midori_rounds_constant_MUX_n40), .ZN(
        Midori_rounds_constant_MUX_n56) );
  NAND3_X1 Midori_rounds_constant_MUX_U63 ( .A1(Midori_rounds_constant_MUX_n51), .A2(Midori_rounds_constant_MUX_n59), .A3(Midori_rounds_constant_MUX_n39), 
        .ZN(Midori_rounds_round_Constant[15]) );
  NAND3_X1 Midori_rounds_constant_MUX_U62 ( .A1(Midori_rounds_constant_MUX_n63), .A2(Midori_rounds_constant_MUX_n38), .A3(Midori_rounds_constant_MUX_n54), 
        .ZN(Midori_rounds_round_Constant[14]) );
  NOR2_X1 Midori_rounds_constant_MUX_U61 ( .A1(Midori_rounds_constant_MUX_n44), 
        .A2(Midori_rounds_constant_MUX_n65), .ZN(
        Midori_rounds_constant_MUX_n54) );
  INV_X1 Midori_rounds_constant_MUX_U60 ( .A(Midori_rounds_constant_MUX_n37), 
        .ZN(Midori_rounds_constant_MUX_n65) );
  INV_X1 Midori_rounds_constant_MUX_U59 ( .A(Midori_rounds_constant_MUX_n53), 
        .ZN(Midori_rounds_constant_MUX_n63) );
  OAI22_X1 Midori_rounds_constant_MUX_U58 ( .A1(Midori_rounds_constant_MUX_n36), .A2(Midori_rounds_constant_MUX_n35), .B1(Midori_rounds_constant_MUX_n34), 
        .B2(Midori_rounds_constant_MUX_n33), .ZN(
        Midori_rounds_constant_MUX_n53) );
  NAND4_X1 Midori_rounds_constant_MUX_U57 ( .A1(Midori_rounds_constant_MUX_n38), .A2(Midori_rounds_constant_MUX_n32), .A3(Midori_rounds_constant_MUX_n61), 
        .A4(Midori_rounds_constant_MUX_n31), .ZN(
        Midori_rounds_round_Constant[13]) );
  NOR2_X1 Midori_rounds_constant_MUX_U56 ( .A1(Midori_rounds_constant_MUX_n49), 
        .A2(Midori_rounds_constant_MUX_n30), .ZN(
        Midori_rounds_constant_MUX_n61) );
  AOI21_X1 Midori_rounds_constant_MUX_U55 ( .B1(Midori_rounds_constant_MUX_n29), .B2(Midori_rounds_constant_MUX_n28), .A(Midori_rounds_constant_MUX_n34), 
        .ZN(Midori_rounds_constant_MUX_n49) );
  INV_X1 Midori_rounds_constant_MUX_U54 ( .A(Midori_rounds_constant_MUX_n52), 
        .ZN(Midori_rounds_constant_MUX_n32) );
  INV_X1 Midori_rounds_constant_MUX_U53 ( .A(Midori_rounds_constant_MUX_n27), 
        .ZN(Midori_rounds_constant_MUX_n38) );
  NAND3_X1 Midori_rounds_constant_MUX_U52 ( .A1(Midori_rounds_constant_MUX_n37), .A2(Midori_rounds_constant_MUX_n62), .A3(Midori_rounds_constant_MUX_n58), 
        .ZN(Midori_rounds_round_Constant[12]) );
  NOR2_X1 Midori_rounds_constant_MUX_U51 ( .A1(Midori_rounds_constant_MUX_n27), 
        .A2(Midori_rounds_constant_MUX_n48), .ZN(
        Midori_rounds_constant_MUX_n58) );
  NOR3_X1 Midori_rounds_constant_MUX_U50 ( .A1(Midori_rounds_constant_MUX_n67), 
        .A2(Midori_rounds_constant_MUX_n57), .A3(
        Midori_rounds_constant_MUX_n30), .ZN(Midori_rounds_constant_MUX_n37)
         );
  OAI211_X1 Midori_rounds_constant_MUX_U49 ( .C1(
        Midori_rounds_constant_MUX_n33), .C2(Midori_rounds_constant_MUX_n41), 
        .A(Midori_rounds_constant_MUX_n26), .B(Midori_rounds_constant_MUX_n59), 
        .ZN(Midori_rounds_constant_MUX_n57) );
  INV_X1 Midori_rounds_constant_MUX_U48 ( .A(Midori_rounds_constant_MUX_n25), 
        .ZN(Midori_rounds_constant_MUX_n59) );
  OAI22_X1 Midori_rounds_constant_MUX_U47 ( .A1(Midori_rounds_constant_MUX_n36), .A2(Midori_rounds_constant_MUX_n24), .B1(Midori_rounds_constant_MUX_n34), 
        .B2(Midori_rounds_constant_MUX_n43), .ZN(
        Midori_rounds_constant_MUX_n25) );
  OR2_X1 Midori_rounds_constant_MUX_U46 ( .A1(Midori_rounds_constant_MUX_n42), 
        .A2(Midori_rounds_constant_MUX_n28), .ZN(
        Midori_rounds_constant_MUX_n26) );
  INV_X1 Midori_rounds_constant_MUX_U45 ( .A(Midori_rounds_constant_MUX_n60), 
        .ZN(Midori_rounds_round_Constant[11]) );
  NOR3_X1 Midori_rounds_constant_MUX_U44 ( .A1(Midori_rounds_constant_MUX_n67), 
        .A2(Midori_rounds_constant_MUX_n27), .A3(
        Midori_rounds_constant_MUX_n64), .ZN(Midori_rounds_constant_MUX_n60)
         );
  NOR3_X1 Midori_rounds_constant_MUX_U43 ( .A1(Midori_rounds_constant_MUX_n36), 
        .A2(Midori_rounds_constant_MUX_n23), .A3(round_Signal[3]), .ZN(
        Midori_rounds_constant_MUX_n64) );
  OAI211_X1 Midori_rounds_constant_MUX_U42 ( .C1(
        Midori_rounds_constant_MUX_n34), .C2(Midori_rounds_constant_MUX_n24), 
        .A(Midori_rounds_constant_MUX_n22), .B(Midori_rounds_constant_MUX_n51), 
        .ZN(Midori_rounds_constant_MUX_n27) );
  INV_X1 Midori_rounds_constant_MUX_U41 ( .A(Midori_rounds_constant_MUX_n21), 
        .ZN(Midori_rounds_constant_MUX_n51) );
  OAI22_X1 Midori_rounds_constant_MUX_U40 ( .A1(Midori_rounds_constant_MUX_n36), .A2(Midori_rounds_constant_MUX_n33), .B1(Midori_rounds_constant_MUX_n35), 
        .B2(Midori_rounds_constant_MUX_n34), .ZN(
        Midori_rounds_constant_MUX_n21) );
  OR2_X1 Midori_rounds_constant_MUX_U39 ( .A1(Midori_rounds_constant_MUX_n36), 
        .A2(Midori_rounds_constant_MUX_n43), .ZN(
        Midori_rounds_constant_MUX_n22) );
  NAND2_X1 Midori_rounds_constant_MUX_U38 ( .A1(round_Signal[2]), .A2(
        Midori_rounds_n1267), .ZN(Midori_rounds_constant_MUX_n36) );
  NAND2_X1 Midori_rounds_constant_MUX_U37 ( .A1(Midori_rounds_constant_MUX_n46), .A2(Midori_rounds_constant_MUX_n39), .ZN(Midori_rounds_round_Constant[10])
         );
  NOR3_X1 Midori_rounds_constant_MUX_U36 ( .A1(Midori_rounds_constant_MUX_n67), 
        .A2(Midori_rounds_constant_MUX_n52), .A3(
        Midori_rounds_constant_MUX_n20), .ZN(Midori_rounds_constant_MUX_n39)
         );
  OAI21_X1 Midori_rounds_constant_MUX_U35 ( .B1(Midori_rounds_constant_MUX_n35), .B2(Midori_rounds_constant_MUX_n42), .A(Midori_rounds_constant_MUX_n19), 
        .ZN(Midori_rounds_constant_MUX_n67) );
  OAI211_X1 Midori_rounds_constant_MUX_U34 ( .C1(
        Midori_rounds_constant_MUX_n18), .C2(Midori_rounds_n1267), .A(
        round_Signal[2]), .B(Midori_rounds_constant_MUX_n17), .ZN(
        Midori_rounds_constant_MUX_n19) );
  INV_X1 Midori_rounds_constant_MUX_U33 ( .A(Midori_rounds_constant_MUX_n66), 
        .ZN(Midori_rounds_constant_MUX_n46) );
  NAND4_X1 Midori_rounds_constant_MUX_U32 ( .A1(Midori_rounds_constant_MUX_n16), .A2(Midori_rounds_constant_MUX_n62), .A3(Midori_rounds_constant_MUX_n47), 
        .A4(Midori_rounds_constant_MUX_n31), .ZN(
        Midori_rounds_round_Constant[0]) );
  INV_X1 Midori_rounds_constant_MUX_U31 ( .A(Midori_rounds_constant_MUX_n44), 
        .ZN(Midori_rounds_constant_MUX_n31) );
  AOI221_X1 Midori_rounds_constant_MUX_U30 ( .B1(round_Signal[3]), .B2(
        Midori_rounds_constant_MUX_n18), .C1(Midori_rounds_constant_MUX_n15), 
        .C2(enc_dec), .A(Midori_rounds_constant_MUX_n68), .ZN(
        Midori_rounds_constant_MUX_n44) );
  OR2_X1 Midori_rounds_constant_MUX_U29 ( .A1(Midori_rounds_constant_MUX_n23), 
        .A2(Midori_rounds_constant_MUX_n34), .ZN(
        Midori_rounds_constant_MUX_n68) );
  NAND2_X1 Midori_rounds_constant_MUX_U28 ( .A1(Midori_rounds_constant_MUX_n14), .A2(Midori_rounds_n1267), .ZN(Midori_rounds_constant_MUX_n34) );
  NOR2_X1 Midori_rounds_constant_MUX_U27 ( .A1(Midori_rounds_constant_MUX_n52), 
        .A2(Midori_rounds_constant_MUX_n48), .ZN(
        Midori_rounds_constant_MUX_n47) );
  OAI22_X1 Midori_rounds_constant_MUX_U26 ( .A1(Midori_rounds_constant_MUX_n24), .A2(Midori_rounds_constant_MUX_n41), .B1(Midori_rounds_constant_MUX_n42), 
        .B2(Midori_rounds_constant_MUX_n13), .ZN(
        Midori_rounds_constant_MUX_n48) );
  OAI22_X1 Midori_rounds_constant_MUX_U25 ( .A1(Midori_rounds_constant_MUX_n43), .A2(Midori_rounds_constant_MUX_n41), .B1(Midori_rounds_constant_MUX_n42), 
        .B2(Midori_rounds_constant_MUX_n40), .ZN(
        Midori_rounds_constant_MUX_n52) );
  NAND2_X1 Midori_rounds_constant_MUX_U24 ( .A1(round_Signal[1]), .A2(
        Midori_rounds_constant_MUX_n12), .ZN(Midori_rounds_constant_MUX_n40)
         );
  NOR2_X1 Midori_rounds_constant_MUX_U23 ( .A1(round_Signal[3]), .A2(enc_dec), 
        .ZN(Midori_rounds_constant_MUX_n12) );
  NAND3_X1 Midori_rounds_constant_MUX_U22 ( .A1(round_Signal[3]), .A2(enc_dec), 
        .A3(Midori_rounds_constant_MUX_n23), .ZN(
        Midori_rounds_constant_MUX_n43) );
  NOR2_X1 Midori_rounds_constant_MUX_U21 ( .A1(Midori_rounds_constant_MUX_n66), 
        .A2(Midori_rounds_constant_MUX_n20), .ZN(
        Midori_rounds_constant_MUX_n62) );
  OAI22_X1 Midori_rounds_constant_MUX_U20 ( .A1(Midori_rounds_constant_MUX_n33), .A2(Midori_rounds_constant_MUX_n42), .B1(Midori_rounds_constant_MUX_n28), 
        .B2(Midori_rounds_constant_MUX_n41), .ZN(
        Midori_rounds_constant_MUX_n20) );
  NAND3_X1 Midori_rounds_constant_MUX_U19 ( .A1(round_Signal[1]), .A2(enc_dec), 
        .A3(Midori_rounds_constant_MUX_n15), .ZN(
        Midori_rounds_constant_MUX_n28) );
  NAND3_X1 Midori_rounds_constant_MUX_U18 ( .A1(Midori_rounds_constant_MUX_n23), .A2(Midori_rounds_constant_MUX_n18), .A3(round_Signal[3]), .ZN(
        Midori_rounds_constant_MUX_n33) );
  OAI22_X1 Midori_rounds_constant_MUX_U17 ( .A1(Midori_rounds_constant_MUX_n24), .A2(Midori_rounds_constant_MUX_n42), .B1(Midori_rounds_constant_MUX_n41), 
        .B2(Midori_rounds_constant_MUX_n13), .ZN(
        Midori_rounds_constant_MUX_n66) );
  NAND2_X1 Midori_rounds_constant_MUX_U16 ( .A1(enc_dec), .A2(
        Midori_rounds_constant_MUX_n17), .ZN(Midori_rounds_constant_MUX_n13)
         );
  NAND3_X1 Midori_rounds_constant_MUX_U15 ( .A1(Midori_rounds_constant_MUX_n15), .A2(Midori_rounds_constant_MUX_n23), .A3(Midori_rounds_constant_MUX_n18), 
        .ZN(Midori_rounds_constant_MUX_n24) );
  INV_X1 Midori_rounds_constant_MUX_U14 ( .A(Midori_rounds_constant_MUX_n30), 
        .ZN(Midori_rounds_constant_MUX_n16) );
  OAI22_X1 Midori_rounds_constant_MUX_U13 ( .A1(Midori_rounds_constant_MUX_n35), .A2(Midori_rounds_constant_MUX_n41), .B1(Midori_rounds_constant_MUX_n29), 
        .B2(Midori_rounds_constant_MUX_n42), .ZN(
        Midori_rounds_constant_MUX_n30) );
  NAND2_X1 Midori_rounds_constant_MUX_U12 ( .A1(Midori_rounds_constant_MUX_n14), .A2(Midori_rounds_constant_MUX_n11), .ZN(Midori_rounds_constant_MUX_n42) );
  INV_X1 Midori_rounds_constant_MUX_U11 ( .A(round_Signal[2]), .ZN(
        Midori_rounds_constant_MUX_n14) );
  NAND2_X1 Midori_rounds_constant_MUX_U10 ( .A1(Midori_rounds_constant_MUX_n18), .A2(Midori_rounds_constant_MUX_n17), .ZN(Midori_rounds_constant_MUX_n29) );
  NOR2_X1 Midori_rounds_constant_MUX_U9 ( .A1(Midori_rounds_constant_MUX_n15), 
        .A2(Midori_rounds_constant_MUX_n23), .ZN(
        Midori_rounds_constant_MUX_n17) );
  INV_X1 Midori_rounds_constant_MUX_U8 ( .A(enc_dec), .ZN(
        Midori_rounds_constant_MUX_n18) );
  NAND2_X1 Midori_rounds_constant_MUX_U7 ( .A1(Midori_rounds_constant_MUX_n11), 
        .A2(round_Signal[2]), .ZN(Midori_rounds_constant_MUX_n41) );
  NAND3_X1 Midori_rounds_constant_MUX_U6 ( .A1(Midori_rounds_constant_MUX_n15), 
        .A2(Midori_rounds_constant_MUX_n23), .A3(enc_dec), .ZN(
        Midori_rounds_constant_MUX_n35) );
  INV_X1 Midori_rounds_constant_MUX_U5 ( .A(round_Signal[1]), .ZN(
        Midori_rounds_constant_MUX_n23) );
  INV_X1 Midori_rounds_constant_MUX_U4 ( .A(round_Signal[3]), .ZN(
        Midori_rounds_constant_MUX_n15) );
  INV_X1 Midori_rounds_constant_MUX_U3 ( .A(Midori_rounds_n1267), .ZN(
        Midori_rounds_constant_MUX_n11) );
  NAND2_X1 Midori_rounds_constant_MUX_U2 ( .A1(Midori_rounds_constant_MUX_n55), 
        .A2(Midori_rounds_constant_MUX_n10), .ZN(
        Midori_rounds_round_Constant[5]) );
  NOR2_X1 Midori_rounds_constant_MUX_U1 ( .A1(Midori_rounds_constant_MUX_n57), 
        .A2(Midori_rounds_constant_MUX_n56), .ZN(
        Midori_rounds_constant_MUX_n10) );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_0_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_0_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_0_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_0_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_0_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_0_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_0_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_0_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_0_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_0_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_0_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_0_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_0_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_0_InputAffine_U7 ( .A(Midori_rounds_n805), .ZN(
        Midori_rounds_sub_Sub_0_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_InputAffine_U6 ( .A(Midori_rounds_n917), .B(
        Midori_rounds_n919), .Z(Midori_rounds_sub_Sub_0_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_InputAffine_U5 ( .A(Midori_rounds_n917), .B(
        Midori_rounds_sub_Sub_0_F_in3[2]), .Z(Midori_rounds_sub_Sub_0_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_InputAffine_U4 ( .A(Midori_rounds_n853), .B(
        Midori_rounds_n855), .Z(Midori_rounds_sub_Sub_0_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_InputAffine_U3 ( .A(Midori_rounds_n853), .B(
        Midori_rounds_sub_Sub_0_F_in2[2]), .Z(Midori_rounds_sub_Sub_0_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_InputAffine_U2 ( .A(Midori_rounds_n789), 
        .B(Midori_rounds_n806), .ZN(Midori_rounds_sub_Sub_0_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_InputAffine_U1 ( .A(Midori_rounds_n789), .B(
        Midori_rounds_sub_Sub_0_F_in1[2]), .Z(Midori_rounds_sub_Sub_0_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U18 ( .A(Midori_rounds_sub_Sub_0_F_n4), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_0_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U17 ( .A(r[2]), .B(
        Midori_rounds_sub_Sub_0_F_q3[3]), .ZN(Midori_rounds_sub_Sub_0_F_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U16 ( .A(Midori_rounds_sub_Sub_0_F_n3), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_0_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U15 ( .A(r[0]), .B(
        Midori_rounds_sub_Sub_0_F_q3[2]), .ZN(Midori_rounds_sub_Sub_0_F_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U14 ( .A(Midori_rounds_sub_Sub_0_F_n2), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_0_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U13 ( .A(r[6]), .B(
        Midori_rounds_sub_Sub_0_F_q3[1]), .ZN(Midori_rounds_sub_Sub_0_F_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U12 ( .A(Midori_rounds_sub_Sub_0_F_n1), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_0_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_U11 ( .A(r[4]), .B(
        Midori_rounds_sub_Sub_0_F_q3[0]), .ZN(Midori_rounds_sub_Sub_0_F_n1) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U10 ( .A(r[3]), .B(
        Midori_rounds_sub_Sub_0_F_q2[3]), .Z(Midori_rounds_sub_Sub_0_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U9 ( .A(r[1]), .B(
        Midori_rounds_sub_Sub_0_F_q2[2]), .Z(Midori_rounds_sub_Sub_0_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U8 ( .A(r[7]), .B(
        Midori_rounds_sub_Sub_0_F_q2[1]), .Z(Midori_rounds_sub_Sub_0_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U7 ( .A(r[5]), .B(
        Midori_rounds_sub_Sub_0_F_q2[0]), .Z(Midori_rounds_sub_Sub_0_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U6 ( .A(r[2]), .B(
        Midori_rounds_sub_Sub_0_F_q1[3]), .Z(Midori_rounds_sub_Sub_0_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U5 ( .A(r[0]), .B(
        Midori_rounds_sub_Sub_0_F_q1[2]), .Z(Midori_rounds_sub_Sub_0_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U4 ( .A(r[6]), .B(
        Midori_rounds_sub_Sub_0_F_q1[1]), .Z(Midori_rounds_sub_Sub_0_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_F_U3 ( .A(r[4]), .B(
        Midori_rounds_sub_Sub_0_F_q1[0]), .Z(Midori_rounds_sub_Sub_0_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_0_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_0_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_0_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_0_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_0_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_0_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_0_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_0_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_0_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_0_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_0_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_0_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_0_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_0_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_0_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_0_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_0_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_0_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_0_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_0_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_0_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_0_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_0_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_0_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_0_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_0_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_0_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_0_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_0_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_0_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_0_G_U3 ( .A(Midori_rounds_sub_Sub_0_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_0_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_0_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[49]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[49]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[49]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_0_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_0_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_0_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .A2(Midori_rounds_sub_Sub_0_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_0_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[3]), .A2(Midori_rounds_sub_Sub_0_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_0_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .A2(Midori_rounds_sub_Sub_0_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_0_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .A2(Midori_rounds_sub_Sub_0_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_0_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq2[3]), .A2(Midori_rounds_sub_Sub_0_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_0_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_0_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_0_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq3[1]), .A2(Midori_rounds_sub_Sub_0_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .A2(Midori_rounds_sub_Sub_0_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_0_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .A2(Midori_rounds_sub_Sub_0_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_0_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[3]), .A2(Midori_rounds_sub_Sub_0_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_0_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .A2(Midori_rounds_sub_Sub_0_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_0_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .A2(Midori_rounds_sub_Sub_0_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_0_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_0_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .A2(Midori_rounds_sub_Sub_0_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_0_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq3[1]), .A2(Midori_rounds_sub_Sub_0_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_0_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_Rq1[3]), .B2(Midori_rounds_sub_Sub_0_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_0_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[3]), .A2(Midori_rounds_sub_Sub_0_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_0_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_Rq3[1]), .C2(Midori_rounds_sub_Sub_0_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_0_Rq1[3]), .B(
        Midori_rounds_sub_Sub_0_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq3[1]), .A2(Midori_rounds_sub_Sub_0_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_0_Rq2[2]), .A(
        Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_0_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_0_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_Rq3[1]), .C2(Midori_rounds_sub_Sub_0_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_0_Rq2[3]), .B(
        Midori_rounds_sub_Sub_0_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq3[1]), .A2(Midori_rounds_sub_Sub_0_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_0_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .C2(Midori_rounds_sub_Sub_0_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_0_Rq3[3]), .B(
        Midori_rounds_sub_Sub_0_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_0_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_Rq1[1]), .A2(Midori_rounds_sub_Sub_0_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_0_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_0_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_0_Rq3[2]), .A(
        Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_0_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_0_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[48]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[48]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[48]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[50]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[50]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[50]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[51]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[51]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[51]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_0_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_0_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_1_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_1_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_1_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_1_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_1_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_1_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_1_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_1_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_1_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_1_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_1_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_1_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_1_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_1_InputAffine_U7 ( .A(Midori_rounds_n808), .ZN(
        Midori_rounds_sub_Sub_1_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_InputAffine_U6 ( .A(Midori_rounds_n921), .B(
        Midori_rounds_n923), .Z(Midori_rounds_sub_Sub_1_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_InputAffine_U5 ( .A(Midori_rounds_n921), .B(
        Midori_rounds_sub_Sub_1_F_in3[2]), .Z(Midori_rounds_sub_Sub_1_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_InputAffine_U4 ( .A(Midori_rounds_n857), .B(
        Midori_rounds_n859), .Z(Midori_rounds_sub_Sub_1_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_InputAffine_U3 ( .A(Midori_rounds_n857), .B(
        Midori_rounds_sub_Sub_1_F_in2[2]), .Z(Midori_rounds_sub_Sub_1_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_InputAffine_U2 ( .A(Midori_rounds_n790), 
        .B(Midori_rounds_n809), .ZN(Midori_rounds_sub_Sub_1_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_InputAffine_U1 ( .A(Midori_rounds_n790), .B(
        Midori_rounds_sub_Sub_1_F_in1[2]), .Z(Midori_rounds_sub_Sub_1_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U18 ( .A(Midori_rounds_sub_Sub_1_F_n12), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_1_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U17 ( .A(r[10]), .B(
        Midori_rounds_sub_Sub_1_F_q3[3]), .ZN(Midori_rounds_sub_Sub_1_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U16 ( .A(Midori_rounds_sub_Sub_1_F_n11), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_1_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U15 ( .A(r[8]), .B(
        Midori_rounds_sub_Sub_1_F_q3[2]), .ZN(Midori_rounds_sub_Sub_1_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U14 ( .A(Midori_rounds_sub_Sub_1_F_n10), 
        .B(r[15]), .ZN(Midori_rounds_sub_Sub_1_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U13 ( .A(r[14]), .B(
        Midori_rounds_sub_Sub_1_F_q3[1]), .ZN(Midori_rounds_sub_Sub_1_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U12 ( .A(Midori_rounds_sub_Sub_1_F_n9), 
        .B(r[13]), .ZN(Midori_rounds_sub_Sub_1_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_U11 ( .A(r[12]), .B(
        Midori_rounds_sub_Sub_1_F_q3[0]), .ZN(Midori_rounds_sub_Sub_1_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U10 ( .A(r[11]), .B(
        Midori_rounds_sub_Sub_1_F_q2[3]), .Z(Midori_rounds_sub_Sub_1_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U9 ( .A(r[9]), .B(
        Midori_rounds_sub_Sub_1_F_q2[2]), .Z(Midori_rounds_sub_Sub_1_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U8 ( .A(r[15]), .B(
        Midori_rounds_sub_Sub_1_F_q2[1]), .Z(Midori_rounds_sub_Sub_1_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U7 ( .A(r[13]), .B(
        Midori_rounds_sub_Sub_1_F_q2[0]), .Z(Midori_rounds_sub_Sub_1_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U6 ( .A(r[10]), .B(
        Midori_rounds_sub_Sub_1_F_q1[3]), .Z(Midori_rounds_sub_Sub_1_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U5 ( .A(r[8]), .B(
        Midori_rounds_sub_Sub_1_F_q1[2]), .Z(Midori_rounds_sub_Sub_1_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U4 ( .A(r[14]), .B(
        Midori_rounds_sub_Sub_1_F_q1[1]), .Z(Midori_rounds_sub_Sub_1_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_F_U3 ( .A(r[12]), .B(
        Midori_rounds_sub_Sub_1_F_q1[0]), .Z(Midori_rounds_sub_Sub_1_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_1_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_1_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_1_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_1_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_1_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_1_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_1_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_1_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_1_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_1_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_1_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_1_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_1_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_1_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_1_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_1_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_1_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_1_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_1_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_1_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_1_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_1_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_1_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_1_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_1_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_1_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_1_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_1_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_1_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_1_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_1_G_U3 ( .A(Midori_rounds_sub_Sub_1_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_1_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_1_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[45]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[45]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[45]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_1_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_1_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_1_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .A2(Midori_rounds_sub_Sub_1_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_1_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[3]), .A2(Midori_rounds_sub_Sub_1_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_1_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .A2(Midori_rounds_sub_Sub_1_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_1_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .A2(Midori_rounds_sub_Sub_1_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_1_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq2[3]), .A2(Midori_rounds_sub_Sub_1_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_1_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_1_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_1_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq3[1]), .A2(Midori_rounds_sub_Sub_1_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .A2(Midori_rounds_sub_Sub_1_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_1_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .A2(Midori_rounds_sub_Sub_1_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_1_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[3]), .A2(Midori_rounds_sub_Sub_1_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_1_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .A2(Midori_rounds_sub_Sub_1_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_1_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .A2(Midori_rounds_sub_Sub_1_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_1_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_1_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .A2(Midori_rounds_sub_Sub_1_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_1_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq3[1]), .A2(Midori_rounds_sub_Sub_1_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_1_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_Rq1[3]), .B2(Midori_rounds_sub_Sub_1_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_1_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[3]), .A2(Midori_rounds_sub_Sub_1_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_1_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_Rq3[1]), .C2(Midori_rounds_sub_Sub_1_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_1_Rq1[3]), .B(
        Midori_rounds_sub_Sub_1_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq3[1]), .A2(Midori_rounds_sub_Sub_1_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_1_Rq2[2]), .A(
        Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_1_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_1_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_Rq3[1]), .C2(Midori_rounds_sub_Sub_1_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_1_Rq2[3]), .B(
        Midori_rounds_sub_Sub_1_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq3[1]), .A2(Midori_rounds_sub_Sub_1_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_1_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .C2(Midori_rounds_sub_Sub_1_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_1_Rq3[3]), .B(
        Midori_rounds_sub_Sub_1_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_1_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_Rq1[1]), .A2(Midori_rounds_sub_Sub_1_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_1_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_1_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_1_Rq3[2]), .A(
        Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_1_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_1_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[44]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[44]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[44]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[46]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[46]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[46]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[47]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[47]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[47]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_1_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_1_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_2_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_2_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_2_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_2_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_2_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_2_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_2_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_2_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_2_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_2_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_2_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_2_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_2_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_2_InputAffine_U7 ( .A(Midori_rounds_n811), .ZN(
        Midori_rounds_sub_Sub_2_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_InputAffine_U6 ( .A(Midori_rounds_n925), .B(
        Midori_rounds_n927), .Z(Midori_rounds_sub_Sub_2_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_InputAffine_U5 ( .A(Midori_rounds_n925), .B(
        Midori_rounds_sub_Sub_2_F_in3[2]), .Z(Midori_rounds_sub_Sub_2_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_InputAffine_U4 ( .A(Midori_rounds_n861), .B(
        Midori_rounds_n863), .Z(Midori_rounds_sub_Sub_2_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_InputAffine_U3 ( .A(Midori_rounds_n861), .B(
        Midori_rounds_sub_Sub_2_F_in2[2]), .Z(Midori_rounds_sub_Sub_2_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_InputAffine_U2 ( .A(Midori_rounds_n791), 
        .B(Midori_rounds_n812), .ZN(Midori_rounds_sub_Sub_2_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_InputAffine_U1 ( .A(Midori_rounds_n791), .B(
        Midori_rounds_sub_Sub_2_F_in1[2]), .Z(Midori_rounds_sub_Sub_2_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U18 ( .A(Midori_rounds_sub_Sub_2_F_n12), 
        .B(r[19]), .ZN(Midori_rounds_sub_Sub_2_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U17 ( .A(r[18]), .B(
        Midori_rounds_sub_Sub_2_F_q3[3]), .ZN(Midori_rounds_sub_Sub_2_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U16 ( .A(Midori_rounds_sub_Sub_2_F_n11), 
        .B(r[17]), .ZN(Midori_rounds_sub_Sub_2_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U15 ( .A(r[16]), .B(
        Midori_rounds_sub_Sub_2_F_q3[2]), .ZN(Midori_rounds_sub_Sub_2_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U14 ( .A(Midori_rounds_sub_Sub_2_F_n10), 
        .B(r[23]), .ZN(Midori_rounds_sub_Sub_2_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U13 ( .A(r[22]), .B(
        Midori_rounds_sub_Sub_2_F_q3[1]), .ZN(Midori_rounds_sub_Sub_2_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U12 ( .A(Midori_rounds_sub_Sub_2_F_n9), 
        .B(r[21]), .ZN(Midori_rounds_sub_Sub_2_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_U11 ( .A(r[20]), .B(
        Midori_rounds_sub_Sub_2_F_q3[0]), .ZN(Midori_rounds_sub_Sub_2_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U10 ( .A(r[19]), .B(
        Midori_rounds_sub_Sub_2_F_q2[3]), .Z(Midori_rounds_sub_Sub_2_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U9 ( .A(r[17]), .B(
        Midori_rounds_sub_Sub_2_F_q2[2]), .Z(Midori_rounds_sub_Sub_2_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U8 ( .A(r[23]), .B(
        Midori_rounds_sub_Sub_2_F_q2[1]), .Z(Midori_rounds_sub_Sub_2_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U7 ( .A(r[21]), .B(
        Midori_rounds_sub_Sub_2_F_q2[0]), .Z(Midori_rounds_sub_Sub_2_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U6 ( .A(r[18]), .B(
        Midori_rounds_sub_Sub_2_F_q1[3]), .Z(Midori_rounds_sub_Sub_2_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U5 ( .A(r[16]), .B(
        Midori_rounds_sub_Sub_2_F_q1[2]), .Z(Midori_rounds_sub_Sub_2_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U4 ( .A(r[22]), .B(
        Midori_rounds_sub_Sub_2_F_q1[1]), .Z(Midori_rounds_sub_Sub_2_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_F_U3 ( .A(r[20]), .B(
        Midori_rounds_sub_Sub_2_F_q1[0]), .Z(Midori_rounds_sub_Sub_2_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_2_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_2_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_2_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_2_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_2_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_2_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_2_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_2_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_2_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_2_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_2_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_2_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_2_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_2_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_2_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_2_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_2_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_2_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_2_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_2_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_2_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_2_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_2_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_2_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_2_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_2_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_2_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_2_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_2_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_2_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_2_G_U3 ( .A(Midori_rounds_sub_Sub_2_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_2_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_2_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_2_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_2_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_2_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .A2(Midori_rounds_sub_Sub_2_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_2_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[3]), .A2(Midori_rounds_sub_Sub_2_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_2_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .A2(Midori_rounds_sub_Sub_2_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_2_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .A2(Midori_rounds_sub_Sub_2_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_2_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq2[3]), .A2(Midori_rounds_sub_Sub_2_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_2_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_2_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_2_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq3[1]), .A2(Midori_rounds_sub_Sub_2_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .A2(Midori_rounds_sub_Sub_2_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_2_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .A2(Midori_rounds_sub_Sub_2_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_2_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[3]), .A2(Midori_rounds_sub_Sub_2_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_2_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .A2(Midori_rounds_sub_Sub_2_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_2_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .A2(Midori_rounds_sub_Sub_2_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_2_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_2_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .A2(Midori_rounds_sub_Sub_2_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_2_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq3[1]), .A2(Midori_rounds_sub_Sub_2_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_2_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_Rq1[3]), .B2(Midori_rounds_sub_Sub_2_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_2_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[3]), .A2(Midori_rounds_sub_Sub_2_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_2_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_Rq3[1]), .C2(Midori_rounds_sub_Sub_2_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_2_Rq1[3]), .B(
        Midori_rounds_sub_Sub_2_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq3[1]), .A2(Midori_rounds_sub_Sub_2_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_2_Rq2[2]), .A(
        Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_2_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_2_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_Rq3[1]), .C2(Midori_rounds_sub_Sub_2_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_2_Rq2[3]), .B(
        Midori_rounds_sub_Sub_2_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq3[1]), .A2(Midori_rounds_sub_Sub_2_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_2_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .C2(Midori_rounds_sub_Sub_2_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_2_Rq3[3]), .B(
        Midori_rounds_sub_Sub_2_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_2_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_Rq1[1]), .A2(Midori_rounds_sub_Sub_2_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_2_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_2_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_2_Rq3[2]), .A(
        Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_2_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_2_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[8])
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[8])
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[8])
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_2_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_2_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_3_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_3_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_3_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_3_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_3_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_3_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_3_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_3_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_3_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_3_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_3_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_3_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_3_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_3_InputAffine_U7 ( .A(Midori_rounds_n814), .ZN(
        Midori_rounds_sub_Sub_3_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_InputAffine_U6 ( .A(Midori_rounds_n929), .B(
        Midori_rounds_n931), .Z(Midori_rounds_sub_Sub_3_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_InputAffine_U5 ( .A(Midori_rounds_n929), .B(
        Midori_rounds_sub_Sub_3_F_in3[2]), .Z(Midori_rounds_sub_Sub_3_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_InputAffine_U4 ( .A(Midori_rounds_n865), .B(
        Midori_rounds_n867), .Z(Midori_rounds_sub_Sub_3_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_InputAffine_U3 ( .A(Midori_rounds_n865), .B(
        Midori_rounds_sub_Sub_3_F_in2[2]), .Z(Midori_rounds_sub_Sub_3_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_InputAffine_U2 ( .A(Midori_rounds_n792), 
        .B(Midori_rounds_n815), .ZN(Midori_rounds_sub_Sub_3_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_InputAffine_U1 ( .A(Midori_rounds_n792), .B(
        Midori_rounds_sub_Sub_3_F_in1[2]), .Z(Midori_rounds_sub_Sub_3_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U18 ( .A(Midori_rounds_sub_Sub_3_F_n12), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_3_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U17 ( .A(r[26]), .B(
        Midori_rounds_sub_Sub_3_F_q3[3]), .ZN(Midori_rounds_sub_Sub_3_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U16 ( .A(Midori_rounds_sub_Sub_3_F_n11), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_3_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U15 ( .A(r[24]), .B(
        Midori_rounds_sub_Sub_3_F_q3[2]), .ZN(Midori_rounds_sub_Sub_3_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U14 ( .A(Midori_rounds_sub_Sub_3_F_n10), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_3_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U13 ( .A(r[30]), .B(
        Midori_rounds_sub_Sub_3_F_q3[1]), .ZN(Midori_rounds_sub_Sub_3_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U12 ( .A(Midori_rounds_sub_Sub_3_F_n9), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_3_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_U11 ( .A(r[28]), .B(
        Midori_rounds_sub_Sub_3_F_q3[0]), .ZN(Midori_rounds_sub_Sub_3_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U10 ( .A(r[27]), .B(
        Midori_rounds_sub_Sub_3_F_q2[3]), .Z(Midori_rounds_sub_Sub_3_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U9 ( .A(r[25]), .B(
        Midori_rounds_sub_Sub_3_F_q2[2]), .Z(Midori_rounds_sub_Sub_3_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U8 ( .A(r[31]), .B(
        Midori_rounds_sub_Sub_3_F_q2[1]), .Z(Midori_rounds_sub_Sub_3_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U7 ( .A(r[29]), .B(
        Midori_rounds_sub_Sub_3_F_q2[0]), .Z(Midori_rounds_sub_Sub_3_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U6 ( .A(r[26]), .B(
        Midori_rounds_sub_Sub_3_F_q1[3]), .Z(Midori_rounds_sub_Sub_3_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U5 ( .A(r[24]), .B(
        Midori_rounds_sub_Sub_3_F_q1[2]), .Z(Midori_rounds_sub_Sub_3_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U4 ( .A(r[30]), .B(
        Midori_rounds_sub_Sub_3_F_q1[1]), .Z(Midori_rounds_sub_Sub_3_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_F_U3 ( .A(r[28]), .B(
        Midori_rounds_sub_Sub_3_F_q1[0]), .Z(Midori_rounds_sub_Sub_3_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_3_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_3_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_3_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_3_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_3_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_3_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_3_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_3_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_3_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_3_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_3_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_3_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_3_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_3_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_3_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_3_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_3_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_3_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_3_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_3_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_3_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_3_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_3_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_3_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_3_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_3_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_3_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_3_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_3_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_3_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_3_G_U3 ( .A(Midori_rounds_sub_Sub_3_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_3_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_3_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_3_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_3_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_3_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .A2(Midori_rounds_sub_Sub_3_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_3_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[3]), .A2(Midori_rounds_sub_Sub_3_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_3_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .A2(Midori_rounds_sub_Sub_3_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_3_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .A2(Midori_rounds_sub_Sub_3_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_3_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq2[3]), .A2(Midori_rounds_sub_Sub_3_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_3_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_3_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_3_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq3[1]), .A2(Midori_rounds_sub_Sub_3_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .A2(Midori_rounds_sub_Sub_3_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_3_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .A2(Midori_rounds_sub_Sub_3_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_3_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[3]), .A2(Midori_rounds_sub_Sub_3_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_3_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .A2(Midori_rounds_sub_Sub_3_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_3_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .A2(Midori_rounds_sub_Sub_3_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_3_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_3_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .A2(Midori_rounds_sub_Sub_3_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_3_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq3[1]), .A2(Midori_rounds_sub_Sub_3_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_3_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_Rq1[3]), .B2(Midori_rounds_sub_Sub_3_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_3_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[3]), .A2(Midori_rounds_sub_Sub_3_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_3_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_Rq3[1]), .C2(Midori_rounds_sub_Sub_3_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_3_Rq1[3]), .B(
        Midori_rounds_sub_Sub_3_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq3[1]), .A2(Midori_rounds_sub_Sub_3_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_3_Rq2[2]), .A(
        Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_3_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_3_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_Rq3[1]), .C2(Midori_rounds_sub_Sub_3_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_3_Rq2[3]), .B(
        Midori_rounds_sub_Sub_3_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq3[1]), .A2(Midori_rounds_sub_Sub_3_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_3_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .C2(Midori_rounds_sub_Sub_3_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_3_Rq3[3]), .B(
        Midori_rounds_sub_Sub_3_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_3_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_Rq1[1]), .A2(Midori_rounds_sub_Sub_3_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_3_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_3_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_3_Rq3[2]), .A(
        Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_3_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_3_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[20]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[20]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[20]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[23]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[23]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[23]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_3_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_3_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_4_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_4_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_4_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_4_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_4_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_4_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_4_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_4_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_4_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_4_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_4_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_4_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_4_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_4_InputAffine_U7 ( .A(Midori_rounds_n817), .ZN(
        Midori_rounds_sub_Sub_4_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_InputAffine_U6 ( .A(Midori_rounds_n933), .B(
        Midori_rounds_n935), .Z(Midori_rounds_sub_Sub_4_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_InputAffine_U5 ( .A(Midori_rounds_n933), .B(
        Midori_rounds_sub_Sub_4_F_in3[2]), .Z(Midori_rounds_sub_Sub_4_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_InputAffine_U4 ( .A(Midori_rounds_n869), .B(
        Midori_rounds_n871), .Z(Midori_rounds_sub_Sub_4_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_InputAffine_U3 ( .A(Midori_rounds_n869), .B(
        Midori_rounds_sub_Sub_4_F_in2[2]), .Z(Midori_rounds_sub_Sub_4_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_InputAffine_U2 ( .A(Midori_rounds_n793), 
        .B(Midori_rounds_n818), .ZN(Midori_rounds_sub_Sub_4_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_InputAffine_U1 ( .A(Midori_rounds_n793), .B(
        Midori_rounds_sub_Sub_4_F_in1[2]), .Z(Midori_rounds_sub_Sub_4_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U18 ( .A(Midori_rounds_sub_Sub_4_F_n12), 
        .B(r[35]), .ZN(Midori_rounds_sub_Sub_4_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U17 ( .A(r[34]), .B(
        Midori_rounds_sub_Sub_4_F_q3[3]), .ZN(Midori_rounds_sub_Sub_4_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U16 ( .A(Midori_rounds_sub_Sub_4_F_n11), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_4_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U15 ( .A(r[32]), .B(
        Midori_rounds_sub_Sub_4_F_q3[2]), .ZN(Midori_rounds_sub_Sub_4_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U14 ( .A(Midori_rounds_sub_Sub_4_F_n10), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_4_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U13 ( .A(r[38]), .B(
        Midori_rounds_sub_Sub_4_F_q3[1]), .ZN(Midori_rounds_sub_Sub_4_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U12 ( .A(Midori_rounds_sub_Sub_4_F_n9), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_4_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_U11 ( .A(r[36]), .B(
        Midori_rounds_sub_Sub_4_F_q3[0]), .ZN(Midori_rounds_sub_Sub_4_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U10 ( .A(r[35]), .B(
        Midori_rounds_sub_Sub_4_F_q2[3]), .Z(Midori_rounds_sub_Sub_4_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U9 ( .A(r[33]), .B(
        Midori_rounds_sub_Sub_4_F_q2[2]), .Z(Midori_rounds_sub_Sub_4_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U8 ( .A(r[39]), .B(
        Midori_rounds_sub_Sub_4_F_q2[1]), .Z(Midori_rounds_sub_Sub_4_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U7 ( .A(r[37]), .B(
        Midori_rounds_sub_Sub_4_F_q2[0]), .Z(Midori_rounds_sub_Sub_4_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U6 ( .A(r[34]), .B(
        Midori_rounds_sub_Sub_4_F_q1[3]), .Z(Midori_rounds_sub_Sub_4_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U5 ( .A(r[32]), .B(
        Midori_rounds_sub_Sub_4_F_q1[2]), .Z(Midori_rounds_sub_Sub_4_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U4 ( .A(r[38]), .B(
        Midori_rounds_sub_Sub_4_F_q1[1]), .Z(Midori_rounds_sub_Sub_4_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_F_U3 ( .A(r[36]), .B(
        Midori_rounds_sub_Sub_4_F_q1[0]), .Z(Midori_rounds_sub_Sub_4_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_4_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_4_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_4_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_4_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_4_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_4_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_4_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_4_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_4_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_4_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_4_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_4_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_4_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_4_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_4_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_4_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_4_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_4_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_4_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_4_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_4_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_4_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_4_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_4_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_4_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_4_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_4_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_4_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_4_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_4_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_4_G_U3 ( .A(Midori_rounds_sub_Sub_4_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_4_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_4_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[37]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[37]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[37]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_4_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_4_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_4_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .A2(Midori_rounds_sub_Sub_4_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_4_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[3]), .A2(Midori_rounds_sub_Sub_4_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_4_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .A2(Midori_rounds_sub_Sub_4_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_4_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .A2(Midori_rounds_sub_Sub_4_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_4_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq2[3]), .A2(Midori_rounds_sub_Sub_4_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_4_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_4_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_4_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq3[1]), .A2(Midori_rounds_sub_Sub_4_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .A2(Midori_rounds_sub_Sub_4_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_4_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .A2(Midori_rounds_sub_Sub_4_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_4_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[3]), .A2(Midori_rounds_sub_Sub_4_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_4_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .A2(Midori_rounds_sub_Sub_4_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_4_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .A2(Midori_rounds_sub_Sub_4_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_4_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_4_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .A2(Midori_rounds_sub_Sub_4_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_4_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq3[1]), .A2(Midori_rounds_sub_Sub_4_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_4_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_Rq1[3]), .B2(Midori_rounds_sub_Sub_4_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_4_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[3]), .A2(Midori_rounds_sub_Sub_4_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_4_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_Rq3[1]), .C2(Midori_rounds_sub_Sub_4_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_4_Rq1[3]), .B(
        Midori_rounds_sub_Sub_4_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq3[1]), .A2(Midori_rounds_sub_Sub_4_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_4_Rq2[2]), .A(
        Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_4_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_4_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_Rq3[1]), .C2(Midori_rounds_sub_Sub_4_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_4_Rq2[3]), .B(
        Midori_rounds_sub_Sub_4_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq3[1]), .A2(Midori_rounds_sub_Sub_4_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_4_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .C2(Midori_rounds_sub_Sub_4_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_4_Rq3[3]), .B(
        Midori_rounds_sub_Sub_4_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_4_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_Rq1[1]), .A2(Midori_rounds_sub_Sub_4_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_4_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_4_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_4_Rq3[2]), .A(
        Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_4_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_4_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[36]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[36]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[36]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[38]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[38]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[38]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[39]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[39]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[39]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_4_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_4_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_5_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_5_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_5_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_5_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_5_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_5_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_5_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_5_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_5_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_5_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_5_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_5_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_5_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_5_InputAffine_U7 ( .A(Midori_rounds_n820), .ZN(
        Midori_rounds_sub_Sub_5_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_InputAffine_U6 ( .A(Midori_rounds_n937), .B(
        Midori_rounds_n939), .Z(Midori_rounds_sub_Sub_5_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_InputAffine_U5 ( .A(Midori_rounds_n937), .B(
        Midori_rounds_sub_Sub_5_F_in3[2]), .Z(Midori_rounds_sub_Sub_5_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_InputAffine_U4 ( .A(Midori_rounds_n873), .B(
        Midori_rounds_n875), .Z(Midori_rounds_sub_Sub_5_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_InputAffine_U3 ( .A(Midori_rounds_n873), .B(
        Midori_rounds_sub_Sub_5_F_in2[2]), .Z(Midori_rounds_sub_Sub_5_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_InputAffine_U2 ( .A(Midori_rounds_n794), 
        .B(Midori_rounds_n821), .ZN(Midori_rounds_sub_Sub_5_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_InputAffine_U1 ( .A(Midori_rounds_n794), .B(
        Midori_rounds_sub_Sub_5_F_in1[2]), .Z(Midori_rounds_sub_Sub_5_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U18 ( .A(Midori_rounds_sub_Sub_5_F_n12), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_5_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U17 ( .A(r[42]), .B(
        Midori_rounds_sub_Sub_5_F_q3[3]), .ZN(Midori_rounds_sub_Sub_5_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U16 ( .A(Midori_rounds_sub_Sub_5_F_n11), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_5_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U15 ( .A(r[40]), .B(
        Midori_rounds_sub_Sub_5_F_q3[2]), .ZN(Midori_rounds_sub_Sub_5_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U14 ( .A(Midori_rounds_sub_Sub_5_F_n10), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_5_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U13 ( .A(r[46]), .B(
        Midori_rounds_sub_Sub_5_F_q3[1]), .ZN(Midori_rounds_sub_Sub_5_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U12 ( .A(Midori_rounds_sub_Sub_5_F_n9), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_5_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_U11 ( .A(r[44]), .B(
        Midori_rounds_sub_Sub_5_F_q3[0]), .ZN(Midori_rounds_sub_Sub_5_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U10 ( .A(r[43]), .B(
        Midori_rounds_sub_Sub_5_F_q2[3]), .Z(Midori_rounds_sub_Sub_5_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U9 ( .A(r[41]), .B(
        Midori_rounds_sub_Sub_5_F_q2[2]), .Z(Midori_rounds_sub_Sub_5_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U8 ( .A(r[47]), .B(
        Midori_rounds_sub_Sub_5_F_q2[1]), .Z(Midori_rounds_sub_Sub_5_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U7 ( .A(r[45]), .B(
        Midori_rounds_sub_Sub_5_F_q2[0]), .Z(Midori_rounds_sub_Sub_5_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U6 ( .A(r[42]), .B(
        Midori_rounds_sub_Sub_5_F_q1[3]), .Z(Midori_rounds_sub_Sub_5_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U5 ( .A(r[40]), .B(
        Midori_rounds_sub_Sub_5_F_q1[2]), .Z(Midori_rounds_sub_Sub_5_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U4 ( .A(r[46]), .B(
        Midori_rounds_sub_Sub_5_F_q1[1]), .Z(Midori_rounds_sub_Sub_5_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_F_U3 ( .A(r[44]), .B(
        Midori_rounds_sub_Sub_5_F_q1[0]), .Z(Midori_rounds_sub_Sub_5_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_5_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_5_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_5_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_5_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_5_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_5_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_5_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_5_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_5_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_5_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_5_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_5_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_5_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_5_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_5_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_5_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_5_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_5_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_5_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_5_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_5_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_5_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_5_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_5_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_5_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_5_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_5_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_5_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_5_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_5_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_5_G_U3 ( .A(Midori_rounds_sub_Sub_5_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_5_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_5_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[57]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[57]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[57]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_5_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_5_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_5_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .A2(Midori_rounds_sub_Sub_5_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_5_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[3]), .A2(Midori_rounds_sub_Sub_5_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_5_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .A2(Midori_rounds_sub_Sub_5_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_5_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .A2(Midori_rounds_sub_Sub_5_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_5_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq2[3]), .A2(Midori_rounds_sub_Sub_5_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_5_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_5_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_5_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq3[1]), .A2(Midori_rounds_sub_Sub_5_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .A2(Midori_rounds_sub_Sub_5_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_5_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .A2(Midori_rounds_sub_Sub_5_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_5_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[3]), .A2(Midori_rounds_sub_Sub_5_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_5_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .A2(Midori_rounds_sub_Sub_5_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_5_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .A2(Midori_rounds_sub_Sub_5_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_5_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_5_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .A2(Midori_rounds_sub_Sub_5_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_5_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq3[1]), .A2(Midori_rounds_sub_Sub_5_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_5_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_Rq1[3]), .B2(Midori_rounds_sub_Sub_5_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_5_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[3]), .A2(Midori_rounds_sub_Sub_5_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_5_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_Rq3[1]), .C2(Midori_rounds_sub_Sub_5_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_5_Rq1[3]), .B(
        Midori_rounds_sub_Sub_5_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq3[1]), .A2(Midori_rounds_sub_Sub_5_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_5_Rq2[2]), .A(
        Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_5_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_5_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_Rq3[1]), .C2(Midori_rounds_sub_Sub_5_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_5_Rq2[3]), .B(
        Midori_rounds_sub_Sub_5_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq3[1]), .A2(Midori_rounds_sub_Sub_5_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_5_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .C2(Midori_rounds_sub_Sub_5_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_5_Rq3[3]), .B(
        Midori_rounds_sub_Sub_5_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_5_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_Rq1[1]), .A2(Midori_rounds_sub_Sub_5_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_5_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_5_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_5_Rq3[2]), .A(
        Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_5_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_5_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[56]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[56]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[56]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[58]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[58]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[58]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[59]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[59]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[59]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_5_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_5_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_6_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_6_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_6_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_6_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_6_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_6_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_6_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_6_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_6_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_6_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_6_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_6_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_6_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_6_InputAffine_U7 ( .A(Midori_rounds_n823), .ZN(
        Midori_rounds_sub_Sub_6_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_InputAffine_U6 ( .A(Midori_rounds_n941), .B(
        Midori_rounds_n943), .Z(Midori_rounds_sub_Sub_6_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_InputAffine_U5 ( .A(Midori_rounds_n941), .B(
        Midori_rounds_sub_Sub_6_F_in3[2]), .Z(Midori_rounds_sub_Sub_6_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_InputAffine_U4 ( .A(Midori_rounds_n877), .B(
        Midori_rounds_n879), .Z(Midori_rounds_sub_Sub_6_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_InputAffine_U3 ( .A(Midori_rounds_n877), .B(
        Midori_rounds_sub_Sub_6_F_in2[2]), .Z(Midori_rounds_sub_Sub_6_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_InputAffine_U2 ( .A(Midori_rounds_n795), 
        .B(Midori_rounds_n824), .ZN(Midori_rounds_sub_Sub_6_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_InputAffine_U1 ( .A(Midori_rounds_n795), .B(
        Midori_rounds_sub_Sub_6_F_in1[2]), .Z(Midori_rounds_sub_Sub_6_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U18 ( .A(Midori_rounds_sub_Sub_6_F_n12), 
        .B(r[51]), .ZN(Midori_rounds_sub_Sub_6_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U17 ( .A(r[50]), .B(
        Midori_rounds_sub_Sub_6_F_q3[3]), .ZN(Midori_rounds_sub_Sub_6_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U16 ( .A(Midori_rounds_sub_Sub_6_F_n11), 
        .B(r[49]), .ZN(Midori_rounds_sub_Sub_6_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U15 ( .A(r[48]), .B(
        Midori_rounds_sub_Sub_6_F_q3[2]), .ZN(Midori_rounds_sub_Sub_6_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U14 ( .A(Midori_rounds_sub_Sub_6_F_n10), 
        .B(r[55]), .ZN(Midori_rounds_sub_Sub_6_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U13 ( .A(r[54]), .B(
        Midori_rounds_sub_Sub_6_F_q3[1]), .ZN(Midori_rounds_sub_Sub_6_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U12 ( .A(Midori_rounds_sub_Sub_6_F_n9), 
        .B(r[53]), .ZN(Midori_rounds_sub_Sub_6_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_U11 ( .A(r[52]), .B(
        Midori_rounds_sub_Sub_6_F_q3[0]), .ZN(Midori_rounds_sub_Sub_6_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U10 ( .A(r[51]), .B(
        Midori_rounds_sub_Sub_6_F_q2[3]), .Z(Midori_rounds_sub_Sub_6_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U9 ( .A(r[49]), .B(
        Midori_rounds_sub_Sub_6_F_q2[2]), .Z(Midori_rounds_sub_Sub_6_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U8 ( .A(r[55]), .B(
        Midori_rounds_sub_Sub_6_F_q2[1]), .Z(Midori_rounds_sub_Sub_6_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U7 ( .A(r[53]), .B(
        Midori_rounds_sub_Sub_6_F_q2[0]), .Z(Midori_rounds_sub_Sub_6_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U6 ( .A(r[50]), .B(
        Midori_rounds_sub_Sub_6_F_q1[3]), .Z(Midori_rounds_sub_Sub_6_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U5 ( .A(r[48]), .B(
        Midori_rounds_sub_Sub_6_F_q1[2]), .Z(Midori_rounds_sub_Sub_6_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U4 ( .A(r[54]), .B(
        Midori_rounds_sub_Sub_6_F_q1[1]), .Z(Midori_rounds_sub_Sub_6_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_F_U3 ( .A(r[52]), .B(
        Midori_rounds_sub_Sub_6_F_q1[0]), .Z(Midori_rounds_sub_Sub_6_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_6_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_6_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_6_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_6_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_6_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_6_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_6_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_6_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_6_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_6_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_6_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_6_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_6_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_6_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_6_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_6_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_6_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_6_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_6_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_6_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_6_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_6_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_6_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_6_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_6_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_6_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_6_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_6_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_6_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_6_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_6_G_U3 ( .A(Midori_rounds_sub_Sub_6_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_6_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_6_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_6_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_6_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_6_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .A2(Midori_rounds_sub_Sub_6_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_6_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[3]), .A2(Midori_rounds_sub_Sub_6_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_6_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .A2(Midori_rounds_sub_Sub_6_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_6_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .A2(Midori_rounds_sub_Sub_6_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_6_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq2[3]), .A2(Midori_rounds_sub_Sub_6_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_6_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_6_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_6_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq3[1]), .A2(Midori_rounds_sub_Sub_6_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .A2(Midori_rounds_sub_Sub_6_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_6_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .A2(Midori_rounds_sub_Sub_6_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_6_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[3]), .A2(Midori_rounds_sub_Sub_6_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_6_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .A2(Midori_rounds_sub_Sub_6_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_6_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .A2(Midori_rounds_sub_Sub_6_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_6_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_6_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .A2(Midori_rounds_sub_Sub_6_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_6_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq3[1]), .A2(Midori_rounds_sub_Sub_6_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_6_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_Rq1[3]), .B2(Midori_rounds_sub_Sub_6_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_6_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[3]), .A2(Midori_rounds_sub_Sub_6_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_6_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_Rq3[1]), .C2(Midori_rounds_sub_Sub_6_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_6_Rq1[3]), .B(
        Midori_rounds_sub_Sub_6_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq3[1]), .A2(Midori_rounds_sub_Sub_6_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_6_Rq2[2]), .A(
        Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_6_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_6_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_Rq3[1]), .C2(Midori_rounds_sub_Sub_6_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_6_Rq2[3]), .B(
        Midori_rounds_sub_Sub_6_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq3[1]), .A2(Midori_rounds_sub_Sub_6_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_6_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .C2(Midori_rounds_sub_Sub_6_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_6_Rq3[3]), .B(
        Midori_rounds_sub_Sub_6_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_6_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_Rq1[1]), .A2(Midori_rounds_sub_Sub_6_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_6_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_6_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_6_Rq3[2]), .A(
        Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_6_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_6_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[28]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[28]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[28]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[30]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[30]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[30]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[31]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[31]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[31]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_6_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_6_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_7_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_7_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_7_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_7_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_7_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_7_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_7_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_7_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_7_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_7_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_7_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_7_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_7_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_7_InputAffine_U7 ( .A(Midori_rounds_n826), .ZN(
        Midori_rounds_sub_Sub_7_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_InputAffine_U6 ( .A(Midori_rounds_n945), .B(
        Midori_rounds_n947), .Z(Midori_rounds_sub_Sub_7_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_InputAffine_U5 ( .A(Midori_rounds_n945), .B(
        Midori_rounds_sub_Sub_7_F_in3[2]), .Z(Midori_rounds_sub_Sub_7_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_InputAffine_U4 ( .A(Midori_rounds_n881), .B(
        Midori_rounds_n883), .Z(Midori_rounds_sub_Sub_7_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_InputAffine_U3 ( .A(Midori_rounds_n881), .B(
        Midori_rounds_sub_Sub_7_F_in2[2]), .Z(Midori_rounds_sub_Sub_7_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_InputAffine_U2 ( .A(Midori_rounds_n796), 
        .B(Midori_rounds_n827), .ZN(Midori_rounds_sub_Sub_7_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_InputAffine_U1 ( .A(Midori_rounds_n796), .B(
        Midori_rounds_sub_Sub_7_F_in1[2]), .Z(Midori_rounds_sub_Sub_7_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U18 ( .A(Midori_rounds_sub_Sub_7_F_n12), 
        .B(r[59]), .ZN(Midori_rounds_sub_Sub_7_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U17 ( .A(r[58]), .B(
        Midori_rounds_sub_Sub_7_F_q3[3]), .ZN(Midori_rounds_sub_Sub_7_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U16 ( .A(Midori_rounds_sub_Sub_7_F_n11), 
        .B(r[57]), .ZN(Midori_rounds_sub_Sub_7_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U15 ( .A(r[56]), .B(
        Midori_rounds_sub_Sub_7_F_q3[2]), .ZN(Midori_rounds_sub_Sub_7_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U14 ( .A(Midori_rounds_sub_Sub_7_F_n10), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_7_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U13 ( .A(r[62]), .B(
        Midori_rounds_sub_Sub_7_F_q3[1]), .ZN(Midori_rounds_sub_Sub_7_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U12 ( .A(Midori_rounds_sub_Sub_7_F_n9), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_7_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_U11 ( .A(r[60]), .B(
        Midori_rounds_sub_Sub_7_F_q3[0]), .ZN(Midori_rounds_sub_Sub_7_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U10 ( .A(r[59]), .B(
        Midori_rounds_sub_Sub_7_F_q2[3]), .Z(Midori_rounds_sub_Sub_7_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U9 ( .A(r[57]), .B(
        Midori_rounds_sub_Sub_7_F_q2[2]), .Z(Midori_rounds_sub_Sub_7_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U8 ( .A(r[63]), .B(
        Midori_rounds_sub_Sub_7_F_q2[1]), .Z(Midori_rounds_sub_Sub_7_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U7 ( .A(r[61]), .B(
        Midori_rounds_sub_Sub_7_F_q2[0]), .Z(Midori_rounds_sub_Sub_7_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U6 ( .A(r[58]), .B(
        Midori_rounds_sub_Sub_7_F_q1[3]), .Z(Midori_rounds_sub_Sub_7_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U5 ( .A(r[56]), .B(
        Midori_rounds_sub_Sub_7_F_q1[2]), .Z(Midori_rounds_sub_Sub_7_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U4 ( .A(r[62]), .B(
        Midori_rounds_sub_Sub_7_F_q1[1]), .Z(Midori_rounds_sub_Sub_7_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_F_U3 ( .A(r[60]), .B(
        Midori_rounds_sub_Sub_7_F_q1[0]), .Z(Midori_rounds_sub_Sub_7_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_7_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_7_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_7_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_7_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_7_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_7_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_7_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_7_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_7_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_7_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_7_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_7_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_7_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_7_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_7_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_7_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_7_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_7_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_7_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_7_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_7_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_7_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_7_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_7_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_7_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_7_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_7_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_7_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_7_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_7_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_7_G_U3 ( .A(Midori_rounds_sub_Sub_7_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_7_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_7_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_7_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_7_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_7_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .A2(Midori_rounds_sub_Sub_7_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_7_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[3]), .A2(Midori_rounds_sub_Sub_7_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_7_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .A2(Midori_rounds_sub_Sub_7_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_7_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .A2(Midori_rounds_sub_Sub_7_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_7_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq2[3]), .A2(Midori_rounds_sub_Sub_7_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_7_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_7_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_7_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq3[1]), .A2(Midori_rounds_sub_Sub_7_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .A2(Midori_rounds_sub_Sub_7_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_7_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .A2(Midori_rounds_sub_Sub_7_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_7_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[3]), .A2(Midori_rounds_sub_Sub_7_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_7_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .A2(Midori_rounds_sub_Sub_7_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_7_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .A2(Midori_rounds_sub_Sub_7_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_7_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_7_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .A2(Midori_rounds_sub_Sub_7_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_7_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq3[1]), .A2(Midori_rounds_sub_Sub_7_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_7_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_Rq1[3]), .B2(Midori_rounds_sub_Sub_7_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_7_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[3]), .A2(Midori_rounds_sub_Sub_7_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_7_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_Rq3[1]), .C2(Midori_rounds_sub_Sub_7_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_7_Rq1[3]), .B(
        Midori_rounds_sub_Sub_7_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq3[1]), .A2(Midori_rounds_sub_Sub_7_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_7_Rq2[2]), .A(
        Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_7_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_7_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_Rq3[1]), .C2(Midori_rounds_sub_Sub_7_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_7_Rq2[3]), .B(
        Midori_rounds_sub_Sub_7_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq3[1]), .A2(Midori_rounds_sub_Sub_7_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_7_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .C2(Midori_rounds_sub_Sub_7_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_7_Rq3[3]), .B(
        Midori_rounds_sub_Sub_7_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_7_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_Rq1[1]), .A2(Midori_rounds_sub_Sub_7_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_7_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_7_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_7_Rq3[2]), .A(
        Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_7_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_7_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[0])
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[0])
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[0])
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[11]), .ZN(Midori_rounds_SR_Result1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[14]), .ZN(Midori_rounds_SR_Result2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[17]), .ZN(Midori_rounds_SR_Result3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[20]), .ZN(Midori_rounds_SR_Result1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[23]), .ZN(Midori_rounds_SR_Result2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[26]), .ZN(Midori_rounds_SR_Result3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_7_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_7_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_8_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_8_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_8_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_8_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_8_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_8_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_8_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_8_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_8_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_8_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_8_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_8_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_8_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_8_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_8_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_8_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_8_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_8_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_8_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_8_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_8_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_8_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_8_InputAffine_U7 ( .A(Midori_rounds_n829), .ZN(
        Midori_rounds_sub_Sub_8_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_InputAffine_U6 ( .A(Midori_rounds_n949), .B(
        Midori_rounds_n951), .Z(Midori_rounds_sub_Sub_8_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_InputAffine_U5 ( .A(Midori_rounds_n949), .B(
        Midori_rounds_sub_Sub_8_F_in3[2]), .Z(Midori_rounds_sub_Sub_8_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_InputAffine_U4 ( .A(Midori_rounds_n885), .B(
        Midori_rounds_n887), .Z(Midori_rounds_sub_Sub_8_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_InputAffine_U3 ( .A(Midori_rounds_n885), .B(
        Midori_rounds_sub_Sub_8_F_in2[2]), .Z(Midori_rounds_sub_Sub_8_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_InputAffine_U2 ( .A(Midori_rounds_n797), 
        .B(Midori_rounds_n830), .ZN(Midori_rounds_sub_Sub_8_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_InputAffine_U1 ( .A(Midori_rounds_n797), .B(
        Midori_rounds_sub_Sub_8_F_in1[2]), .Z(Midori_rounds_sub_Sub_8_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U18 ( .A(Midori_rounds_sub_Sub_8_F_n12), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_8_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U17 ( .A(r[66]), .B(
        Midori_rounds_sub_Sub_8_F_q3[3]), .ZN(Midori_rounds_sub_Sub_8_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U16 ( .A(Midori_rounds_sub_Sub_8_F_n11), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_8_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U15 ( .A(r[64]), .B(
        Midori_rounds_sub_Sub_8_F_q3[2]), .ZN(Midori_rounds_sub_Sub_8_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U14 ( .A(Midori_rounds_sub_Sub_8_F_n10), 
        .B(r[71]), .ZN(Midori_rounds_sub_Sub_8_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U13 ( .A(r[70]), .B(
        Midori_rounds_sub_Sub_8_F_q3[1]), .ZN(Midori_rounds_sub_Sub_8_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U12 ( .A(Midori_rounds_sub_Sub_8_F_n9), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_8_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_U11 ( .A(r[68]), .B(
        Midori_rounds_sub_Sub_8_F_q3[0]), .ZN(Midori_rounds_sub_Sub_8_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U10 ( .A(r[67]), .B(
        Midori_rounds_sub_Sub_8_F_q2[3]), .Z(Midori_rounds_sub_Sub_8_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U9 ( .A(r[65]), .B(
        Midori_rounds_sub_Sub_8_F_q2[2]), .Z(Midori_rounds_sub_Sub_8_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U8 ( .A(r[71]), .B(
        Midori_rounds_sub_Sub_8_F_q2[1]), .Z(Midori_rounds_sub_Sub_8_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U7 ( .A(r[69]), .B(
        Midori_rounds_sub_Sub_8_F_q2[0]), .Z(Midori_rounds_sub_Sub_8_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U6 ( .A(r[66]), .B(
        Midori_rounds_sub_Sub_8_F_q1[3]), .Z(Midori_rounds_sub_Sub_8_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U5 ( .A(r[64]), .B(
        Midori_rounds_sub_Sub_8_F_q1[2]), .Z(Midori_rounds_sub_Sub_8_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U4 ( .A(r[70]), .B(
        Midori_rounds_sub_Sub_8_F_q1[1]), .Z(Midori_rounds_sub_Sub_8_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_8_F_U3 ( .A(r[68]), .B(
        Midori_rounds_sub_Sub_8_F_q1[0]), .Z(Midori_rounds_sub_Sub_8_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_8_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_8_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_8_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_8_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_8_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_8_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_8_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_8_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_8_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_8_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_8_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_8_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_8_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_8_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_8_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_8_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_8_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_8_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_8_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_8_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_8_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_8_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_8_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_8_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_8_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_8_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_8_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_8_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_8_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_8_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_8_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_8_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_8_G_U3 ( .A(Midori_rounds_sub_Sub_8_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_8_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_8_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_8_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_8_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_8_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_8_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_8_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .A2(Midori_rounds_sub_Sub_8_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_8_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[3]), .A2(Midori_rounds_sub_Sub_8_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_8_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_8_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .A2(Midori_rounds_sub_Sub_8_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_8_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .A2(Midori_rounds_sub_Sub_8_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_8_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq2[3]), .A2(Midori_rounds_sub_Sub_8_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_8_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_8_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_8_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_8_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq3[1]), .A2(Midori_rounds_sub_Sub_8_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .A2(Midori_rounds_sub_Sub_8_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_8_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .A2(Midori_rounds_sub_Sub_8_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_8_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[3]), .A2(Midori_rounds_sub_Sub_8_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_8_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_8_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .A2(Midori_rounds_sub_Sub_8_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_8_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .A2(Midori_rounds_sub_Sub_8_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_8_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_8_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .A2(Midori_rounds_sub_Sub_8_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_8_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_8_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq3[1]), .A2(Midori_rounds_sub_Sub_8_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_8_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_Rq1[3]), .B2(Midori_rounds_sub_Sub_8_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_8_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[3]), .A2(Midori_rounds_sub_Sub_8_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_8_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_8_Rq3[1]), .C2(Midori_rounds_sub_Sub_8_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_8_Rq1[3]), .B(
        Midori_rounds_sub_Sub_8_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq3[1]), .A2(Midori_rounds_sub_Sub_8_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_8_Rq2[2]), .A(
        Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_8_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_8_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_8_Rq3[1]), .C2(Midori_rounds_sub_Sub_8_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_8_Rq2[3]), .B(
        Midori_rounds_sub_Sub_8_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq3[1]), .A2(Midori_rounds_sub_Sub_8_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_8_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .C2(Midori_rounds_sub_Sub_8_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_8_Rq3[3]), .B(
        Midori_rounds_sub_Sub_8_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_8_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_8_Rq1[1]), .A2(Midori_rounds_sub_Sub_8_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_8_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_8_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_8_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_8_Rq3[2]), .A(
        Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_8_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_8_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_8_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_8_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[12]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[12]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[12]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[14]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[14]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[14]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[15]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[15]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[15]) );
  XNOR2_X1 Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_8_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_8_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_8_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq1_reg_3_ ( .D(Midori_rounds_sub_Sub_9_q1[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq1_reg_2_ ( .D(Midori_rounds_sub_Sub_9_q1[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq1_reg_1_ ( .D(Midori_rounds_sub_Sub_9_q1[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq1_reg_0_ ( .D(Midori_rounds_sub_Sub_9_q1[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq2_reg_3_ ( .D(Midori_rounds_sub_Sub_9_q2[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq2_reg_2_ ( .D(Midori_rounds_sub_Sub_9_q2[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq2_reg_1_ ( .D(Midori_rounds_sub_Sub_9_q2[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq2_reg_0_ ( .D(Midori_rounds_sub_Sub_9_q2[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq3_reg_3_ ( .D(Midori_rounds_sub_Sub_9_q3[3]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq3_reg_2_ ( .D(Midori_rounds_sub_Sub_9_q3[2]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq3_reg_1_ ( .D(Midori_rounds_sub_Sub_9_q3[1]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_Rq3_reg_0_ ( .D(Midori_rounds_sub_Sub_9_q3[0]), .CK(clk), .Q(Midori_rounds_sub_Sub_9_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_9_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_9_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_9_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_9_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_9_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_9_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_9_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_9_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_9_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_9_InputAffine_U7 ( .A(Midori_rounds_n832), .ZN(
        Midori_rounds_sub_Sub_9_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_InputAffine_U6 ( .A(Midori_rounds_n953), .B(
        Midori_rounds_n955), .Z(Midori_rounds_sub_Sub_9_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_InputAffine_U5 ( .A(Midori_rounds_n953), .B(
        Midori_rounds_sub_Sub_9_F_in3[2]), .Z(Midori_rounds_sub_Sub_9_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_InputAffine_U4 ( .A(Midori_rounds_n889), .B(
        Midori_rounds_n891), .Z(Midori_rounds_sub_Sub_9_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_InputAffine_U3 ( .A(Midori_rounds_n889), .B(
        Midori_rounds_sub_Sub_9_F_in2[2]), .Z(Midori_rounds_sub_Sub_9_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_InputAffine_U2 ( .A(Midori_rounds_n798), 
        .B(Midori_rounds_n833), .ZN(Midori_rounds_sub_Sub_9_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_InputAffine_U1 ( .A(Midori_rounds_n798), .B(
        Midori_rounds_sub_Sub_9_F_in1[2]), .Z(Midori_rounds_sub_Sub_9_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U18 ( .A(Midori_rounds_sub_Sub_9_F_n12), 
        .B(r[75]), .ZN(Midori_rounds_sub_Sub_9_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U17 ( .A(r[74]), .B(
        Midori_rounds_sub_Sub_9_F_q3[3]), .ZN(Midori_rounds_sub_Sub_9_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U16 ( .A(Midori_rounds_sub_Sub_9_F_n11), 
        .B(r[73]), .ZN(Midori_rounds_sub_Sub_9_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U15 ( .A(r[72]), .B(
        Midori_rounds_sub_Sub_9_F_q3[2]), .ZN(Midori_rounds_sub_Sub_9_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U14 ( .A(Midori_rounds_sub_Sub_9_F_n10), 
        .B(r[79]), .ZN(Midori_rounds_sub_Sub_9_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U13 ( .A(r[78]), .B(
        Midori_rounds_sub_Sub_9_F_q3[1]), .ZN(Midori_rounds_sub_Sub_9_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U12 ( .A(Midori_rounds_sub_Sub_9_F_n9), 
        .B(r[77]), .ZN(Midori_rounds_sub_Sub_9_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_U11 ( .A(r[76]), .B(
        Midori_rounds_sub_Sub_9_F_q3[0]), .ZN(Midori_rounds_sub_Sub_9_F_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U10 ( .A(r[75]), .B(
        Midori_rounds_sub_Sub_9_F_q2[3]), .Z(Midori_rounds_sub_Sub_9_q2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U9 ( .A(r[73]), .B(
        Midori_rounds_sub_Sub_9_F_q2[2]), .Z(Midori_rounds_sub_Sub_9_q2[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U8 ( .A(r[79]), .B(
        Midori_rounds_sub_Sub_9_F_q2[1]), .Z(Midori_rounds_sub_Sub_9_q2[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U7 ( .A(r[77]), .B(
        Midori_rounds_sub_Sub_9_F_q2[0]), .Z(Midori_rounds_sub_Sub_9_q2[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U6 ( .A(r[74]), .B(
        Midori_rounds_sub_Sub_9_F_q1[3]), .Z(Midori_rounds_sub_Sub_9_q1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U5 ( .A(r[72]), .B(
        Midori_rounds_sub_Sub_9_F_q1[2]), .Z(Midori_rounds_sub_Sub_9_q1[2]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U4 ( .A(r[78]), .B(
        Midori_rounds_sub_Sub_9_F_q1[1]), .Z(Midori_rounds_sub_Sub_9_q1[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_9_F_U3 ( .A(r[76]), .B(
        Midori_rounds_sub_Sub_9_F_q1[0]), .Z(Midori_rounds_sub_Sub_9_q1[0]) );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_9_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_9_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_9_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_9_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_9_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_9_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_9_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_9_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_9_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_9_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_9_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_9_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_9_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_9_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_9_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_9_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_9_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_9_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_9_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_9_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_9_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_9_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_9_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_9_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_9_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_9_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_9_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_9_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_9_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_9_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_9_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_9_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_9_G_U3 ( .A(Midori_rounds_sub_Sub_9_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_9_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_9_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_9_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_9_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_9_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_9_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_9_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .A2(Midori_rounds_sub_Sub_9_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_9_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[3]), .A2(Midori_rounds_sub_Sub_9_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_9_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_9_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .A2(Midori_rounds_sub_Sub_9_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_9_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .A2(Midori_rounds_sub_Sub_9_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_9_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq2[3]), .A2(Midori_rounds_sub_Sub_9_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_9_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_9_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_9_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_9_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq3[1]), .A2(Midori_rounds_sub_Sub_9_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .A2(Midori_rounds_sub_Sub_9_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_9_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .A2(Midori_rounds_sub_Sub_9_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_9_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[3]), .A2(Midori_rounds_sub_Sub_9_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_9_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_9_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .A2(Midori_rounds_sub_Sub_9_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_9_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .A2(Midori_rounds_sub_Sub_9_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_9_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_9_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .A2(Midori_rounds_sub_Sub_9_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_9_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_9_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq3[1]), .A2(Midori_rounds_sub_Sub_9_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_9_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_Rq1[3]), .B2(Midori_rounds_sub_Sub_9_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_9_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[3]), .A2(Midori_rounds_sub_Sub_9_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_9_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_9_Rq3[1]), .C2(Midori_rounds_sub_Sub_9_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_9_Rq1[3]), .B(
        Midori_rounds_sub_Sub_9_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq3[1]), .A2(Midori_rounds_sub_Sub_9_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_9_Rq2[2]), .A(
        Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_9_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_9_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_9_Rq3[1]), .C2(Midori_rounds_sub_Sub_9_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_9_Rq2[3]), .B(
        Midori_rounds_sub_Sub_9_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq3[1]), .A2(Midori_rounds_sub_Sub_9_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_9_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .C2(Midori_rounds_sub_Sub_9_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_9_Rq3[3]), .B(
        Midori_rounds_sub_Sub_9_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_9_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_9_Rq1[1]), .A2(Midori_rounds_sub_Sub_9_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_9_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_9_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_9_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_9_Rq3[2]), .A(
        Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_9_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_9_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_9_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_9_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[18]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[18]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[18]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_9_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_9_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_9_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq1_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_q1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq1_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_q1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_q1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq1_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_q1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq2_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_q2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq2_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_q2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_q2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq2_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_q2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq3_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_q3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq3_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_q3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_q3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_Rq3_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_q3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_10_InputAffine_U7 ( .A(Midori_rounds_n835), 
        .ZN(Midori_rounds_sub_Sub_10_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_10_InputAffine_U6 ( .A(Midori_rounds_n957), 
        .B(Midori_rounds_n959), .Z(Midori_rounds_sub_Sub_10_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_10_InputAffine_U5 ( .A(Midori_rounds_n957), 
        .B(Midori_rounds_sub_Sub_10_F_in3[2]), .Z(
        Midori_rounds_sub_Sub_10_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_10_InputAffine_U4 ( .A(Midori_rounds_n893), 
        .B(Midori_rounds_n895), .Z(Midori_rounds_sub_Sub_10_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_10_InputAffine_U3 ( .A(Midori_rounds_n893), 
        .B(Midori_rounds_sub_Sub_10_F_in2[2]), .Z(
        Midori_rounds_sub_Sub_10_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_InputAffine_U2 ( .A(Midori_rounds_n799), 
        .B(Midori_rounds_n836), .ZN(Midori_rounds_sub_Sub_10_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_10_InputAffine_U1 ( .A(Midori_rounds_n799), 
        .B(Midori_rounds_sub_Sub_10_F_in1[2]), .Z(
        Midori_rounds_sub_Sub_10_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U18 ( .A(Midori_rounds_sub_Sub_10_F_n12), 
        .B(r[83]), .ZN(Midori_rounds_sub_Sub_10_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U17 ( .A(r[82]), .B(
        Midori_rounds_sub_Sub_10_F_q3[3]), .ZN(Midori_rounds_sub_Sub_10_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U16 ( .A(Midori_rounds_sub_Sub_10_F_n11), 
        .B(r[81]), .ZN(Midori_rounds_sub_Sub_10_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U15 ( .A(r[80]), .B(
        Midori_rounds_sub_Sub_10_F_q3[2]), .ZN(Midori_rounds_sub_Sub_10_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U14 ( .A(Midori_rounds_sub_Sub_10_F_n10), 
        .B(r[87]), .ZN(Midori_rounds_sub_Sub_10_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U13 ( .A(r[86]), .B(
        Midori_rounds_sub_Sub_10_F_q3[1]), .ZN(Midori_rounds_sub_Sub_10_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U12 ( .A(Midori_rounds_sub_Sub_10_F_n9), 
        .B(r[85]), .ZN(Midori_rounds_sub_Sub_10_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_U11 ( .A(r[84]), .B(
        Midori_rounds_sub_Sub_10_F_q3[0]), .ZN(Midori_rounds_sub_Sub_10_F_n9)
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U10 ( .A(r[83]), .B(
        Midori_rounds_sub_Sub_10_F_q2[3]), .Z(Midori_rounds_sub_Sub_10_q2[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U9 ( .A(r[81]), .B(
        Midori_rounds_sub_Sub_10_F_q2[2]), .Z(Midori_rounds_sub_Sub_10_q2[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U8 ( .A(r[87]), .B(
        Midori_rounds_sub_Sub_10_F_q2[1]), .Z(Midori_rounds_sub_Sub_10_q2[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U7 ( .A(r[85]), .B(
        Midori_rounds_sub_Sub_10_F_q2[0]), .Z(Midori_rounds_sub_Sub_10_q2[0])
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U6 ( .A(r[82]), .B(
        Midori_rounds_sub_Sub_10_F_q1[3]), .Z(Midori_rounds_sub_Sub_10_q1[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U5 ( .A(r[80]), .B(
        Midori_rounds_sub_Sub_10_F_q1[2]), .Z(Midori_rounds_sub_Sub_10_q1[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U4 ( .A(r[86]), .B(
        Midori_rounds_sub_Sub_10_F_q1[1]), .Z(Midori_rounds_sub_Sub_10_q1[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_10_F_U3 ( .A(r[84]), .B(
        Midori_rounds_sub_Sub_10_F_q1[0]), .Z(Midori_rounds_sub_Sub_10_q1[0])
         );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_10_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_10_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_10_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_10_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_10_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_10_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_10_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_10_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_10_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_10_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_10_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_10_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_10_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_10_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_10_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_10_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_10_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_10_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_10_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_10_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_10_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_10_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_10_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_10_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_10_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_10_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_10_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_10_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_10_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_10_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_10_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_10_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_10_G_U3 ( .A(Midori_rounds_sub_Sub_10_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_10_G_n2) );
  DFF_X1 Midori_rounds_sub_Sub_10_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[53]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[53]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_G_n2), .CK(clk), .Q(
        Midori_rounds_SR_Result1[53]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_10_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_10_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_10_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_10_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_10_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .A2(Midori_rounds_sub_Sub_10_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_10_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[3]), .A2(Midori_rounds_sub_Sub_10_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_10_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_10_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .A2(Midori_rounds_sub_Sub_10_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_10_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .A2(Midori_rounds_sub_Sub_10_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_10_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq2[3]), .A2(Midori_rounds_sub_Sub_10_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_10_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_10_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_10_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_10_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq3[1]), .A2(Midori_rounds_sub_Sub_10_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .A2(Midori_rounds_sub_Sub_10_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_10_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .A2(Midori_rounds_sub_Sub_10_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_10_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[3]), .A2(Midori_rounds_sub_Sub_10_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_10_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_10_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .A2(Midori_rounds_sub_Sub_10_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_10_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .A2(Midori_rounds_sub_Sub_10_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_10_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_10_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .A2(Midori_rounds_sub_Sub_10_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_10_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_10_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq3[1]), .A2(Midori_rounds_sub_Sub_10_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_10_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_Rq1[3]), .B2(Midori_rounds_sub_Sub_10_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_10_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[3]), .A2(Midori_rounds_sub_Sub_10_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_10_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_10_Rq3[1]), .C2(Midori_rounds_sub_Sub_10_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_10_Rq1[3]), .B(
        Midori_rounds_sub_Sub_10_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq3[1]), .A2(Midori_rounds_sub_Sub_10_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_10_Rq2[2]), .A(
        Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_10_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_10_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_10_Rq3[1]), .C2(Midori_rounds_sub_Sub_10_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_10_Rq2[3]), .B(
        Midori_rounds_sub_Sub_10_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq3[1]), .A2(Midori_rounds_sub_Sub_10_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_10_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .C2(Midori_rounds_sub_Sub_10_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_10_Rq3[3]), .B(
        Midori_rounds_sub_Sub_10_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_10_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_10_Rq1[1]), .A2(Midori_rounds_sub_Sub_10_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_10_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_10_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_10_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_10_Rq3[2]), .A(
        Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_10_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_10_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_10_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_10_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[52]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[52]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[52]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[54]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[54]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[54]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[55]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[55]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[55]) );
  XNOR2_X1 Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_10_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_10_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_10_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq1_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_q1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq1_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_q1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_q1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq1_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_q1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq2_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_q2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq2_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_q2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_q2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq2_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_q2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq3_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_q3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq3_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_q3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_q3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_Rq3_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_q3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_11_InputAffine_U7 ( .A(Midori_rounds_n838), 
        .ZN(Midori_rounds_sub_Sub_11_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_11_InputAffine_U6 ( .A(Midori_rounds_n961), 
        .B(Midori_rounds_n963), .Z(Midori_rounds_sub_Sub_11_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_11_InputAffine_U5 ( .A(Midori_rounds_n961), 
        .B(Midori_rounds_sub_Sub_11_F_in3[2]), .Z(
        Midori_rounds_sub_Sub_11_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_11_InputAffine_U4 ( .A(Midori_rounds_n897), 
        .B(Midori_rounds_n899), .Z(Midori_rounds_sub_Sub_11_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_11_InputAffine_U3 ( .A(Midori_rounds_n897), 
        .B(Midori_rounds_sub_Sub_11_F_in2[2]), .Z(
        Midori_rounds_sub_Sub_11_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_InputAffine_U2 ( .A(Midori_rounds_n800), 
        .B(Midori_rounds_n839), .ZN(Midori_rounds_sub_Sub_11_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_11_InputAffine_U1 ( .A(Midori_rounds_n800), 
        .B(Midori_rounds_sub_Sub_11_F_in1[2]), .Z(
        Midori_rounds_sub_Sub_11_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U18 ( .A(Midori_rounds_sub_Sub_11_F_n12), 
        .B(r[91]), .ZN(Midori_rounds_sub_Sub_11_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U17 ( .A(r[90]), .B(
        Midori_rounds_sub_Sub_11_F_q3[3]), .ZN(Midori_rounds_sub_Sub_11_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U16 ( .A(Midori_rounds_sub_Sub_11_F_n11), 
        .B(r[89]), .ZN(Midori_rounds_sub_Sub_11_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U15 ( .A(r[88]), .B(
        Midori_rounds_sub_Sub_11_F_q3[2]), .ZN(Midori_rounds_sub_Sub_11_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U14 ( .A(Midori_rounds_sub_Sub_11_F_n10), 
        .B(r[95]), .ZN(Midori_rounds_sub_Sub_11_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U13 ( .A(r[94]), .B(
        Midori_rounds_sub_Sub_11_F_q3[1]), .ZN(Midori_rounds_sub_Sub_11_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U12 ( .A(Midori_rounds_sub_Sub_11_F_n9), 
        .B(r[93]), .ZN(Midori_rounds_sub_Sub_11_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_U11 ( .A(r[92]), .B(
        Midori_rounds_sub_Sub_11_F_q3[0]), .ZN(Midori_rounds_sub_Sub_11_F_n9)
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U10 ( .A(r[91]), .B(
        Midori_rounds_sub_Sub_11_F_q2[3]), .Z(Midori_rounds_sub_Sub_11_q2[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U9 ( .A(r[89]), .B(
        Midori_rounds_sub_Sub_11_F_q2[2]), .Z(Midori_rounds_sub_Sub_11_q2[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U8 ( .A(r[95]), .B(
        Midori_rounds_sub_Sub_11_F_q2[1]), .Z(Midori_rounds_sub_Sub_11_q2[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U7 ( .A(r[93]), .B(
        Midori_rounds_sub_Sub_11_F_q2[0]), .Z(Midori_rounds_sub_Sub_11_q2[0])
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U6 ( .A(r[90]), .B(
        Midori_rounds_sub_Sub_11_F_q1[3]), .Z(Midori_rounds_sub_Sub_11_q1[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U5 ( .A(r[88]), .B(
        Midori_rounds_sub_Sub_11_F_q1[2]), .Z(Midori_rounds_sub_Sub_11_q1[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U4 ( .A(r[94]), .B(
        Midori_rounds_sub_Sub_11_F_q1[1]), .Z(Midori_rounds_sub_Sub_11_q1[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_11_F_U3 ( .A(r[92]), .B(
        Midori_rounds_sub_Sub_11_F_q1[0]), .Z(Midori_rounds_sub_Sub_11_q1[0])
         );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_11_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_11_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_11_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_11_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_11_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_11_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_11_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_11_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_11_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_11_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_11_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_11_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_11_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_11_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_11_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_11_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_11_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_11_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_11_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_11_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_11_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_11_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_11_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_11_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_11_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_11_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_11_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_11_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_11_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_11_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_11_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_11_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_11_G_U3 ( .A(Midori_rounds_sub_Sub_11_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_11_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_11_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[41]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[41]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[41]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_11_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_11_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_11_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_11_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_11_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .A2(Midori_rounds_sub_Sub_11_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_11_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[3]), .A2(Midori_rounds_sub_Sub_11_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_11_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_11_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .A2(Midori_rounds_sub_Sub_11_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_11_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .A2(Midori_rounds_sub_Sub_11_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_11_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq2[3]), .A2(Midori_rounds_sub_Sub_11_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_11_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_11_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_11_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_11_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq3[1]), .A2(Midori_rounds_sub_Sub_11_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .A2(Midori_rounds_sub_Sub_11_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_11_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .A2(Midori_rounds_sub_Sub_11_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_11_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[3]), .A2(Midori_rounds_sub_Sub_11_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_11_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_11_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .A2(Midori_rounds_sub_Sub_11_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_11_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .A2(Midori_rounds_sub_Sub_11_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_11_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_11_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .A2(Midori_rounds_sub_Sub_11_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_11_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_11_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq3[1]), .A2(Midori_rounds_sub_Sub_11_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_11_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_Rq1[3]), .B2(Midori_rounds_sub_Sub_11_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_11_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[3]), .A2(Midori_rounds_sub_Sub_11_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_11_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_11_Rq3[1]), .C2(Midori_rounds_sub_Sub_11_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_11_Rq1[3]), .B(
        Midori_rounds_sub_Sub_11_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq3[1]), .A2(Midori_rounds_sub_Sub_11_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_11_Rq2[2]), .A(
        Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_11_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_11_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_11_Rq3[1]), .C2(Midori_rounds_sub_Sub_11_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_11_Rq2[3]), .B(
        Midori_rounds_sub_Sub_11_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq3[1]), .A2(Midori_rounds_sub_Sub_11_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_11_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .C2(Midori_rounds_sub_Sub_11_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_11_Rq3[3]), .B(
        Midori_rounds_sub_Sub_11_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_11_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_11_Rq1[1]), .A2(Midori_rounds_sub_Sub_11_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_11_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_11_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_11_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_11_Rq3[2]), .A(
        Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_11_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_11_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_11_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_11_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[40]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[40]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[40]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[42]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[42]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[42]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[43]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[43]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[43]) );
  XNOR2_X1 Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_11_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_11_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_11_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq1_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_q1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq1_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_q1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_q1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq1_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_q1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq2_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_q2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq2_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_q2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_q2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq2_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_q2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq3_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_q3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq3_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_q3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_q3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_Rq3_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_q3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_12_InputAffine_U7 ( .A(Midori_rounds_n841), 
        .ZN(Midori_rounds_sub_Sub_12_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_12_InputAffine_U6 ( .A(Midori_rounds_n965), 
        .B(Midori_rounds_n967), .Z(Midori_rounds_sub_Sub_12_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_12_InputAffine_U5 ( .A(Midori_rounds_n965), 
        .B(Midori_rounds_sub_Sub_12_F_in3[2]), .Z(
        Midori_rounds_sub_Sub_12_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_12_InputAffine_U4 ( .A(Midori_rounds_n901), 
        .B(Midori_rounds_n903), .Z(Midori_rounds_sub_Sub_12_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_12_InputAffine_U3 ( .A(Midori_rounds_n901), 
        .B(Midori_rounds_sub_Sub_12_F_in2[2]), .Z(
        Midori_rounds_sub_Sub_12_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_InputAffine_U2 ( .A(Midori_rounds_n801), 
        .B(Midori_rounds_n842), .ZN(Midori_rounds_sub_Sub_12_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_12_InputAffine_U1 ( .A(Midori_rounds_n801), 
        .B(Midori_rounds_sub_Sub_12_F_in1[2]), .Z(
        Midori_rounds_sub_Sub_12_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U18 ( .A(Midori_rounds_sub_Sub_12_F_n12), 
        .B(r[99]), .ZN(Midori_rounds_sub_Sub_12_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U17 ( .A(r[98]), .B(
        Midori_rounds_sub_Sub_12_F_q3[3]), .ZN(Midori_rounds_sub_Sub_12_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U16 ( .A(Midori_rounds_sub_Sub_12_F_n11), 
        .B(r[97]), .ZN(Midori_rounds_sub_Sub_12_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U15 ( .A(r[96]), .B(
        Midori_rounds_sub_Sub_12_F_q3[2]), .ZN(Midori_rounds_sub_Sub_12_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U14 ( .A(Midori_rounds_sub_Sub_12_F_n10), 
        .B(r[103]), .ZN(Midori_rounds_sub_Sub_12_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U13 ( .A(r[102]), .B(
        Midori_rounds_sub_Sub_12_F_q3[1]), .ZN(Midori_rounds_sub_Sub_12_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U12 ( .A(Midori_rounds_sub_Sub_12_F_n9), 
        .B(r[101]), .ZN(Midori_rounds_sub_Sub_12_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_U11 ( .A(r[100]), .B(
        Midori_rounds_sub_Sub_12_F_q3[0]), .ZN(Midori_rounds_sub_Sub_12_F_n9)
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U10 ( .A(r[99]), .B(
        Midori_rounds_sub_Sub_12_F_q2[3]), .Z(Midori_rounds_sub_Sub_12_q2[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U9 ( .A(r[97]), .B(
        Midori_rounds_sub_Sub_12_F_q2[2]), .Z(Midori_rounds_sub_Sub_12_q2[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U8 ( .A(r[103]), .B(
        Midori_rounds_sub_Sub_12_F_q2[1]), .Z(Midori_rounds_sub_Sub_12_q2[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U7 ( .A(r[101]), .B(
        Midori_rounds_sub_Sub_12_F_q2[0]), .Z(Midori_rounds_sub_Sub_12_q2[0])
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U6 ( .A(r[98]), .B(
        Midori_rounds_sub_Sub_12_F_q1[3]), .Z(Midori_rounds_sub_Sub_12_q1[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U5 ( .A(r[96]), .B(
        Midori_rounds_sub_Sub_12_F_q1[2]), .Z(Midori_rounds_sub_Sub_12_q1[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U4 ( .A(r[102]), .B(
        Midori_rounds_sub_Sub_12_F_q1[1]), .Z(Midori_rounds_sub_Sub_12_q1[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_12_F_U3 ( .A(r[100]), .B(
        Midori_rounds_sub_Sub_12_F_q1[0]), .Z(Midori_rounds_sub_Sub_12_q1[0])
         );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_12_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_12_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_12_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_12_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_12_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_12_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_12_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_12_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_12_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_12_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_12_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_12_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_12_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_12_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_12_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_12_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_12_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_12_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_12_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_12_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_12_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_12_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_12_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_12_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_12_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_12_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_12_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_12_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_12_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_12_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_12_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_12_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_12_G_U3 ( .A(Midori_rounds_sub_Sub_12_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_12_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_12_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_12_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_12_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_12_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_12_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_12_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .A2(Midori_rounds_sub_Sub_12_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_12_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[3]), .A2(Midori_rounds_sub_Sub_12_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_12_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_12_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .A2(Midori_rounds_sub_Sub_12_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_12_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .A2(Midori_rounds_sub_Sub_12_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_12_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq2[3]), .A2(Midori_rounds_sub_Sub_12_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_12_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_12_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_12_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_12_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq3[1]), .A2(Midori_rounds_sub_Sub_12_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .A2(Midori_rounds_sub_Sub_12_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_12_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .A2(Midori_rounds_sub_Sub_12_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_12_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[3]), .A2(Midori_rounds_sub_Sub_12_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_12_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_12_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .A2(Midori_rounds_sub_Sub_12_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_12_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .A2(Midori_rounds_sub_Sub_12_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_12_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_12_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .A2(Midori_rounds_sub_Sub_12_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_12_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_12_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq3[1]), .A2(Midori_rounds_sub_Sub_12_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_12_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_Rq1[3]), .B2(Midori_rounds_sub_Sub_12_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_12_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[3]), .A2(Midori_rounds_sub_Sub_12_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_12_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_12_Rq3[1]), .C2(Midori_rounds_sub_Sub_12_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_12_Rq1[3]), .B(
        Midori_rounds_sub_Sub_12_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq3[1]), .A2(Midori_rounds_sub_Sub_12_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_12_Rq2[2]), .A(
        Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_12_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_12_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_12_Rq3[1]), .C2(Midori_rounds_sub_Sub_12_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_12_Rq2[3]), .B(
        Midori_rounds_sub_Sub_12_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq3[1]), .A2(Midori_rounds_sub_Sub_12_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_12_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .C2(Midori_rounds_sub_Sub_12_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_12_Rq3[3]), .B(
        Midori_rounds_sub_Sub_12_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_12_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_12_Rq1[1]), .A2(Midori_rounds_sub_Sub_12_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_12_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_12_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_12_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_12_Rq3[2]), .A(
        Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_12_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_12_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_12_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_12_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[24]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[24]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[24]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[27]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[27]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[27]) );
  XNOR2_X1 Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_12_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_12_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_12_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq1_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_q1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq1_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_q1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_q1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq1_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_q1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq2_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_q2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq2_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_q2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_q2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq2_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_q2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq3_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_q3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq3_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_q3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_q3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_Rq3_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_q3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_13_InputAffine_U7 ( .A(Midori_rounds_n844), 
        .ZN(Midori_rounds_sub_Sub_13_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_13_InputAffine_U6 ( .A(Midori_rounds_n969), 
        .B(Midori_rounds_n971), .Z(Midori_rounds_sub_Sub_13_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_13_InputAffine_U5 ( .A(Midori_rounds_n969), 
        .B(Midori_rounds_sub_Sub_13_F_in3[2]), .Z(
        Midori_rounds_sub_Sub_13_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_13_InputAffine_U4 ( .A(Midori_rounds_n905), 
        .B(Midori_rounds_n907), .Z(Midori_rounds_sub_Sub_13_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_13_InputAffine_U3 ( .A(Midori_rounds_n905), 
        .B(Midori_rounds_sub_Sub_13_F_in2[2]), .Z(
        Midori_rounds_sub_Sub_13_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_InputAffine_U2 ( .A(Midori_rounds_n802), 
        .B(Midori_rounds_n845), .ZN(Midori_rounds_sub_Sub_13_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_13_InputAffine_U1 ( .A(Midori_rounds_n802), 
        .B(Midori_rounds_sub_Sub_13_F_in1[2]), .Z(
        Midori_rounds_sub_Sub_13_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U18 ( .A(Midori_rounds_sub_Sub_13_F_n12), 
        .B(r[107]), .ZN(Midori_rounds_sub_Sub_13_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U17 ( .A(r[106]), .B(
        Midori_rounds_sub_Sub_13_F_q3[3]), .ZN(Midori_rounds_sub_Sub_13_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U16 ( .A(Midori_rounds_sub_Sub_13_F_n11), 
        .B(r[105]), .ZN(Midori_rounds_sub_Sub_13_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U15 ( .A(r[104]), .B(
        Midori_rounds_sub_Sub_13_F_q3[2]), .ZN(Midori_rounds_sub_Sub_13_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U14 ( .A(Midori_rounds_sub_Sub_13_F_n10), 
        .B(r[111]), .ZN(Midori_rounds_sub_Sub_13_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U13 ( .A(r[110]), .B(
        Midori_rounds_sub_Sub_13_F_q3[1]), .ZN(Midori_rounds_sub_Sub_13_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U12 ( .A(Midori_rounds_sub_Sub_13_F_n9), 
        .B(r[109]), .ZN(Midori_rounds_sub_Sub_13_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_U11 ( .A(r[108]), .B(
        Midori_rounds_sub_Sub_13_F_q3[0]), .ZN(Midori_rounds_sub_Sub_13_F_n9)
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U10 ( .A(r[107]), .B(
        Midori_rounds_sub_Sub_13_F_q2[3]), .Z(Midori_rounds_sub_Sub_13_q2[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U9 ( .A(r[105]), .B(
        Midori_rounds_sub_Sub_13_F_q2[2]), .Z(Midori_rounds_sub_Sub_13_q2[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U8 ( .A(r[111]), .B(
        Midori_rounds_sub_Sub_13_F_q2[1]), .Z(Midori_rounds_sub_Sub_13_q2[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U7 ( .A(r[109]), .B(
        Midori_rounds_sub_Sub_13_F_q2[0]), .Z(Midori_rounds_sub_Sub_13_q2[0])
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U6 ( .A(r[106]), .B(
        Midori_rounds_sub_Sub_13_F_q1[3]), .Z(Midori_rounds_sub_Sub_13_q1[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U5 ( .A(r[104]), .B(
        Midori_rounds_sub_Sub_13_F_q1[2]), .Z(Midori_rounds_sub_Sub_13_q1[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U4 ( .A(r[110]), .B(
        Midori_rounds_sub_Sub_13_F_q1[1]), .Z(Midori_rounds_sub_Sub_13_q1[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_13_F_U3 ( .A(r[108]), .B(
        Midori_rounds_sub_Sub_13_F_q1[0]), .Z(Midori_rounds_sub_Sub_13_q1[0])
         );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_13_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_13_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_13_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_13_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_13_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_13_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_13_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_13_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_13_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_13_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_13_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_13_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_13_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_13_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_13_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_13_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_13_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_13_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_13_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_13_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_13_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_13_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_13_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_13_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_13_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_13_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_13_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_13_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_13_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_13_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_13_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_13_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_13_G_U3 ( .A(Midori_rounds_sub_Sub_13_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_13_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_13_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_13_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_13_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_13_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_13_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_13_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .A2(Midori_rounds_sub_Sub_13_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_13_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[3]), .A2(Midori_rounds_sub_Sub_13_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_13_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_13_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .A2(Midori_rounds_sub_Sub_13_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_13_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .A2(Midori_rounds_sub_Sub_13_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_13_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq2[3]), .A2(Midori_rounds_sub_Sub_13_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_13_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_13_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_13_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_13_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq3[1]), .A2(Midori_rounds_sub_Sub_13_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .A2(Midori_rounds_sub_Sub_13_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_13_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .A2(Midori_rounds_sub_Sub_13_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_13_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[3]), .A2(Midori_rounds_sub_Sub_13_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_13_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_13_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .A2(Midori_rounds_sub_Sub_13_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_13_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .A2(Midori_rounds_sub_Sub_13_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_13_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_13_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .A2(Midori_rounds_sub_Sub_13_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_13_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_13_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq3[1]), .A2(Midori_rounds_sub_Sub_13_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_13_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_Rq1[3]), .B2(Midori_rounds_sub_Sub_13_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_13_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[3]), .A2(Midori_rounds_sub_Sub_13_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_13_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_13_Rq3[1]), .C2(Midori_rounds_sub_Sub_13_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_13_Rq1[3]), .B(
        Midori_rounds_sub_Sub_13_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq3[1]), .A2(Midori_rounds_sub_Sub_13_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_13_Rq2[2]), .A(
        Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_13_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_13_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_13_Rq3[1]), .C2(Midori_rounds_sub_Sub_13_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_13_Rq2[3]), .B(
        Midori_rounds_sub_Sub_13_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq3[1]), .A2(Midori_rounds_sub_Sub_13_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_13_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .C2(Midori_rounds_sub_Sub_13_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_13_Rq3[3]), .B(
        Midori_rounds_sub_Sub_13_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_13_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_13_Rq1[1]), .A2(Midori_rounds_sub_Sub_13_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_13_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_13_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_13_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_13_Rq3[2]), .A(
        Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_13_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_13_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_13_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_13_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[2]), .ZN(Midori_rounds_SR_Result1[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[5]), .ZN(Midori_rounds_SR_Result2[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[8]), .ZN(Midori_rounds_SR_Result3[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[6]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[6]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[6]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_13_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_13_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_13_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq1_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_q1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq1_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_q1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_q1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq1_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_q1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq2_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_q2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq2_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_q2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_q2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq2_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_q2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq3_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_q3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq3_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_q3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_q3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_Rq3_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_q3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_14_InputAffine_U7 ( .A(Midori_rounds_n847), 
        .ZN(Midori_rounds_sub_Sub_14_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_14_InputAffine_U6 ( .A(Midori_rounds_n973), 
        .B(Midori_rounds_n975), .Z(Midori_rounds_sub_Sub_14_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_14_InputAffine_U5 ( .A(Midori_rounds_n973), 
        .B(Midori_rounds_sub_Sub_14_F_in3[2]), .Z(
        Midori_rounds_sub_Sub_14_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_14_InputAffine_U4 ( .A(Midori_rounds_n909), 
        .B(Midori_rounds_n911), .Z(Midori_rounds_sub_Sub_14_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_14_InputAffine_U3 ( .A(Midori_rounds_n909), 
        .B(Midori_rounds_sub_Sub_14_F_in2[2]), .Z(
        Midori_rounds_sub_Sub_14_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_InputAffine_U2 ( .A(Midori_rounds_n803), 
        .B(Midori_rounds_n848), .ZN(Midori_rounds_sub_Sub_14_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_14_InputAffine_U1 ( .A(Midori_rounds_n803), 
        .B(Midori_rounds_sub_Sub_14_F_in1[2]), .Z(
        Midori_rounds_sub_Sub_14_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U18 ( .A(Midori_rounds_sub_Sub_14_F_n12), 
        .B(r[115]), .ZN(Midori_rounds_sub_Sub_14_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U17 ( .A(r[114]), .B(
        Midori_rounds_sub_Sub_14_F_q3[3]), .ZN(Midori_rounds_sub_Sub_14_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U16 ( .A(Midori_rounds_sub_Sub_14_F_n11), 
        .B(r[113]), .ZN(Midori_rounds_sub_Sub_14_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U15 ( .A(r[112]), .B(
        Midori_rounds_sub_Sub_14_F_q3[2]), .ZN(Midori_rounds_sub_Sub_14_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U14 ( .A(Midori_rounds_sub_Sub_14_F_n10), 
        .B(r[119]), .ZN(Midori_rounds_sub_Sub_14_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U13 ( .A(r[118]), .B(
        Midori_rounds_sub_Sub_14_F_q3[1]), .ZN(Midori_rounds_sub_Sub_14_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U12 ( .A(Midori_rounds_sub_Sub_14_F_n9), 
        .B(r[117]), .ZN(Midori_rounds_sub_Sub_14_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_U11 ( .A(r[116]), .B(
        Midori_rounds_sub_Sub_14_F_q3[0]), .ZN(Midori_rounds_sub_Sub_14_F_n9)
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U10 ( .A(r[115]), .B(
        Midori_rounds_sub_Sub_14_F_q2[3]), .Z(Midori_rounds_sub_Sub_14_q2[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U9 ( .A(r[113]), .B(
        Midori_rounds_sub_Sub_14_F_q2[2]), .Z(Midori_rounds_sub_Sub_14_q2[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U8 ( .A(r[119]), .B(
        Midori_rounds_sub_Sub_14_F_q2[1]), .Z(Midori_rounds_sub_Sub_14_q2[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U7 ( .A(r[117]), .B(
        Midori_rounds_sub_Sub_14_F_q2[0]), .Z(Midori_rounds_sub_Sub_14_q2[0])
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U6 ( .A(r[114]), .B(
        Midori_rounds_sub_Sub_14_F_q1[3]), .Z(Midori_rounds_sub_Sub_14_q1[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U5 ( .A(r[112]), .B(
        Midori_rounds_sub_Sub_14_F_q1[2]), .Z(Midori_rounds_sub_Sub_14_q1[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U4 ( .A(r[118]), .B(
        Midori_rounds_sub_Sub_14_F_q1[1]), .Z(Midori_rounds_sub_Sub_14_q1[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_14_F_U3 ( .A(r[116]), .B(
        Midori_rounds_sub_Sub_14_F_q1[0]), .Z(Midori_rounds_sub_Sub_14_q1[0])
         );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_14_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_14_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_14_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_14_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_14_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_14_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_14_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_14_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_14_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_14_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_14_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_14_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_14_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_14_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_14_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_14_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_14_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_14_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_14_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_14_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_14_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_14_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_14_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_14_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_14_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_14_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_14_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_14_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_14_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_14_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_14_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_14_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_14_G_U3 ( .A(Midori_rounds_sub_Sub_14_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_14_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_14_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_14_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_14_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_14_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_14_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_14_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .A2(Midori_rounds_sub_Sub_14_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_14_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[3]), .A2(Midori_rounds_sub_Sub_14_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_14_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_14_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .A2(Midori_rounds_sub_Sub_14_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_14_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .A2(Midori_rounds_sub_Sub_14_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_14_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq2[3]), .A2(Midori_rounds_sub_Sub_14_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_14_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_14_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_14_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_14_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq3[1]), .A2(Midori_rounds_sub_Sub_14_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .A2(Midori_rounds_sub_Sub_14_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_14_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .A2(Midori_rounds_sub_Sub_14_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_14_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[3]), .A2(Midori_rounds_sub_Sub_14_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_14_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_14_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .A2(Midori_rounds_sub_Sub_14_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_14_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .A2(Midori_rounds_sub_Sub_14_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_14_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_14_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .A2(Midori_rounds_sub_Sub_14_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_14_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_14_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq3[1]), .A2(Midori_rounds_sub_Sub_14_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_14_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_Rq1[3]), .B2(Midori_rounds_sub_Sub_14_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_14_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[3]), .A2(Midori_rounds_sub_Sub_14_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_14_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_14_Rq3[1]), .C2(Midori_rounds_sub_Sub_14_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_14_Rq1[3]), .B(
        Midori_rounds_sub_Sub_14_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq3[1]), .A2(Midori_rounds_sub_Sub_14_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_14_Rq2[2]), .A(
        Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_14_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_14_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_14_Rq3[1]), .C2(Midori_rounds_sub_Sub_14_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_14_Rq2[3]), .B(
        Midori_rounds_sub_Sub_14_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq3[1]), .A2(Midori_rounds_sub_Sub_14_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_14_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .C2(Midori_rounds_sub_Sub_14_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_14_Rq3[3]), .B(
        Midori_rounds_sub_Sub_14_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_14_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_14_Rq1[1]), .A2(Midori_rounds_sub_Sub_14_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_14_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_14_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_14_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_14_Rq3[2]), .A(
        Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_14_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_14_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_14_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_14_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[32]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[32]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[32]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[34]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[34]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[34]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[35]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[35]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[35]) );
  XNOR2_X1 Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_14_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_14_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_14_G_InstXOR2_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq1_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_q1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq1_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_q1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_q1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq1_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_q1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq2_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_q2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq2_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_q2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_q2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq2_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_q2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq3_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_q3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq3[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq3_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_q3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_q3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_Rq3_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_q3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_Rq3[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_F_in3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_F_in3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_F_in3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_F_in3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_F_in2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in2_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_F_in2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_F_in2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_F_in2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_F_in1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in1_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_F_in1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_F_in1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_in1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_F_in1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .QN() );
  INV_X1 Midori_rounds_sub_Sub_15_InputAffine_U7 ( .A(Midori_rounds_n850), 
        .ZN(Midori_rounds_sub_Sub_15_F_in1[0]) );
  XOR2_X1 Midori_rounds_sub_Sub_15_InputAffine_U6 ( .A(Midori_rounds_n977), 
        .B(Midori_rounds_n979), .Z(Midori_rounds_sub_Sub_15_F_in3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_15_InputAffine_U5 ( .A(Midori_rounds_n977), 
        .B(Midori_rounds_sub_Sub_15_F_in3[2]), .Z(
        Midori_rounds_sub_Sub_15_F_in3[1]) );
  XOR2_X1 Midori_rounds_sub_Sub_15_InputAffine_U4 ( .A(Midori_rounds_n913), 
        .B(Midori_rounds_n915), .Z(Midori_rounds_sub_Sub_15_F_in2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_15_InputAffine_U3 ( .A(Midori_rounds_n913), 
        .B(Midori_rounds_sub_Sub_15_F_in2[2]), .Z(
        Midori_rounds_sub_Sub_15_F_in2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_InputAffine_U2 ( .A(Midori_rounds_n804), 
        .B(Midori_rounds_n851), .ZN(Midori_rounds_sub_Sub_15_F_in1[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_15_InputAffine_U1 ( .A(Midori_rounds_n804), 
        .B(Midori_rounds_sub_Sub_15_F_in1[2]), .Z(
        Midori_rounds_sub_Sub_15_F_in1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U18 ( .A(Midori_rounds_sub_Sub_15_F_n12), 
        .B(r[123]), .ZN(Midori_rounds_sub_Sub_15_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U17 ( .A(r[122]), .B(
        Midori_rounds_sub_Sub_15_F_q3[3]), .ZN(Midori_rounds_sub_Sub_15_F_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U16 ( .A(Midori_rounds_sub_Sub_15_F_n11), 
        .B(r[121]), .ZN(Midori_rounds_sub_Sub_15_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U15 ( .A(r[120]), .B(
        Midori_rounds_sub_Sub_15_F_q3[2]), .ZN(Midori_rounds_sub_Sub_15_F_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U14 ( .A(Midori_rounds_sub_Sub_15_F_n10), 
        .B(r[127]), .ZN(Midori_rounds_sub_Sub_15_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U13 ( .A(r[126]), .B(
        Midori_rounds_sub_Sub_15_F_q3[1]), .ZN(Midori_rounds_sub_Sub_15_F_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U12 ( .A(Midori_rounds_sub_Sub_15_F_n9), 
        .B(r[125]), .ZN(Midori_rounds_sub_Sub_15_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_U11 ( .A(r[124]), .B(
        Midori_rounds_sub_Sub_15_F_q3[0]), .ZN(Midori_rounds_sub_Sub_15_F_n9)
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U10 ( .A(r[123]), .B(
        Midori_rounds_sub_Sub_15_F_q2[3]), .Z(Midori_rounds_sub_Sub_15_q2[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U9 ( .A(r[121]), .B(
        Midori_rounds_sub_Sub_15_F_q2[2]), .Z(Midori_rounds_sub_Sub_15_q2[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U8 ( .A(r[127]), .B(
        Midori_rounds_sub_Sub_15_F_q2[1]), .Z(Midori_rounds_sub_Sub_15_q2[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U7 ( .A(r[125]), .B(
        Midori_rounds_sub_Sub_15_F_q2[0]), .Z(Midori_rounds_sub_Sub_15_q2[0])
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U6 ( .A(r[122]), .B(
        Midori_rounds_sub_Sub_15_F_q1[3]), .Z(Midori_rounds_sub_Sub_15_q1[3])
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U5 ( .A(r[120]), .B(
        Midori_rounds_sub_Sub_15_F_q1[2]), .Z(Midori_rounds_sub_Sub_15_q1[2])
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U4 ( .A(r[126]), .B(
        Midori_rounds_sub_Sub_15_F_q1[1]), .Z(Midori_rounds_sub_Sub_15_q1[1])
         );
  XOR2_X1 Midori_rounds_sub_Sub_15_F_U3 ( .A(r[124]), .B(
        Midori_rounds_sub_Sub_15_F_q1[0]), .Z(Midori_rounds_sub_Sub_15_q1[0])
         );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[26]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_27_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[27]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[27]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_28_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[28]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[28]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_29_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[29]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_30_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[30]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[30]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_31_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[31]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[31]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_32_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[32]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[32]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_33_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[33]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_34_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[34]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[34]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_F_CF_Reg_reg_35_ ( .D(
        Midori_rounds_sub_Sub_15_F_CF_Out[35]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_F_CF_Reg[35]), .QN() );
  AND2_X1 Midori_rounds_sub_Sub_15_F_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_Inst_1__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[1]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_F_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_1__CF_Inst_n3) );
  OR2_X1 Midori_rounds_sub_Sub_15_F_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_F_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_3__CF_Inst_n3) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_4__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_4__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[4]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_4__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_4__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_5__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_5__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[5]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_5__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_5__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_8__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_9__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_9__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[9]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_9__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_9__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[10]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_10__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_11__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_11__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[11]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_11__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_11__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_n6) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_12__CF_Inst_n5) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_13__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[13]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_13__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_14__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_15__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_15__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[15]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_15__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_15__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_Inst_17__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[17]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_17__CF_Inst_n6) );
  AOI211_X1 Midori_rounds_sub_Sub_15_F_Inst_18__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_18__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[18]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_18__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_19__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_20__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_15_F_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .B(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .S(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .Z(
        Midori_rounds_sub_Sub_15_F_CF_Out[21]) );
  AOI21_X1 Midori_rounds_sub_Sub_15_F_Inst_22__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_Inst_22__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[22]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_22__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_22__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_15_F_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_15_F_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .C2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_24__CF_Inst_n3) );
  MUX2_X1 Midori_rounds_sub_Sub_15_F_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_15_F_CF_Out[25]) );
  AOI21_X1 Midori_rounds_sub_Sub_15_F_Inst_26__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_Inst_26__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[26]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_26__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_26__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[0]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[27]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_n8), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_27__CF_Inst_n8) );
  AOI21_X1 Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[28]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_28__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A(
        Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[29]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_29__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[0]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[30]) );
  AOI22_X1 Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .A2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .B1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_30__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_15_F_Inst_31__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_Inst_31__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[31]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_31__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_31__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_15_F_Inst_32__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .C2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[3]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_32__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[32]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_32__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .A2(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_32__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[0]), .B(
        Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[33]) );
  AOI221_X1 Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n10), .C1(
        Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n9), .C2(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n11) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in1_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_33__CF_Inst_n10) );
  MUX2_X1 Midori_rounds_sub_Sub_15_F_Inst_34__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in2_reg[1]), .B(
        Midori_rounds_sub_Sub_15_F_in2_reg[2]), .S(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .Z(
        Midori_rounds_sub_Sub_15_F_CF_Out[34]) );
  AOI21_X1 Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_F_CF_Out[35]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_F_in3_reg[1]), .B2(
        Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_in3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_Inst_35__CF_Inst_n4) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_15_F_q1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_15_F_q2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_15_F_q3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_15_F_q1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_15_F_q2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_15_F_q3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_15_F_q1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_15_F_q2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_15_F_q3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression1_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[29]), .ZN(
        Midori_rounds_sub_Sub_15_F_q1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[27]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[28]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression2_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[32]), .ZN(
        Midori_rounds_sub_Sub_15_F_q2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[30]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[31]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression3_n3), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[35]), .ZN(
        Midori_rounds_sub_Sub_15_F_q3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_15_F_CF_Reg[33]), .B(
        Midori_rounds_sub_Sub_15_F_CF_Reg[34]), .ZN(
        Midori_rounds_sub_Sub_15_F_InstXOR_3__Compression3_n3) );
  INV_X1 Midori_rounds_sub_Sub_15_G_U3 ( .A(Midori_rounds_sub_Sub_15_Rq1[0]), 
        .ZN(Midori_rounds_sub_Sub_15_G_n1) );
  DFF_X1 Midori_rounds_sub_Sub_15_G_out3_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_Rq3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[61]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_out2_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_Rq2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[61]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_out1_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_G_n1), .CK(clk), .Q(
        Midori_rounds_SR_Result1[61]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_15_G_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_15_G_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_15_G_CF_Reg[26]), .QN() );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_0__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[3]), .A2(
        Midori_rounds_sub_Sub_15_G_Inst_0__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[0]) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_0__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq1[1]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_0__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_1__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_Inst_1__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_15_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[1]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .A2(Midori_rounds_sub_Sub_15_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_1__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_15_G_Inst_2__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[3]), .A2(Midori_rounds_sub_Sub_15_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_15_G_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_Inst_3__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_15_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .A2(Midori_rounds_sub_Sub_15_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_3__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_15_G_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .A2(Midori_rounds_sub_Sub_15_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_CF_Out[4]) );
  OR2_X1 Midori_rounds_sub_Sub_15_G_Inst_5__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq2[3]), .A2(Midori_rounds_sub_Sub_15_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_15_G_CF_Out[5]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_6__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .A2(
        Midori_rounds_sub_Sub_15_G_Inst_6__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[6]) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_6__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_6__CF_Inst_n2) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_15_G_Inst_7__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[7]) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_7__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_7__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_Inst_8__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_15_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_8__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq3[1]), .A2(Midori_rounds_sub_Sub_15_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_8__CF_Inst_n3) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .A2(Midori_rounds_sub_Sub_15_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_CF_Out[9]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_Inst_10__CF_Inst_n6), .B(
        Midori_rounds_sub_Sub_15_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[10]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_10__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .A2(Midori_rounds_sub_Sub_15_Rq1[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_10__CF_Inst_n6) );
  OR2_X1 Midori_rounds_sub_Sub_15_G_Inst_11__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[3]), .A2(Midori_rounds_sub_Sub_15_Rq3[1]), 
        .ZN(Midori_rounds_sub_Sub_15_G_CF_Out[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_Inst_12__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_15_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .A2(Midori_rounds_sub_Sub_15_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_12__CF_Inst_n3) );
  AND2_X1 Midori_rounds_sub_Sub_15_G_Inst_13__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .A2(Midori_rounds_sub_Sub_15_Rq2[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_CF_Out[13]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_14__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_Rq2[3]), .A2(
        Midori_rounds_sub_Sub_15_G_Inst_14__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[14]) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_14__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_14__CF_Inst_n2) );
  AND2_X1 Midori_rounds_sub_Sub_15_G_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .A2(Midori_rounds_sub_Sub_15_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_CF_Out[15]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_16__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_Rq3[3]), .A2(
        Midori_rounds_sub_Sub_15_G_Inst_16__CF_Inst_n2), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[16]) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_16__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_16__CF_Inst_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_17__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_Inst_17__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_15_Rq3[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[17]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_17__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq3[1]), .A2(Midori_rounds_sub_Sub_15_Rq3[3]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_17__CF_Inst_n3) );
  OAI21_X1 Midori_rounds_sub_Sub_15_G_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_Rq1[3]), .B2(Midori_rounds_sub_Sub_15_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_15_G_Inst_18__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[3]), .A2(Midori_rounds_sub_Sub_15_Rq1[1]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_18__CF_Inst_n9) );
  AOI21_X1 Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[19]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_Rq1[3]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_19__CF_Inst_n4) );
  AOI211_X1 Midori_rounds_sub_Sub_15_G_Inst_20__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_15_Rq3[1]), .C2(Midori_rounds_sub_Sub_15_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_15_Rq1[3]), .B(
        Midori_rounds_sub_Sub_15_G_Inst_20__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[20]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_20__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq3[1]), .A2(Midori_rounds_sub_Sub_15_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_20__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[21]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .B2(
        Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq1[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_21__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_15_Rq2[2]), .A(
        Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[22]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_15_Rq2[1]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq2[3]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_22__CF_Inst_n10) );
  AOI211_X1 Midori_rounds_sub_Sub_15_G_Inst_23__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_15_Rq3[1]), .C2(Midori_rounds_sub_Sub_15_Rq3[2]), 
        .A(Midori_rounds_sub_Sub_15_Rq2[3]), .B(
        Midori_rounds_sub_Sub_15_G_Inst_23__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[23]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_23__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq3[1]), .A2(Midori_rounds_sub_Sub_15_Rq3[2]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_23__CF_Inst_n3) );
  AOI211_X1 Midori_rounds_sub_Sub_15_G_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .C2(Midori_rounds_sub_Sub_15_Rq1[2]), 
        .A(Midori_rounds_sub_Sub_15_Rq3[3]), .B(
        Midori_rounds_sub_Sub_15_G_Inst_24__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[24]) );
  NOR2_X1 Midori_rounds_sub_Sub_15_G_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_15_Rq1[1]), .A2(Midori_rounds_sub_Sub_15_Rq1[2]), 
        .ZN(Midori_rounds_sub_Sub_15_G_Inst_24__CF_Inst_n3) );
  AOI21_X1 Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_n3), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[25]) );
  OAI21_X1 Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_15_Rq2[1]), .B2(
        Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_n4), .A(
        Midori_rounds_sub_Sub_15_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_n3) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq2[2]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_25__CF_Inst_n4) );
  OAI21_X1 Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_U3 ( .B1(
        Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_n10), .B2(
        Midori_rounds_sub_Sub_15_Rq3[2]), .A(
        Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_15_G_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_n10), .A2(
        Midori_rounds_sub_Sub_15_Rq3[1]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_n9) );
  INV_X1 Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_15_Rq3[3]), .ZN(
        Midori_rounds_sub_Sub_15_G_Inst_26__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[60]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[60]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[60]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[62]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[62]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[62]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR2_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[63]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[63]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[63]) );
  XNOR2_X1 Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_15_G_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_15_G_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_15_G_InstXOR2_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U24 ( .A(Midori_rounds_mul_input1[61]), .B(
        Midori_rounds_mul1_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result1[21]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U23 ( .A(Midori_rounds_mul_input1[60]), .B(
        Midori_rounds_mul1_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result1[20]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U22 ( .A(Midori_rounds_mul_input1[51]), .B(
        Midori_rounds_mul1_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result1[43]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U21 ( .A(Midori_rounds_mul_input1[50]), .B(
        Midori_rounds_mul1_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result1[42]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U20 ( .A(Midori_rounds_mul_input1[49]), .B(
        Midori_rounds_mul1_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result1[41]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U19 ( .A(Midori_rounds_mul_input1[48]), .B(
        Midori_rounds_mul1_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result1[40]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U18 ( .A(Midori_rounds_mul_input1[55]), .B(
        Midori_rounds_mul1_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result1[3]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U17 ( .A(Midori_rounds_mul_input1[63]), .B(
        Midori_rounds_mul_input1[59]), .ZN(Midori_rounds_mul1_MC1_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U16 ( .A(Midori_rounds_mul_input1[54]), .B(
        Midori_rounds_mul1_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result1[2]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U15 ( .A(Midori_rounds_mul_input1[62]), .B(
        Midori_rounds_mul_input1[58]), .ZN(Midori_rounds_mul1_MC1_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U14 ( .A(Midori_rounds_mul_input1[53]), .B(
        Midori_rounds_mul1_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result1[1]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U13 ( .A(Midori_rounds_mul_input1[57]), .B(
        Midori_rounds_mul_input1[61]), .ZN(Midori_rounds_mul1_MC1_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U12 ( .A(Midori_rounds_mul_input1[59]), .B(
        Midori_rounds_mul1_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result1[63]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U11 ( .A(Midori_rounds_mul_input1[58]), .B(
        Midori_rounds_mul1_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result1[62]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U10 ( .A(Midori_rounds_mul_input1[57]), .B(
        Midori_rounds_mul1_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result1[61]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U9 ( .A(Midori_rounds_mul_input1[49]), .B(
        Midori_rounds_mul_input1[53]), .ZN(Midori_rounds_mul1_MC1_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U8 ( .A(Midori_rounds_mul_input1[56]), .B(
        Midori_rounds_mul1_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result1[60]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U7 ( .A(Midori_rounds_mul_input1[52]), .B(
        Midori_rounds_mul_input1[48]), .ZN(Midori_rounds_mul1_MC1_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U6 ( .A(Midori_rounds_mul_input1[63]), .B(
        Midori_rounds_mul1_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result1[23]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U5 ( .A(Midori_rounds_mul_input1[51]), .B(
        Midori_rounds_mul_input1[55]), .ZN(Midori_rounds_mul1_MC1_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U4 ( .A(Midori_rounds_mul_input1[62]), .B(
        Midori_rounds_mul1_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result1[22]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U3 ( .A(Midori_rounds_mul_input1[50]), .B(
        Midori_rounds_mul_input1[54]), .ZN(Midori_rounds_mul1_MC1_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U2 ( .A(Midori_rounds_mul_input1[52]), .B(
        Midori_rounds_mul1_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result1[0]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U1 ( .A(Midori_rounds_mul_input1[60]), .B(
        Midori_rounds_mul_input1[56]), .ZN(Midori_rounds_mul1_MC1_n19) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U24 ( .A(Midori_rounds_mul_input1[45]), .B(
        Midori_rounds_mul1_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result1[45]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U23 ( .A(Midori_rounds_mul_input1[44]), .B(
        Midori_rounds_mul1_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result1[44]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U22 ( .A(Midori_rounds_mul_input1[35]), .B(
        Midori_rounds_mul1_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result1[19]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U21 ( .A(Midori_rounds_mul_input1[34]), .B(
        Midori_rounds_mul1_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result1[18]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U20 ( .A(Midori_rounds_mul_input1[33]), .B(
        Midori_rounds_mul1_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result1[17]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U19 ( .A(Midori_rounds_mul_input1[32]), .B(
        Midori_rounds_mul1_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result1[16]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U18 ( .A(Midori_rounds_mul_input1[39]), .B(
        Midori_rounds_mul1_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result1[59]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U17 ( .A(Midori_rounds_mul_input1[47]), .B(
        Midori_rounds_mul_input1[43]), .ZN(Midori_rounds_mul1_MC2_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U16 ( .A(Midori_rounds_mul_input1[38]), .B(
        Midori_rounds_mul1_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result1[58]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U15 ( .A(Midori_rounds_mul_input1[46]), .B(
        Midori_rounds_mul_input1[42]), .ZN(Midori_rounds_mul1_MC2_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U14 ( .A(Midori_rounds_mul_input1[37]), .B(
        Midori_rounds_mul1_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result1[57]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U13 ( .A(Midori_rounds_mul_input1[41]), .B(
        Midori_rounds_mul_input1[45]), .ZN(Midori_rounds_mul1_MC2_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U12 ( .A(Midori_rounds_mul_input1[43]), .B(
        Midori_rounds_mul1_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result1[7]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U11 ( .A(Midori_rounds_mul_input1[42]), .B(
        Midori_rounds_mul1_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result1[6]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U10 ( .A(Midori_rounds_mul_input1[41]), .B(
        Midori_rounds_mul1_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result1[5]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U9 ( .A(Midori_rounds_mul_input1[33]), .B(
        Midori_rounds_mul_input1[37]), .ZN(Midori_rounds_mul1_MC2_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U8 ( .A(Midori_rounds_mul_input1[40]), .B(
        Midori_rounds_mul1_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result1[4]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U7 ( .A(Midori_rounds_mul_input1[36]), .B(
        Midori_rounds_mul_input1[32]), .ZN(Midori_rounds_mul1_MC2_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U6 ( .A(Midori_rounds_mul_input1[47]), .B(
        Midori_rounds_mul1_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result1[47]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U5 ( .A(Midori_rounds_mul_input1[35]), .B(
        Midori_rounds_mul_input1[39]), .ZN(Midori_rounds_mul1_MC2_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U4 ( .A(Midori_rounds_mul_input1[46]), .B(
        Midori_rounds_mul1_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result1[46]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U3 ( .A(Midori_rounds_mul_input1[34]), .B(
        Midori_rounds_mul_input1[38]), .ZN(Midori_rounds_mul1_MC2_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U2 ( .A(Midori_rounds_mul_input1[36]), .B(
        Midori_rounds_mul1_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result1[56]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U1 ( .A(Midori_rounds_mul_input1[44]), .B(
        Midori_rounds_mul_input1[40]), .ZN(Midori_rounds_mul1_MC2_n19) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U24 ( .A(Midori_rounds_mul_input1[29]), .B(
        Midori_rounds_mul1_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result1[49]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U23 ( .A(Midori_rounds_mul_input1[28]), .B(
        Midori_rounds_mul1_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result1[48]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U22 ( .A(Midori_rounds_mul_input1[19]), .B(
        Midori_rounds_mul1_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result1[15]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U21 ( .A(Midori_rounds_mul_input1[18]), .B(
        Midori_rounds_mul1_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result1[14]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U20 ( .A(Midori_rounds_mul_input1[17]), .B(
        Midori_rounds_mul1_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result1[13]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U19 ( .A(Midori_rounds_mul_input1[16]), .B(
        Midori_rounds_mul1_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result1[12]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U18 ( .A(Midori_rounds_mul_input1[23]), .B(
        Midori_rounds_mul1_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result1[39]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U17 ( .A(Midori_rounds_mul_input1[31]), .B(
        Midori_rounds_mul_input1[27]), .ZN(Midori_rounds_mul1_MC3_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U16 ( .A(Midori_rounds_mul_input1[22]), .B(
        Midori_rounds_mul1_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result1[38]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U15 ( .A(Midori_rounds_mul_input1[30]), .B(
        Midori_rounds_mul_input1[26]), .ZN(Midori_rounds_mul1_MC3_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U14 ( .A(Midori_rounds_mul_input1[21]), .B(
        Midori_rounds_mul1_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result1[37]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U13 ( .A(Midori_rounds_mul_input1[25]), .B(
        Midori_rounds_mul_input1[29]), .ZN(Midori_rounds_mul1_MC3_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U12 ( .A(Midori_rounds_mul_input1[27]), .B(
        Midori_rounds_mul1_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result1[27]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U11 ( .A(Midori_rounds_mul_input1[26]), .B(
        Midori_rounds_mul1_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result1[26]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U10 ( .A(Midori_rounds_mul_input1[25]), .B(
        Midori_rounds_mul1_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result1[25]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U9 ( .A(Midori_rounds_mul_input1[17]), .B(
        Midori_rounds_mul_input1[21]), .ZN(Midori_rounds_mul1_MC3_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U8 ( .A(Midori_rounds_mul_input1[24]), .B(
        Midori_rounds_mul1_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result1[24]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U7 ( .A(Midori_rounds_mul_input1[20]), .B(
        Midori_rounds_mul_input1[16]), .ZN(Midori_rounds_mul1_MC3_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U6 ( .A(Midori_rounds_mul_input1[31]), .B(
        Midori_rounds_mul1_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result1[51]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U5 ( .A(Midori_rounds_mul_input1[19]), .B(
        Midori_rounds_mul_input1[23]), .ZN(Midori_rounds_mul1_MC3_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U4 ( .A(Midori_rounds_mul_input1[30]), .B(
        Midori_rounds_mul1_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result1[50]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U3 ( .A(Midori_rounds_mul_input1[18]), .B(
        Midori_rounds_mul_input1[22]), .ZN(Midori_rounds_mul1_MC3_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U2 ( .A(Midori_rounds_mul_input1[20]), .B(
        Midori_rounds_mul1_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result1[36]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U1 ( .A(Midori_rounds_mul_input1[28]), .B(
        Midori_rounds_mul_input1[24]), .ZN(Midori_rounds_mul1_MC3_n19) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U24 ( .A(Midori_rounds_mul_input1[13]), .B(
        Midori_rounds_mul1_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result1[9]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U23 ( .A(Midori_rounds_mul_input1[12]), .B(
        Midori_rounds_mul1_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result1[8]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U22 ( .A(Midori_rounds_mul_input1[3]), .B(
        Midori_rounds_mul1_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result1[55]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U21 ( .A(Midori_rounds_mul_input1[2]), .B(
        Midori_rounds_mul1_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result1[54]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U20 ( .A(Midori_rounds_mul_input1[1]), .B(
        Midori_rounds_mul1_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result1[53]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U19 ( .A(Midori_rounds_mul_input1[0]), .B(
        Midori_rounds_mul1_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result1[52]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U18 ( .A(Midori_rounds_mul_input1[7]), .B(
        Midori_rounds_mul1_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result1[31]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U17 ( .A(Midori_rounds_mul_input1[15]), .B(
        Midori_rounds_mul_input1[11]), .ZN(Midori_rounds_mul1_MC4_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U16 ( .A(Midori_rounds_mul_input1[6]), .B(
        Midori_rounds_mul1_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result1[30]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U15 ( .A(Midori_rounds_mul_input1[14]), .B(
        Midori_rounds_mul_input1[10]), .ZN(Midori_rounds_mul1_MC4_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U14 ( .A(Midori_rounds_mul_input1[5]), .B(
        Midori_rounds_mul1_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result1[29]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U13 ( .A(Midori_rounds_mul_input1[9]), .B(
        Midori_rounds_mul_input1[13]), .ZN(Midori_rounds_mul1_MC4_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U12 ( .A(Midori_rounds_mul_input1[11]), .B(
        Midori_rounds_mul1_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result1[35]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U11 ( .A(Midori_rounds_mul_input1[10]), .B(
        Midori_rounds_mul1_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result1[34]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U10 ( .A(Midori_rounds_mul_input1[9]), .B(
        Midori_rounds_mul1_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result1[33]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U9 ( .A(Midori_rounds_mul_input1[1]), .B(
        Midori_rounds_mul_input1[5]), .ZN(Midori_rounds_mul1_MC4_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U8 ( .A(Midori_rounds_mul_input1[8]), .B(
        Midori_rounds_mul1_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result1[32]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U7 ( .A(Midori_rounds_mul_input1[4]), .B(
        Midori_rounds_mul_input1[0]), .ZN(Midori_rounds_mul1_MC4_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U6 ( .A(Midori_rounds_mul_input1[15]), .B(
        Midori_rounds_mul1_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result1[11]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U5 ( .A(Midori_rounds_mul_input1[3]), .B(
        Midori_rounds_mul_input1[7]), .ZN(Midori_rounds_mul1_MC4_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U4 ( .A(Midori_rounds_mul_input1[14]), .B(
        Midori_rounds_mul1_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result1[10]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U3 ( .A(Midori_rounds_mul_input1[2]), .B(
        Midori_rounds_mul_input1[6]), .ZN(Midori_rounds_mul1_MC4_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U2 ( .A(Midori_rounds_mul_input1[4]), .B(
        Midori_rounds_mul1_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result1[28]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U1 ( .A(Midori_rounds_mul_input1[12]), .B(
        Midori_rounds_mul_input1[8]), .ZN(Midori_rounds_mul1_MC4_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U24 ( .A(Midori_rounds_mul_input2[61]), .B(
        Midori_rounds_mul2_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result2[21]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U23 ( .A(Midori_rounds_mul_input2[60]), .B(
        Midori_rounds_mul2_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result2[20]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U22 ( .A(Midori_rounds_mul_input2[51]), .B(
        Midori_rounds_mul2_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result2[43]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U21 ( .A(Midori_rounds_mul_input2[50]), .B(
        Midori_rounds_mul2_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result2[42]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U20 ( .A(Midori_rounds_mul_input2[49]), .B(
        Midori_rounds_mul2_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result2[41]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U19 ( .A(Midori_rounds_mul_input2[48]), .B(
        Midori_rounds_mul2_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result2[40]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U18 ( .A(Midori_rounds_mul_input2[55]), .B(
        Midori_rounds_mul2_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result2[3]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U17 ( .A(Midori_rounds_mul_input2[63]), .B(
        Midori_rounds_mul_input2[59]), .ZN(Midori_rounds_mul2_MC1_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U16 ( .A(Midori_rounds_mul_input2[54]), .B(
        Midori_rounds_mul2_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result2[2]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U15 ( .A(Midori_rounds_mul_input2[62]), .B(
        Midori_rounds_mul_input2[58]), .ZN(Midori_rounds_mul2_MC1_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U14 ( .A(Midori_rounds_mul_input2[53]), .B(
        Midori_rounds_mul2_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result2[1]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U13 ( .A(Midori_rounds_mul_input2[57]), .B(
        Midori_rounds_mul_input2[61]), .ZN(Midori_rounds_mul2_MC1_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U12 ( .A(Midori_rounds_mul_input2[59]), .B(
        Midori_rounds_mul2_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result2[63]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U11 ( .A(Midori_rounds_mul_input2[58]), .B(
        Midori_rounds_mul2_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result2[62]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U10 ( .A(Midori_rounds_mul_input2[57]), .B(
        Midori_rounds_mul2_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result2[61]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U9 ( .A(Midori_rounds_mul_input2[49]), .B(
        Midori_rounds_mul_input2[53]), .ZN(Midori_rounds_mul2_MC1_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U8 ( .A(Midori_rounds_mul_input2[56]), .B(
        Midori_rounds_mul2_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result2[60]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U7 ( .A(Midori_rounds_mul_input2[52]), .B(
        Midori_rounds_mul_input2[48]), .ZN(Midori_rounds_mul2_MC1_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U6 ( .A(Midori_rounds_mul_input2[63]), .B(
        Midori_rounds_mul2_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result2[23]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U5 ( .A(Midori_rounds_mul_input2[51]), .B(
        Midori_rounds_mul_input2[55]), .ZN(Midori_rounds_mul2_MC1_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U4 ( .A(Midori_rounds_mul_input2[62]), .B(
        Midori_rounds_mul2_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result2[22]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U3 ( .A(Midori_rounds_mul_input2[50]), .B(
        Midori_rounds_mul_input2[54]), .ZN(Midori_rounds_mul2_MC1_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U2 ( .A(Midori_rounds_mul_input2[52]), .B(
        Midori_rounds_mul2_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result2[0]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U1 ( .A(Midori_rounds_mul_input2[60]), .B(
        Midori_rounds_mul_input2[56]), .ZN(Midori_rounds_mul2_MC1_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U24 ( .A(Midori_rounds_mul_input2[45]), .B(
        Midori_rounds_mul2_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result2[45]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U23 ( .A(Midori_rounds_mul_input2[44]), .B(
        Midori_rounds_mul2_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result2[44]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U22 ( .A(Midori_rounds_mul_input2[35]), .B(
        Midori_rounds_mul2_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result2[19]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U21 ( .A(Midori_rounds_mul_input2[34]), .B(
        Midori_rounds_mul2_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result2[18]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U20 ( .A(Midori_rounds_mul_input2[33]), .B(
        Midori_rounds_mul2_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result2[17]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U19 ( .A(Midori_rounds_mul_input2[32]), .B(
        Midori_rounds_mul2_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result2[16]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U18 ( .A(Midori_rounds_mul_input2[39]), .B(
        Midori_rounds_mul2_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result2[59]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U17 ( .A(Midori_rounds_mul_input2[47]), .B(
        Midori_rounds_mul_input2[43]), .ZN(Midori_rounds_mul2_MC2_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U16 ( .A(Midori_rounds_mul_input2[38]), .B(
        Midori_rounds_mul2_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result2[58]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U15 ( .A(Midori_rounds_mul_input2[46]), .B(
        Midori_rounds_mul_input2[42]), .ZN(Midori_rounds_mul2_MC2_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U14 ( .A(Midori_rounds_mul_input2[37]), .B(
        Midori_rounds_mul2_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result2[57]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U13 ( .A(Midori_rounds_mul_input2[41]), .B(
        Midori_rounds_mul_input2[45]), .ZN(Midori_rounds_mul2_MC2_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U12 ( .A(Midori_rounds_mul_input2[43]), .B(
        Midori_rounds_mul2_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result2[7]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U11 ( .A(Midori_rounds_mul_input2[42]), .B(
        Midori_rounds_mul2_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result2[6]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U10 ( .A(Midori_rounds_mul_input2[41]), .B(
        Midori_rounds_mul2_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result2[5]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U9 ( .A(Midori_rounds_mul_input2[33]), .B(
        Midori_rounds_mul_input2[37]), .ZN(Midori_rounds_mul2_MC2_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U8 ( .A(Midori_rounds_mul_input2[40]), .B(
        Midori_rounds_mul2_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result2[4]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U7 ( .A(Midori_rounds_mul_input2[36]), .B(
        Midori_rounds_mul_input2[32]), .ZN(Midori_rounds_mul2_MC2_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U6 ( .A(Midori_rounds_mul_input2[47]), .B(
        Midori_rounds_mul2_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result2[47]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U5 ( .A(Midori_rounds_mul_input2[35]), .B(
        Midori_rounds_mul_input2[39]), .ZN(Midori_rounds_mul2_MC2_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U4 ( .A(Midori_rounds_mul_input2[46]), .B(
        Midori_rounds_mul2_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result2[46]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U3 ( .A(Midori_rounds_mul_input2[34]), .B(
        Midori_rounds_mul_input2[38]), .ZN(Midori_rounds_mul2_MC2_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U2 ( .A(Midori_rounds_mul_input2[36]), .B(
        Midori_rounds_mul2_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result2[56]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U1 ( .A(Midori_rounds_mul_input2[44]), .B(
        Midori_rounds_mul_input2[40]), .ZN(Midori_rounds_mul2_MC2_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U24 ( .A(Midori_rounds_mul_input2[29]), .B(
        Midori_rounds_mul2_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result2[49]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U23 ( .A(Midori_rounds_mul_input2[28]), .B(
        Midori_rounds_mul2_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result2[48]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U22 ( .A(Midori_rounds_mul_input2[19]), .B(
        Midori_rounds_mul2_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result2[15]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U21 ( .A(Midori_rounds_mul_input2[18]), .B(
        Midori_rounds_mul2_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result2[14]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U20 ( .A(Midori_rounds_mul_input2[17]), .B(
        Midori_rounds_mul2_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result2[13]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U19 ( .A(Midori_rounds_mul_input2[16]), .B(
        Midori_rounds_mul2_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result2[12]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U18 ( .A(Midori_rounds_mul_input2[23]), .B(
        Midori_rounds_mul2_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result2[39]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U17 ( .A(Midori_rounds_mul_input2[31]), .B(
        Midori_rounds_mul_input2[27]), .ZN(Midori_rounds_mul2_MC3_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U16 ( .A(Midori_rounds_mul_input2[22]), .B(
        Midori_rounds_mul2_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result2[38]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U15 ( .A(Midori_rounds_mul_input2[30]), .B(
        Midori_rounds_mul_input2[26]), .ZN(Midori_rounds_mul2_MC3_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U14 ( .A(Midori_rounds_mul_input2[21]), .B(
        Midori_rounds_mul2_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result2[37]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U13 ( .A(Midori_rounds_mul_input2[25]), .B(
        Midori_rounds_mul_input2[29]), .ZN(Midori_rounds_mul2_MC3_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U12 ( .A(Midori_rounds_mul_input2[27]), .B(
        Midori_rounds_mul2_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result2[27]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U11 ( .A(Midori_rounds_mul_input2[26]), .B(
        Midori_rounds_mul2_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result2[26]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U10 ( .A(Midori_rounds_mul_input2[25]), .B(
        Midori_rounds_mul2_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result2[25]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U9 ( .A(Midori_rounds_mul_input2[17]), .B(
        Midori_rounds_mul_input2[21]), .ZN(Midori_rounds_mul2_MC3_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U8 ( .A(Midori_rounds_mul_input2[24]), .B(
        Midori_rounds_mul2_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result2[24]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U7 ( .A(Midori_rounds_mul_input2[20]), .B(
        Midori_rounds_mul_input2[16]), .ZN(Midori_rounds_mul2_MC3_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U6 ( .A(Midori_rounds_mul_input2[31]), .B(
        Midori_rounds_mul2_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result2[51]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U5 ( .A(Midori_rounds_mul_input2[19]), .B(
        Midori_rounds_mul_input2[23]), .ZN(Midori_rounds_mul2_MC3_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U4 ( .A(Midori_rounds_mul_input2[30]), .B(
        Midori_rounds_mul2_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result2[50]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U3 ( .A(Midori_rounds_mul_input2[18]), .B(
        Midori_rounds_mul_input2[22]), .ZN(Midori_rounds_mul2_MC3_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U2 ( .A(Midori_rounds_mul_input2[20]), .B(
        Midori_rounds_mul2_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result2[36]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U1 ( .A(Midori_rounds_mul_input2[28]), .B(
        Midori_rounds_mul_input2[24]), .ZN(Midori_rounds_mul2_MC3_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U24 ( .A(Midori_rounds_mul_input2[13]), .B(
        Midori_rounds_mul2_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result2[9]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U23 ( .A(Midori_rounds_mul_input2[12]), .B(
        Midori_rounds_mul2_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result2[8]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U22 ( .A(Midori_rounds_mul_input2[3]), .B(
        Midori_rounds_mul2_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result2[55]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U21 ( .A(Midori_rounds_mul_input2[2]), .B(
        Midori_rounds_mul2_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result2[54]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U20 ( .A(Midori_rounds_mul_input2[1]), .B(
        Midori_rounds_mul2_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result2[53]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U19 ( .A(Midori_rounds_mul_input2[0]), .B(
        Midori_rounds_mul2_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result2[52]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U18 ( .A(Midori_rounds_mul_input2[7]), .B(
        Midori_rounds_mul2_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result2[31]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U17 ( .A(Midori_rounds_mul_input2[15]), .B(
        Midori_rounds_mul_input2[11]), .ZN(Midori_rounds_mul2_MC4_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U16 ( .A(Midori_rounds_mul_input2[6]), .B(
        Midori_rounds_mul2_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result2[30]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U15 ( .A(Midori_rounds_mul_input2[14]), .B(
        Midori_rounds_mul_input2[10]), .ZN(Midori_rounds_mul2_MC4_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U14 ( .A(Midori_rounds_mul_input2[5]), .B(
        Midori_rounds_mul2_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result2[29]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U13 ( .A(Midori_rounds_mul_input2[9]), .B(
        Midori_rounds_mul_input2[13]), .ZN(Midori_rounds_mul2_MC4_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U12 ( .A(Midori_rounds_mul_input2[11]), .B(
        Midori_rounds_mul2_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result2[35]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U11 ( .A(Midori_rounds_mul_input2[10]), .B(
        Midori_rounds_mul2_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result2[34]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U10 ( .A(Midori_rounds_mul_input2[9]), .B(
        Midori_rounds_mul2_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result2[33]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U9 ( .A(Midori_rounds_mul_input2[1]), .B(
        Midori_rounds_mul_input2[5]), .ZN(Midori_rounds_mul2_MC4_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U8 ( .A(Midori_rounds_mul_input2[8]), .B(
        Midori_rounds_mul2_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result2[32]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U7 ( .A(Midori_rounds_mul_input2[4]), .B(
        Midori_rounds_mul_input2[0]), .ZN(Midori_rounds_mul2_MC4_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U6 ( .A(Midori_rounds_mul_input2[15]), .B(
        Midori_rounds_mul2_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result2[11]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U5 ( .A(Midori_rounds_mul_input2[3]), .B(
        Midori_rounds_mul_input2[7]), .ZN(Midori_rounds_mul2_MC4_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U4 ( .A(Midori_rounds_mul_input2[14]), .B(
        Midori_rounds_mul2_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result2[10]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U3 ( .A(Midori_rounds_mul_input2[2]), .B(
        Midori_rounds_mul_input2[6]), .ZN(Midori_rounds_mul2_MC4_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U2 ( .A(Midori_rounds_mul_input2[4]), .B(
        Midori_rounds_mul2_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result2[28]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U1 ( .A(Midori_rounds_mul_input2[12]), .B(
        Midori_rounds_mul_input2[8]), .ZN(Midori_rounds_mul2_MC4_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U24 ( .A(Midori_rounds_mul_input3[61]), .B(
        Midori_rounds_mul3_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result3[21]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U23 ( .A(Midori_rounds_mul_input3[60]), .B(
        Midori_rounds_mul3_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result3[20]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U22 ( .A(Midori_rounds_mul_input3[51]), .B(
        Midori_rounds_mul3_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result3[43]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U21 ( .A(Midori_rounds_mul_input3[50]), .B(
        Midori_rounds_mul3_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result3[42]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U20 ( .A(Midori_rounds_mul_input3[49]), .B(
        Midori_rounds_mul3_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result3[41]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U19 ( .A(Midori_rounds_mul_input3[48]), .B(
        Midori_rounds_mul3_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result3[40]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U18 ( .A(Midori_rounds_mul_input3[55]), .B(
        Midori_rounds_mul3_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result3[3]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U17 ( .A(Midori_rounds_mul_input3[63]), .B(
        Midori_rounds_mul_input3[59]), .ZN(Midori_rounds_mul3_MC1_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U16 ( .A(Midori_rounds_mul_input3[54]), .B(
        Midori_rounds_mul3_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result3[2]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U15 ( .A(Midori_rounds_mul_input3[62]), .B(
        Midori_rounds_mul_input3[58]), .ZN(Midori_rounds_mul3_MC1_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U14 ( .A(Midori_rounds_mul_input3[53]), .B(
        Midori_rounds_mul3_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result3[1]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U13 ( .A(Midori_rounds_mul_input3[57]), .B(
        Midori_rounds_mul_input3[61]), .ZN(Midori_rounds_mul3_MC1_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U12 ( .A(Midori_rounds_mul_input3[59]), .B(
        Midori_rounds_mul3_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result3[63]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U11 ( .A(Midori_rounds_mul_input3[58]), .B(
        Midori_rounds_mul3_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result3[62]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U10 ( .A(Midori_rounds_mul_input3[57]), .B(
        Midori_rounds_mul3_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result3[61]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U9 ( .A(Midori_rounds_mul_input3[49]), .B(
        Midori_rounds_mul_input3[53]), .ZN(Midori_rounds_mul3_MC1_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U8 ( .A(Midori_rounds_mul_input3[56]), .B(
        Midori_rounds_mul3_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result3[60]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U7 ( .A(Midori_rounds_mul_input3[52]), .B(
        Midori_rounds_mul_input3[48]), .ZN(Midori_rounds_mul3_MC1_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U6 ( .A(Midori_rounds_mul_input3[63]), .B(
        Midori_rounds_mul3_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result3[23]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U5 ( .A(Midori_rounds_mul_input3[51]), .B(
        Midori_rounds_mul_input3[55]), .ZN(Midori_rounds_mul3_MC1_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U4 ( .A(Midori_rounds_mul_input3[62]), .B(
        Midori_rounds_mul3_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result3[22]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U3 ( .A(Midori_rounds_mul_input3[50]), .B(
        Midori_rounds_mul_input3[54]), .ZN(Midori_rounds_mul3_MC1_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U2 ( .A(Midori_rounds_mul_input3[52]), .B(
        Midori_rounds_mul3_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result3[0]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U1 ( .A(Midori_rounds_mul_input3[60]), .B(
        Midori_rounds_mul_input3[56]), .ZN(Midori_rounds_mul3_MC1_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U24 ( .A(Midori_rounds_mul_input3[45]), .B(
        Midori_rounds_mul3_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result3[45]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U23 ( .A(Midori_rounds_mul_input3[44]), .B(
        Midori_rounds_mul3_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result3[44]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U22 ( .A(Midori_rounds_mul_input3[35]), .B(
        Midori_rounds_mul3_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result3[19]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U21 ( .A(Midori_rounds_mul_input3[34]), .B(
        Midori_rounds_mul3_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result3[18]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U20 ( .A(Midori_rounds_mul_input3[33]), .B(
        Midori_rounds_mul3_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result3[17]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U19 ( .A(Midori_rounds_mul_input3[32]), .B(
        Midori_rounds_mul3_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result3[16]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U18 ( .A(Midori_rounds_mul_input3[39]), .B(
        Midori_rounds_mul3_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result3[59]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U17 ( .A(Midori_rounds_mul_input3[47]), .B(
        Midori_rounds_mul_input3[43]), .ZN(Midori_rounds_mul3_MC2_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U16 ( .A(Midori_rounds_mul_input3[38]), .B(
        Midori_rounds_mul3_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result3[58]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U15 ( .A(Midori_rounds_mul_input3[46]), .B(
        Midori_rounds_mul_input3[42]), .ZN(Midori_rounds_mul3_MC2_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U14 ( .A(Midori_rounds_mul_input3[37]), .B(
        Midori_rounds_mul3_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result3[57]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U13 ( .A(Midori_rounds_mul_input3[41]), .B(
        Midori_rounds_mul_input3[45]), .ZN(Midori_rounds_mul3_MC2_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U12 ( .A(Midori_rounds_mul_input3[43]), .B(
        Midori_rounds_mul3_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result3[7]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U11 ( .A(Midori_rounds_mul_input3[42]), .B(
        Midori_rounds_mul3_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result3[6]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U10 ( .A(Midori_rounds_mul_input3[41]), .B(
        Midori_rounds_mul3_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result3[5]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U9 ( .A(Midori_rounds_mul_input3[33]), .B(
        Midori_rounds_mul_input3[37]), .ZN(Midori_rounds_mul3_MC2_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U8 ( .A(Midori_rounds_mul_input3[40]), .B(
        Midori_rounds_mul3_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result3[4]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U7 ( .A(Midori_rounds_mul_input3[36]), .B(
        Midori_rounds_mul_input3[32]), .ZN(Midori_rounds_mul3_MC2_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U6 ( .A(Midori_rounds_mul_input3[47]), .B(
        Midori_rounds_mul3_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result3[47]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U5 ( .A(Midori_rounds_mul_input3[35]), .B(
        Midori_rounds_mul_input3[39]), .ZN(Midori_rounds_mul3_MC2_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U4 ( .A(Midori_rounds_mul_input3[46]), .B(
        Midori_rounds_mul3_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result3[46]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U3 ( .A(Midori_rounds_mul_input3[34]), .B(
        Midori_rounds_mul_input3[38]), .ZN(Midori_rounds_mul3_MC2_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U2 ( .A(Midori_rounds_mul_input3[36]), .B(
        Midori_rounds_mul3_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result3[56]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U1 ( .A(Midori_rounds_mul_input3[44]), .B(
        Midori_rounds_mul_input3[40]), .ZN(Midori_rounds_mul3_MC2_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U24 ( .A(Midori_rounds_mul_input3[29]), .B(
        Midori_rounds_mul3_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result3[49]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U23 ( .A(Midori_rounds_mul_input3[28]), .B(
        Midori_rounds_mul3_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result3[48]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U22 ( .A(Midori_rounds_mul_input3[19]), .B(
        Midori_rounds_mul3_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result3[15]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U21 ( .A(Midori_rounds_mul_input3[18]), .B(
        Midori_rounds_mul3_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result3[14]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U20 ( .A(Midori_rounds_mul_input3[17]), .B(
        Midori_rounds_mul3_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result3[13]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U19 ( .A(Midori_rounds_mul_input3[16]), .B(
        Midori_rounds_mul3_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result3[12]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U18 ( .A(Midori_rounds_mul_input3[23]), .B(
        Midori_rounds_mul3_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result3[39]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U17 ( .A(Midori_rounds_mul_input3[31]), .B(
        Midori_rounds_mul_input3[27]), .ZN(Midori_rounds_mul3_MC3_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U16 ( .A(Midori_rounds_mul_input3[22]), .B(
        Midori_rounds_mul3_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result3[38]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U15 ( .A(Midori_rounds_mul_input3[30]), .B(
        Midori_rounds_mul_input3[26]), .ZN(Midori_rounds_mul3_MC3_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U14 ( .A(Midori_rounds_mul_input3[21]), .B(
        Midori_rounds_mul3_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result3[37]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U13 ( .A(Midori_rounds_mul_input3[25]), .B(
        Midori_rounds_mul_input3[29]), .ZN(Midori_rounds_mul3_MC3_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U12 ( .A(Midori_rounds_mul_input3[27]), .B(
        Midori_rounds_mul3_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result3[27]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U11 ( .A(Midori_rounds_mul_input3[26]), .B(
        Midori_rounds_mul3_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result3[26]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U10 ( .A(Midori_rounds_mul_input3[25]), .B(
        Midori_rounds_mul3_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result3[25]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U9 ( .A(Midori_rounds_mul_input3[17]), .B(
        Midori_rounds_mul_input3[21]), .ZN(Midori_rounds_mul3_MC3_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U8 ( .A(Midori_rounds_mul_input3[24]), .B(
        Midori_rounds_mul3_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result3[24]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U7 ( .A(Midori_rounds_mul_input3[20]), .B(
        Midori_rounds_mul_input3[16]), .ZN(Midori_rounds_mul3_MC3_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U6 ( .A(Midori_rounds_mul_input3[31]), .B(
        Midori_rounds_mul3_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result3[51]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U5 ( .A(Midori_rounds_mul_input3[19]), .B(
        Midori_rounds_mul_input3[23]), .ZN(Midori_rounds_mul3_MC3_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U4 ( .A(Midori_rounds_mul_input3[30]), .B(
        Midori_rounds_mul3_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result3[50]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U3 ( .A(Midori_rounds_mul_input3[18]), .B(
        Midori_rounds_mul_input3[22]), .ZN(Midori_rounds_mul3_MC3_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U2 ( .A(Midori_rounds_mul_input3[20]), .B(
        Midori_rounds_mul3_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result3[36]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U1 ( .A(Midori_rounds_mul_input3[28]), .B(
        Midori_rounds_mul_input3[24]), .ZN(Midori_rounds_mul3_MC3_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U24 ( .A(Midori_rounds_mul_input3[13]), .B(
        Midori_rounds_mul3_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result3[9]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U23 ( .A(Midori_rounds_mul_input3[12]), .B(
        Midori_rounds_mul3_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result3[8]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U22 ( .A(Midori_rounds_mul_input3[3]), .B(
        Midori_rounds_mul3_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result3[55]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U21 ( .A(Midori_rounds_mul_input3[2]), .B(
        Midori_rounds_mul3_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result3[54]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U20 ( .A(Midori_rounds_mul_input3[1]), .B(
        Midori_rounds_mul3_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result3[53]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U19 ( .A(Midori_rounds_mul_input3[0]), .B(
        Midori_rounds_mul3_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result3[52]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U18 ( .A(Midori_rounds_mul_input3[7]), .B(
        Midori_rounds_mul3_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result3[31]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U17 ( .A(Midori_rounds_mul_input3[15]), .B(
        Midori_rounds_mul_input3[11]), .ZN(Midori_rounds_mul3_MC4_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U16 ( .A(Midori_rounds_mul_input3[6]), .B(
        Midori_rounds_mul3_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result3[30]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U15 ( .A(Midori_rounds_mul_input3[14]), .B(
        Midori_rounds_mul_input3[10]), .ZN(Midori_rounds_mul3_MC4_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U14 ( .A(Midori_rounds_mul_input3[5]), .B(
        Midori_rounds_mul3_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result3[29]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U13 ( .A(Midori_rounds_mul_input3[9]), .B(
        Midori_rounds_mul_input3[13]), .ZN(Midori_rounds_mul3_MC4_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U12 ( .A(Midori_rounds_mul_input3[11]), .B(
        Midori_rounds_mul3_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result3[35]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U11 ( .A(Midori_rounds_mul_input3[10]), .B(
        Midori_rounds_mul3_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result3[34]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U10 ( .A(Midori_rounds_mul_input3[9]), .B(
        Midori_rounds_mul3_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result3[33]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U9 ( .A(Midori_rounds_mul_input3[1]), .B(
        Midori_rounds_mul_input3[5]), .ZN(Midori_rounds_mul3_MC4_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U8 ( .A(Midori_rounds_mul_input3[8]), .B(
        Midori_rounds_mul3_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result3[32]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U7 ( .A(Midori_rounds_mul_input3[4]), .B(
        Midori_rounds_mul_input3[0]), .ZN(Midori_rounds_mul3_MC4_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U6 ( .A(Midori_rounds_mul_input3[15]), .B(
        Midori_rounds_mul3_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result3[11]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U5 ( .A(Midori_rounds_mul_input3[3]), .B(
        Midori_rounds_mul_input3[7]), .ZN(Midori_rounds_mul3_MC4_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U4 ( .A(Midori_rounds_mul_input3[14]), .B(
        Midori_rounds_mul3_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result3[10]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U3 ( .A(Midori_rounds_mul_input3[2]), .B(
        Midori_rounds_mul_input3[6]), .ZN(Midori_rounds_mul3_MC4_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U2 ( .A(Midori_rounds_mul_input3[4]), .B(
        Midori_rounds_mul3_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result3[28]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U1 ( .A(Midori_rounds_mul_input3[12]), .B(
        Midori_rounds_mul_input3[8]), .ZN(Midori_rounds_mul3_MC4_n19) );
endmodule
